
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_671 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_671;

architecture SYN_full_adder_arch of FullAdder_671 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_670 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_670;

architecture SYN_full_adder_arch of FullAdder_670 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_669 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_669;

architecture SYN_full_adder_arch of FullAdder_669 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_668 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_668;

architecture SYN_full_adder_arch of FullAdder_668 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_667 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_667;

architecture SYN_full_adder_arch of FullAdder_667 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_666 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_666;

architecture SYN_full_adder_arch of FullAdder_666 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_665 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_665;

architecture SYN_full_adder_arch of FullAdder_665 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_664 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_664;

architecture SYN_full_adder_arch of FullAdder_664 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_663 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_663;

architecture SYN_full_adder_arch of FullAdder_663 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_662 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_662;

architecture SYN_full_adder_arch of FullAdder_662 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_661 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_661;

architecture SYN_full_adder_arch of FullAdder_661 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_660 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_660;

architecture SYN_full_adder_arch of FullAdder_660 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_659 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_659;

architecture SYN_full_adder_arch of FullAdder_659 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_658 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_658;

architecture SYN_full_adder_arch of FullAdder_658 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_657 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_657;

architecture SYN_full_adder_arch of FullAdder_657 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_656 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_656;

architecture SYN_full_adder_arch of FullAdder_656 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_655 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_655;

architecture SYN_full_adder_arch of FullAdder_655 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_654 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_654;

architecture SYN_full_adder_arch of FullAdder_654 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_653 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_653;

architecture SYN_full_adder_arch of FullAdder_653 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_652 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_652;

architecture SYN_full_adder_arch of FullAdder_652 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_651 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_651;

architecture SYN_full_adder_arch of FullAdder_651 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_650 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_650;

architecture SYN_full_adder_arch of FullAdder_650 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_649 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_649;

architecture SYN_full_adder_arch of FullAdder_649 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_648 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_648;

architecture SYN_full_adder_arch of FullAdder_648 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_647 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_647;

architecture SYN_full_adder_arch of FullAdder_647 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_646 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_646;

architecture SYN_full_adder_arch of FullAdder_646 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_645 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_645;

architecture SYN_full_adder_arch of FullAdder_645 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_644 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_644;

architecture SYN_full_adder_arch of FullAdder_644 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_643 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_643;

architecture SYN_full_adder_arch of FullAdder_643 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_642 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_642;

architecture SYN_full_adder_arch of FullAdder_642 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_641 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_641;

architecture SYN_full_adder_arch of FullAdder_641 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_640 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_640;

architecture SYN_full_adder_arch of FullAdder_640 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_639 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_639;

architecture SYN_full_adder_arch of FullAdder_639 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_638 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_638;

architecture SYN_full_adder_arch of FullAdder_638 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_637 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_637;

architecture SYN_full_adder_arch of FullAdder_637 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_636 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_636;

architecture SYN_full_adder_arch of FullAdder_636 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_635 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_635;

architecture SYN_full_adder_arch of FullAdder_635 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_634 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_634;

architecture SYN_full_adder_arch of FullAdder_634 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_633 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_633;

architecture SYN_full_adder_arch of FullAdder_633 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_632 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_632;

architecture SYN_full_adder_arch of FullAdder_632 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_631 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_631;

architecture SYN_full_adder_arch of FullAdder_631 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_630 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_630;

architecture SYN_full_adder_arch of FullAdder_630 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_629 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_629;

architecture SYN_full_adder_arch of FullAdder_629 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_628 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_628;

architecture SYN_full_adder_arch of FullAdder_628 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_627 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_627;

architecture SYN_full_adder_arch of FullAdder_627 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_626 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_626;

architecture SYN_full_adder_arch of FullAdder_626 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_625 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_625;

architecture SYN_full_adder_arch of FullAdder_625 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_624 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_624;

architecture SYN_full_adder_arch of FullAdder_624 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_623 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_623;

architecture SYN_full_adder_arch of FullAdder_623 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_622 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_622;

architecture SYN_full_adder_arch of FullAdder_622 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_621 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_621;

architecture SYN_full_adder_arch of FullAdder_621 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_620 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_620;

architecture SYN_full_adder_arch of FullAdder_620 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_619 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_619;

architecture SYN_full_adder_arch of FullAdder_619 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_618 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_618;

architecture SYN_full_adder_arch of FullAdder_618 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_617 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_617;

architecture SYN_full_adder_arch of FullAdder_617 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_616 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_616;

architecture SYN_full_adder_arch of FullAdder_616 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => ci, Z => s);
   U1 : INV_X1 port map( A => b, ZN => n6);
   U2 : CLKBUF_X1 port map( A => n8, Z => n4);
   U4 : CLKBUF_X1 port map( A => a, Z => n5);
   U5 : XNOR2_X1 port map( A => a, B => n6, ZN => n8);
   U6 : INV_X1 port map( A => n7, ZN => co);
   U7 : AOI22_X1 port map( A1 => b, A2 => n5, B1 => n8, B2 => ci, ZN => n7);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_615 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_615;

architecture SYN_full_adder_arch of FullAdder_615 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n5, B => n7, Z => s);
   U1 : INV_X1 port map( A => b, ZN => n4);
   U2 : XNOR2_X1 port map( A => a, B => n4, ZN => n7);
   U4 : CLKBUF_X1 port map( A => ci, Z => n5);
   U5 : AOI22_X1 port map( A1 => b, A2 => a, B1 => ci, B2 => n7, ZN => n6);
   U6 : INV_X1 port map( A => n6, ZN => co);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_614 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_614;

architecture SYN_full_adder_arch of FullAdder_614 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : AOI22_X1 port map( A1 => b, A2 => a, B1 => ci, B2 => n5, ZN => n4);
   U2 : INV_X1 port map( A => n4, ZN => co);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_613 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_613;

architecture SYN_full_adder_arch of FullAdder_613 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => a, B => b, Z => n6);
   U1 : INV_X1 port map( A => n6, ZN => n4);
   U2 : XNOR2_X1 port map( A => ci, B => n4, ZN => s);
   U3 : INV_X1 port map( A => n5, ZN => co);
   U5 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n6, B2 => ci, ZN => n5);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_612 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_612;

architecture SYN_full_adder_arch of FullAdder_612 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => n4, B => ci, Z => s);
   U1 : INV_X1 port map( A => b, ZN => n5);
   U2 : XNOR2_X1 port map( A => n6, B => n5, ZN => n4);
   U4 : XNOR2_X1 port map( A => a, B => n5, ZN => n8);
   U5 : CLKBUF_X1 port map( A => a, Z => n6);
   U6 : AOI22_X1 port map( A1 => b, A2 => n6, B1 => n8, B2 => ci, ZN => n7);
   U7 : INV_X1 port map( A => n7, ZN => co);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_611 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_611;

architecture SYN_full_adder_arch of FullAdder_611 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n5, n6, n7 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n7, Z => s);
   U1 : INV_X1 port map( A => b, ZN => n3);
   U2 : XNOR2_X1 port map( A => a, B => n3, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => co);
   U5 : NAND2_X1 port map( A1 => b, A2 => a, ZN => n5);
   U6 : NAND2_X1 port map( A1 => ci, A2 => n7, ZN => n6);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_610 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_610;

architecture SYN_full_adder_arch of FullAdder_610 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => ci, B2 => n5, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_609 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_609;

architecture SYN_full_adder_arch of FullAdder_609 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U4 : XOR2_X1 port map( A => a, B => b, Z => n9);
   U1 : NAND2_X1 port map( A1 => ci, A2 => n7, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n4, A2 => n9, ZN => n6);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => s);
   U5 : INV_X1 port map( A => ci, ZN => n4);
   U6 : INV_X1 port map( A => n9, ZN => n7);
   U7 : INV_X1 port map( A => n8, ZN => co);
   U8 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n9, B2 => ci, ZN => n8);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_608 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_608;

architecture SYN_full_adder_arch of FullAdder_608 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_607 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_607;

architecture SYN_full_adder_arch of FullAdder_607 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_606 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_606;

architecture SYN_full_adder_arch of FullAdder_606 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_605 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_605;

architecture SYN_full_adder_arch of FullAdder_605 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_604 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_604;

architecture SYN_full_adder_arch of FullAdder_604 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_603 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_603;

architecture SYN_full_adder_arch of FullAdder_603 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_602 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_602;

architecture SYN_full_adder_arch of FullAdder_602 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_601 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_601;

architecture SYN_full_adder_arch of FullAdder_601 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_600 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_600;

architecture SYN_full_adder_arch of FullAdder_600 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_599 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_599;

architecture SYN_full_adder_arch of FullAdder_599 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_598 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_598;

architecture SYN_full_adder_arch of FullAdder_598 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_597 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_597;

architecture SYN_full_adder_arch of FullAdder_597 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_596 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_596;

architecture SYN_full_adder_arch of FullAdder_596 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_595 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_595;

architecture SYN_full_adder_arch of FullAdder_595 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_594 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_594;

architecture SYN_full_adder_arch of FullAdder_594 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_593 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_593;

architecture SYN_full_adder_arch of FullAdder_593 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_592 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_592;

architecture SYN_full_adder_arch of FullAdder_592 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_591 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_591;

architecture SYN_full_adder_arch of FullAdder_591 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_590 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_590;

architecture SYN_full_adder_arch of FullAdder_590 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_589 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_589;

architecture SYN_full_adder_arch of FullAdder_589 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_588 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_588;

architecture SYN_full_adder_arch of FullAdder_588 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_587 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_587;

architecture SYN_full_adder_arch of FullAdder_587 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_586 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_586;

architecture SYN_full_adder_arch of FullAdder_586 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_585 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_585;

architecture SYN_full_adder_arch of FullAdder_585 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_584 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_584;

architecture SYN_full_adder_arch of FullAdder_584 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_583 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_583;

architecture SYN_full_adder_arch of FullAdder_583 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_582 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_582;

architecture SYN_full_adder_arch of FullAdder_582 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_581 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_581;

architecture SYN_full_adder_arch of FullAdder_581 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_580 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_580;

architecture SYN_full_adder_arch of FullAdder_580 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_579 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_579;

architecture SYN_full_adder_arch of FullAdder_579 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_578 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_578;

architecture SYN_full_adder_arch of FullAdder_578 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_577 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_577;

architecture SYN_full_adder_arch of FullAdder_577 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_576 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_576;

architecture SYN_full_adder_arch of FullAdder_576 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_575 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_575;

architecture SYN_full_adder_arch of FullAdder_575 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_574 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_574;

architecture SYN_full_adder_arch of FullAdder_574 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_573 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_573;

architecture SYN_full_adder_arch of FullAdder_573 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_572 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_572;

architecture SYN_full_adder_arch of FullAdder_572 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_571 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_571;

architecture SYN_full_adder_arch of FullAdder_571 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_570 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_570;

architecture SYN_full_adder_arch of FullAdder_570 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_569 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_569;

architecture SYN_full_adder_arch of FullAdder_569 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_568 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_568;

architecture SYN_full_adder_arch of FullAdder_568 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_567 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_567;

architecture SYN_full_adder_arch of FullAdder_567 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_566 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_566;

architecture SYN_full_adder_arch of FullAdder_566 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_565 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_565;

architecture SYN_full_adder_arch of FullAdder_565 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_564 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_564;

architecture SYN_full_adder_arch of FullAdder_564 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_563 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_563;

architecture SYN_full_adder_arch of FullAdder_563 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_562 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_562;

architecture SYN_full_adder_arch of FullAdder_562 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_561 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_561;

architecture SYN_full_adder_arch of FullAdder_561 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_560 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_560;

architecture SYN_full_adder_arch of FullAdder_560 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_559 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_559;

architecture SYN_full_adder_arch of FullAdder_559 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_558 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_558;

architecture SYN_full_adder_arch of FullAdder_558 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_557 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_557;

architecture SYN_full_adder_arch of FullAdder_557 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_556 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_556;

architecture SYN_full_adder_arch of FullAdder_556 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_555 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_555;

architecture SYN_full_adder_arch of FullAdder_555 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_554 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_554;

architecture SYN_full_adder_arch of FullAdder_554 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_553 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_553;

architecture SYN_full_adder_arch of FullAdder_553 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_552 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_552;

architecture SYN_full_adder_arch of FullAdder_552 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_551 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_551;

architecture SYN_full_adder_arch of FullAdder_551 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_550 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_550;

architecture SYN_full_adder_arch of FullAdder_550 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_549 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_549;

architecture SYN_full_adder_arch of FullAdder_549 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_548 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_548;

architecture SYN_full_adder_arch of FullAdder_548 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_547 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_547;

architecture SYN_full_adder_arch of FullAdder_547 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_546 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_546;

architecture SYN_full_adder_arch of FullAdder_546 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_545 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_545;

architecture SYN_full_adder_arch of FullAdder_545 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_544 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_544;

architecture SYN_full_adder_arch of FullAdder_544 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_543 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_543;

architecture SYN_full_adder_arch of FullAdder_543 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_542 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_542;

architecture SYN_full_adder_arch of FullAdder_542 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_541 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_541;

architecture SYN_full_adder_arch of FullAdder_541 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_540 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_540;

architecture SYN_full_adder_arch of FullAdder_540 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_539 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_539;

architecture SYN_full_adder_arch of FullAdder_539 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_538 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_538;

architecture SYN_full_adder_arch of FullAdder_538 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_537 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_537;

architecture SYN_full_adder_arch of FullAdder_537 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_536 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_536;

architecture SYN_full_adder_arch of FullAdder_536 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_535 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_535;

architecture SYN_full_adder_arch of FullAdder_535 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_534 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_534;

architecture SYN_full_adder_arch of FullAdder_534 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_533 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_533;

architecture SYN_full_adder_arch of FullAdder_533 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_532 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_532;

architecture SYN_full_adder_arch of FullAdder_532 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_531 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_531;

architecture SYN_full_adder_arch of FullAdder_531 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_530 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_530;

architecture SYN_full_adder_arch of FullAdder_530 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_529 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_529;

architecture SYN_full_adder_arch of FullAdder_529 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_528 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_528;

architecture SYN_full_adder_arch of FullAdder_528 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_527 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_527;

architecture SYN_full_adder_arch of FullAdder_527 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_526 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_526;

architecture SYN_full_adder_arch of FullAdder_526 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_525 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_525;

architecture SYN_full_adder_arch of FullAdder_525 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_524 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_524;

architecture SYN_full_adder_arch of FullAdder_524 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_523 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_523;

architecture SYN_full_adder_arch of FullAdder_523 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_522 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_522;

architecture SYN_full_adder_arch of FullAdder_522 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_521 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_521;

architecture SYN_full_adder_arch of FullAdder_521 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_520 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_520;

architecture SYN_full_adder_arch of FullAdder_520 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_519 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_519;

architecture SYN_full_adder_arch of FullAdder_519 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_518 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_518;

architecture SYN_full_adder_arch of FullAdder_518 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_517 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_517;

architecture SYN_full_adder_arch of FullAdder_517 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_516 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_516;

architecture SYN_full_adder_arch of FullAdder_516 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_515 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_515;

architecture SYN_full_adder_arch of FullAdder_515 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_514 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_514;

architecture SYN_full_adder_arch of FullAdder_514 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_513 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_513;

architecture SYN_full_adder_arch of FullAdder_513 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_512 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_512;

architecture SYN_full_adder_arch of FullAdder_512 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_511 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_511;

architecture SYN_full_adder_arch of FullAdder_511 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_510 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_510;

architecture SYN_full_adder_arch of FullAdder_510 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_509 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_509;

architecture SYN_full_adder_arch of FullAdder_509 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_508 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_508;

architecture SYN_full_adder_arch of FullAdder_508 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_507 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_507;

architecture SYN_full_adder_arch of FullAdder_507 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_506 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_506;

architecture SYN_full_adder_arch of FullAdder_506 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_505 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_505;

architecture SYN_full_adder_arch of FullAdder_505 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_504 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_504;

architecture SYN_full_adder_arch of FullAdder_504 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_503 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_503;

architecture SYN_full_adder_arch of FullAdder_503 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_502 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_502;

architecture SYN_full_adder_arch of FullAdder_502 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_501 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_501;

architecture SYN_full_adder_arch of FullAdder_501 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_500 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_500;

architecture SYN_full_adder_arch of FullAdder_500 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_499 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_499;

architecture SYN_full_adder_arch of FullAdder_499 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_498 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_498;

architecture SYN_full_adder_arch of FullAdder_498 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_497 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_497;

architecture SYN_full_adder_arch of FullAdder_497 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_496 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_496;

architecture SYN_full_adder_arch of FullAdder_496 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_495 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_495;

architecture SYN_full_adder_arch of FullAdder_495 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_494 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_494;

architecture SYN_full_adder_arch of FullAdder_494 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_493 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_493;

architecture SYN_full_adder_arch of FullAdder_493 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_492 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_492;

architecture SYN_full_adder_arch of FullAdder_492 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_491 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_491;

architecture SYN_full_adder_arch of FullAdder_491 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_490 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_490;

architecture SYN_full_adder_arch of FullAdder_490 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_489 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_489;

architecture SYN_full_adder_arch of FullAdder_489 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_488 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_488;

architecture SYN_full_adder_arch of FullAdder_488 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_487 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_487;

architecture SYN_full_adder_arch of FullAdder_487 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_486 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_486;

architecture SYN_full_adder_arch of FullAdder_486 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_485 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_485;

architecture SYN_full_adder_arch of FullAdder_485 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_484 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_484;

architecture SYN_full_adder_arch of FullAdder_484 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_483 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_483;

architecture SYN_full_adder_arch of FullAdder_483 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_482 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_482;

architecture SYN_full_adder_arch of FullAdder_482 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_481 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_481;

architecture SYN_full_adder_arch of FullAdder_481 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_480 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_480;

architecture SYN_full_adder_arch of FullAdder_480 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_479 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_479;

architecture SYN_full_adder_arch of FullAdder_479 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_478 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_478;

architecture SYN_full_adder_arch of FullAdder_478 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_477 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_477;

architecture SYN_full_adder_arch of FullAdder_477 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_476 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_476;

architecture SYN_full_adder_arch of FullAdder_476 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_475 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_475;

architecture SYN_full_adder_arch of FullAdder_475 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_474 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_474;

architecture SYN_full_adder_arch of FullAdder_474 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_473 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_473;

architecture SYN_full_adder_arch of FullAdder_473 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_472 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_472;

architecture SYN_full_adder_arch of FullAdder_472 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_471 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_471;

architecture SYN_full_adder_arch of FullAdder_471 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_470 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_470;

architecture SYN_full_adder_arch of FullAdder_470 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_469 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_469;

architecture SYN_full_adder_arch of FullAdder_469 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_468 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_468;

architecture SYN_full_adder_arch of FullAdder_468 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_467 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_467;

architecture SYN_full_adder_arch of FullAdder_467 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_466 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_466;

architecture SYN_full_adder_arch of FullAdder_466 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_465 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_465;

architecture SYN_full_adder_arch of FullAdder_465 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_464 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_464;

architecture SYN_full_adder_arch of FullAdder_464 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_463 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_463;

architecture SYN_full_adder_arch of FullAdder_463 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_462 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_462;

architecture SYN_full_adder_arch of FullAdder_462 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_461 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_461;

architecture SYN_full_adder_arch of FullAdder_461 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_460 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_460;

architecture SYN_full_adder_arch of FullAdder_460 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_459 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_459;

architecture SYN_full_adder_arch of FullAdder_459 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_458 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_458;

architecture SYN_full_adder_arch of FullAdder_458 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_457 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_457;

architecture SYN_full_adder_arch of FullAdder_457 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_456 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_456;

architecture SYN_full_adder_arch of FullAdder_456 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_455 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_455;

architecture SYN_full_adder_arch of FullAdder_455 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_454 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_454;

architecture SYN_full_adder_arch of FullAdder_454 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_453 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_453;

architecture SYN_full_adder_arch of FullAdder_453 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_452 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_452;

architecture SYN_full_adder_arch of FullAdder_452 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_451 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_451;

architecture SYN_full_adder_arch of FullAdder_451 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_450 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_450;

architecture SYN_full_adder_arch of FullAdder_450 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_449 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_449;

architecture SYN_full_adder_arch of FullAdder_449 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_448 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_448;

architecture SYN_full_adder_arch of FullAdder_448 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_447 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_447;

architecture SYN_full_adder_arch of FullAdder_447 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_446 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_446;

architecture SYN_full_adder_arch of FullAdder_446 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_445 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_445;

architecture SYN_full_adder_arch of FullAdder_445 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_444 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_444;

architecture SYN_full_adder_arch of FullAdder_444 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_443 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_443;

architecture SYN_full_adder_arch of FullAdder_443 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_442 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_442;

architecture SYN_full_adder_arch of FullAdder_442 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_441 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_441;

architecture SYN_full_adder_arch of FullAdder_441 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_440 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_440;

architecture SYN_full_adder_arch of FullAdder_440 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_439 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_439;

architecture SYN_full_adder_arch of FullAdder_439 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_438 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_438;

architecture SYN_full_adder_arch of FullAdder_438 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_437 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_437;

architecture SYN_full_adder_arch of FullAdder_437 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_436 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_436;

architecture SYN_full_adder_arch of FullAdder_436 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_435 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_435;

architecture SYN_full_adder_arch of FullAdder_435 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_434 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_434;

architecture SYN_full_adder_arch of FullAdder_434 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_433 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_433;

architecture SYN_full_adder_arch of FullAdder_433 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_432 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_432;

architecture SYN_full_adder_arch of FullAdder_432 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_431 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_431;

architecture SYN_full_adder_arch of FullAdder_431 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_430 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_430;

architecture SYN_full_adder_arch of FullAdder_430 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_429 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_429;

architecture SYN_full_adder_arch of FullAdder_429 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_428 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_428;

architecture SYN_full_adder_arch of FullAdder_428 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_427 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_427;

architecture SYN_full_adder_arch of FullAdder_427 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_426 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_426;

architecture SYN_full_adder_arch of FullAdder_426 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_425 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_425;

architecture SYN_full_adder_arch of FullAdder_425 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_424 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_424;

architecture SYN_full_adder_arch of FullAdder_424 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_423 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_423;

architecture SYN_full_adder_arch of FullAdder_423 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_422 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_422;

architecture SYN_full_adder_arch of FullAdder_422 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_421 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_421;

architecture SYN_full_adder_arch of FullAdder_421 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_420 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_420;

architecture SYN_full_adder_arch of FullAdder_420 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_419 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_419;

architecture SYN_full_adder_arch of FullAdder_419 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_418 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_418;

architecture SYN_full_adder_arch of FullAdder_418 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_417 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_417;

architecture SYN_full_adder_arch of FullAdder_417 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_416 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_416;

architecture SYN_full_adder_arch of FullAdder_416 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_415 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_415;

architecture SYN_full_adder_arch of FullAdder_415 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_414 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_414;

architecture SYN_full_adder_arch of FullAdder_414 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_413 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_413;

architecture SYN_full_adder_arch of FullAdder_413 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_412 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_412;

architecture SYN_full_adder_arch of FullAdder_412 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_411 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_411;

architecture SYN_full_adder_arch of FullAdder_411 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_410 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_410;

architecture SYN_full_adder_arch of FullAdder_410 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_409 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_409;

architecture SYN_full_adder_arch of FullAdder_409 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_408 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_408;

architecture SYN_full_adder_arch of FullAdder_408 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_407 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_407;

architecture SYN_full_adder_arch of FullAdder_407 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_406 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_406;

architecture SYN_full_adder_arch of FullAdder_406 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_405 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_405;

architecture SYN_full_adder_arch of FullAdder_405 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_404 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_404;

architecture SYN_full_adder_arch of FullAdder_404 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_403 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_403;

architecture SYN_full_adder_arch of FullAdder_403 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_402 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_402;

architecture SYN_full_adder_arch of FullAdder_402 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_401 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_401;

architecture SYN_full_adder_arch of FullAdder_401 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_400 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_400;

architecture SYN_full_adder_arch of FullAdder_400 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_399 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_399;

architecture SYN_full_adder_arch of FullAdder_399 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_398 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_398;

architecture SYN_full_adder_arch of FullAdder_398 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_397 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_397;

architecture SYN_full_adder_arch of FullAdder_397 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_396 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_396;

architecture SYN_full_adder_arch of FullAdder_396 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_395 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_395;

architecture SYN_full_adder_arch of FullAdder_395 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_394 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_394;

architecture SYN_full_adder_arch of FullAdder_394 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_393 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_393;

architecture SYN_full_adder_arch of FullAdder_393 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_392 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_392;

architecture SYN_full_adder_arch of FullAdder_392 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_391 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_391;

architecture SYN_full_adder_arch of FullAdder_391 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_390 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_390;

architecture SYN_full_adder_arch of FullAdder_390 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_389 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_389;

architecture SYN_full_adder_arch of FullAdder_389 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_388 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_388;

architecture SYN_full_adder_arch of FullAdder_388 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_387 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_387;

architecture SYN_full_adder_arch of FullAdder_387 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_386 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_386;

architecture SYN_full_adder_arch of FullAdder_386 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_385 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_385;

architecture SYN_full_adder_arch of FullAdder_385 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_384 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_384;

architecture SYN_full_adder_arch of FullAdder_384 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_383 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_383;

architecture SYN_full_adder_arch of FullAdder_383 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_382 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_382;

architecture SYN_full_adder_arch of FullAdder_382 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_381 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_381;

architecture SYN_full_adder_arch of FullAdder_381 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_380 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_380;

architecture SYN_full_adder_arch of FullAdder_380 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_379 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_379;

architecture SYN_full_adder_arch of FullAdder_379 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_378 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_378;

architecture SYN_full_adder_arch of FullAdder_378 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_377 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_377;

architecture SYN_full_adder_arch of FullAdder_377 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_376 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_376;

architecture SYN_full_adder_arch of FullAdder_376 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_375 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_375;

architecture SYN_full_adder_arch of FullAdder_375 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_374 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_374;

architecture SYN_full_adder_arch of FullAdder_374 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_373 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_373;

architecture SYN_full_adder_arch of FullAdder_373 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_372 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_372;

architecture SYN_full_adder_arch of FullAdder_372 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_371 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_371;

architecture SYN_full_adder_arch of FullAdder_371 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_370 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_370;

architecture SYN_full_adder_arch of FullAdder_370 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_369 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_369;

architecture SYN_full_adder_arch of FullAdder_369 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_368 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_368;

architecture SYN_full_adder_arch of FullAdder_368 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_367 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_367;

architecture SYN_full_adder_arch of FullAdder_367 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_366 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_366;

architecture SYN_full_adder_arch of FullAdder_366 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_365 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_365;

architecture SYN_full_adder_arch of FullAdder_365 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_364 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_364;

architecture SYN_full_adder_arch of FullAdder_364 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_363 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_363;

architecture SYN_full_adder_arch of FullAdder_363 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_362 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_362;

architecture SYN_full_adder_arch of FullAdder_362 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_361 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_361;

architecture SYN_full_adder_arch of FullAdder_361 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_360 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_360;

architecture SYN_full_adder_arch of FullAdder_360 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_359 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_359;

architecture SYN_full_adder_arch of FullAdder_359 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_358 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_358;

architecture SYN_full_adder_arch of FullAdder_358 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_357 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_357;

architecture SYN_full_adder_arch of FullAdder_357 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_356 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_356;

architecture SYN_full_adder_arch of FullAdder_356 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_355 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_355;

architecture SYN_full_adder_arch of FullAdder_355 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_354 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_354;

architecture SYN_full_adder_arch of FullAdder_354 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_353 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_353;

architecture SYN_full_adder_arch of FullAdder_353 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_352 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_352;

architecture SYN_full_adder_arch of FullAdder_352 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_351 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_351;

architecture SYN_full_adder_arch of FullAdder_351 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_350 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_350;

architecture SYN_full_adder_arch of FullAdder_350 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_349 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_349;

architecture SYN_full_adder_arch of FullAdder_349 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_348 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_348;

architecture SYN_full_adder_arch of FullAdder_348 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_347 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_347;

architecture SYN_full_adder_arch of FullAdder_347 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_346 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_346;

architecture SYN_full_adder_arch of FullAdder_346 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_345 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_345;

architecture SYN_full_adder_arch of FullAdder_345 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_344 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_344;

architecture SYN_full_adder_arch of FullAdder_344 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_343 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_343;

architecture SYN_full_adder_arch of FullAdder_343 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_342 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_342;

architecture SYN_full_adder_arch of FullAdder_342 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_341 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_341;

architecture SYN_full_adder_arch of FullAdder_341 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_340 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_340;

architecture SYN_full_adder_arch of FullAdder_340 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_339 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_339;

architecture SYN_full_adder_arch of FullAdder_339 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_338 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_338;

architecture SYN_full_adder_arch of FullAdder_338 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_337 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_337;

architecture SYN_full_adder_arch of FullAdder_337 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_336 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_336;

architecture SYN_full_adder_arch of FullAdder_336 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_335 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_335;

architecture SYN_full_adder_arch of FullAdder_335 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_334 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_334;

architecture SYN_full_adder_arch of FullAdder_334 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_333 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_333;

architecture SYN_full_adder_arch of FullAdder_333 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_332 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_332;

architecture SYN_full_adder_arch of FullAdder_332 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_331 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_331;

architecture SYN_full_adder_arch of FullAdder_331 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_330 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_330;

architecture SYN_full_adder_arch of FullAdder_330 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_329 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_329;

architecture SYN_full_adder_arch of FullAdder_329 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_328 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_328;

architecture SYN_full_adder_arch of FullAdder_328 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_327 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_327;

architecture SYN_full_adder_arch of FullAdder_327 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_326 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_326;

architecture SYN_full_adder_arch of FullAdder_326 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_325 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_325;

architecture SYN_full_adder_arch of FullAdder_325 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_324 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_324;

architecture SYN_full_adder_arch of FullAdder_324 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_323 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_323;

architecture SYN_full_adder_arch of FullAdder_323 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_322 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_322;

architecture SYN_full_adder_arch of FullAdder_322 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_321 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_321;

architecture SYN_full_adder_arch of FullAdder_321 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_320 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_320;

architecture SYN_full_adder_arch of FullAdder_320 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_319 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_319;

architecture SYN_full_adder_arch of FullAdder_319 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_318 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_318;

architecture SYN_full_adder_arch of FullAdder_318 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_317 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_317;

architecture SYN_full_adder_arch of FullAdder_317 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_316 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_316;

architecture SYN_full_adder_arch of FullAdder_316 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_315 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_315;

architecture SYN_full_adder_arch of FullAdder_315 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_314 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_314;

architecture SYN_full_adder_arch of FullAdder_314 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_313 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_313;

architecture SYN_full_adder_arch of FullAdder_313 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_312 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_312;

architecture SYN_full_adder_arch of FullAdder_312 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_311 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_311;

architecture SYN_full_adder_arch of FullAdder_311 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_310 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_310;

architecture SYN_full_adder_arch of FullAdder_310 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_309 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_309;

architecture SYN_full_adder_arch of FullAdder_309 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_308 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_308;

architecture SYN_full_adder_arch of FullAdder_308 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_307 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_307;

architecture SYN_full_adder_arch of FullAdder_307 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_306 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_306;

architecture SYN_full_adder_arch of FullAdder_306 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_305 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_305;

architecture SYN_full_adder_arch of FullAdder_305 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_304 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_304;

architecture SYN_full_adder_arch of FullAdder_304 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_303 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_303;

architecture SYN_full_adder_arch of FullAdder_303 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_302 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_302;

architecture SYN_full_adder_arch of FullAdder_302 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_301 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_301;

architecture SYN_full_adder_arch of FullAdder_301 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_300 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_300;

architecture SYN_full_adder_arch of FullAdder_300 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_299 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_299;

architecture SYN_full_adder_arch of FullAdder_299 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_298 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_298;

architecture SYN_full_adder_arch of FullAdder_298 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_297 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_297;

architecture SYN_full_adder_arch of FullAdder_297 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_296 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_296;

architecture SYN_full_adder_arch of FullAdder_296 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_295 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_295;

architecture SYN_full_adder_arch of FullAdder_295 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_294 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_294;

architecture SYN_full_adder_arch of FullAdder_294 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_293 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_293;

architecture SYN_full_adder_arch of FullAdder_293 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_292 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_292;

architecture SYN_full_adder_arch of FullAdder_292 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_291 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_291;

architecture SYN_full_adder_arch of FullAdder_291 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_290 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_290;

architecture SYN_full_adder_arch of FullAdder_290 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_289 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_289;

architecture SYN_full_adder_arch of FullAdder_289 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_288 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_288;

architecture SYN_full_adder_arch of FullAdder_288 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_287 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_287;

architecture SYN_full_adder_arch of FullAdder_287 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_286 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_286;

architecture SYN_full_adder_arch of FullAdder_286 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_285 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_285;

architecture SYN_full_adder_arch of FullAdder_285 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_284 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_284;

architecture SYN_full_adder_arch of FullAdder_284 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_283 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_283;

architecture SYN_full_adder_arch of FullAdder_283 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_282 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_282;

architecture SYN_full_adder_arch of FullAdder_282 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_281 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_281;

architecture SYN_full_adder_arch of FullAdder_281 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_280 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_280;

architecture SYN_full_adder_arch of FullAdder_280 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_279 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_279;

architecture SYN_full_adder_arch of FullAdder_279 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_278 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_278;

architecture SYN_full_adder_arch of FullAdder_278 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_277 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_277;

architecture SYN_full_adder_arch of FullAdder_277 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_276 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_276;

architecture SYN_full_adder_arch of FullAdder_276 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_275 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_275;

architecture SYN_full_adder_arch of FullAdder_275 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_274 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_274;

architecture SYN_full_adder_arch of FullAdder_274 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_273 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_273;

architecture SYN_full_adder_arch of FullAdder_273 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_272 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_272;

architecture SYN_full_adder_arch of FullAdder_272 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_271 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_271;

architecture SYN_full_adder_arch of FullAdder_271 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_270 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_270;

architecture SYN_full_adder_arch of FullAdder_270 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_269 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_269;

architecture SYN_full_adder_arch of FullAdder_269 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_268 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_268;

architecture SYN_full_adder_arch of FullAdder_268 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_267 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_267;

architecture SYN_full_adder_arch of FullAdder_267 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_266 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_266;

architecture SYN_full_adder_arch of FullAdder_266 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_265 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_265;

architecture SYN_full_adder_arch of FullAdder_265 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_264 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_264;

architecture SYN_full_adder_arch of FullAdder_264 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_263 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_263;

architecture SYN_full_adder_arch of FullAdder_263 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_262 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_262;

architecture SYN_full_adder_arch of FullAdder_262 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_261 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_261;

architecture SYN_full_adder_arch of FullAdder_261 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_260 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_260;

architecture SYN_full_adder_arch of FullAdder_260 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_259 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_259;

architecture SYN_full_adder_arch of FullAdder_259 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_258 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_258;

architecture SYN_full_adder_arch of FullAdder_258 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_257 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_257;

architecture SYN_full_adder_arch of FullAdder_257 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_256 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_256;

architecture SYN_full_adder_arch of FullAdder_256 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_255 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_255;

architecture SYN_full_adder_arch of FullAdder_255 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_254 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_254;

architecture SYN_full_adder_arch of FullAdder_254 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_253 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_253;

architecture SYN_full_adder_arch of FullAdder_253 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_252 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_252;

architecture SYN_full_adder_arch of FullAdder_252 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_251 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_251;

architecture SYN_full_adder_arch of FullAdder_251 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_250 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_250;

architecture SYN_full_adder_arch of FullAdder_250 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_249 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_249;

architecture SYN_full_adder_arch of FullAdder_249 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_248 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_248;

architecture SYN_full_adder_arch of FullAdder_248 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_247 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_247;

architecture SYN_full_adder_arch of FullAdder_247 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_246 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_246;

architecture SYN_full_adder_arch of FullAdder_246 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_245 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_245;

architecture SYN_full_adder_arch of FullAdder_245 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_244 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_244;

architecture SYN_full_adder_arch of FullAdder_244 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_243 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_243;

architecture SYN_full_adder_arch of FullAdder_243 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_242 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_242;

architecture SYN_full_adder_arch of FullAdder_242 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_241 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_241;

architecture SYN_full_adder_arch of FullAdder_241 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_240 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_240;

architecture SYN_full_adder_arch of FullAdder_240 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_239 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_239;

architecture SYN_full_adder_arch of FullAdder_239 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_238 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_238;

architecture SYN_full_adder_arch of FullAdder_238 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_237 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_237;

architecture SYN_full_adder_arch of FullAdder_237 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_236 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_236;

architecture SYN_full_adder_arch of FullAdder_236 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_235 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_235;

architecture SYN_full_adder_arch of FullAdder_235 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_234 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_234;

architecture SYN_full_adder_arch of FullAdder_234 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_233 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_233;

architecture SYN_full_adder_arch of FullAdder_233 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_232 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_232;

architecture SYN_full_adder_arch of FullAdder_232 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_231 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_231;

architecture SYN_full_adder_arch of FullAdder_231 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_230 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_230;

architecture SYN_full_adder_arch of FullAdder_230 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_229 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_229;

architecture SYN_full_adder_arch of FullAdder_229 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_228 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_228;

architecture SYN_full_adder_arch of FullAdder_228 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_227 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_227;

architecture SYN_full_adder_arch of FullAdder_227 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_226 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_226;

architecture SYN_full_adder_arch of FullAdder_226 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_225 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_225;

architecture SYN_full_adder_arch of FullAdder_225 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_224 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_224;

architecture SYN_full_adder_arch of FullAdder_224 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_223 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_223;

architecture SYN_full_adder_arch of FullAdder_223 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_222 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_222;

architecture SYN_full_adder_arch of FullAdder_222 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_221 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_221;

architecture SYN_full_adder_arch of FullAdder_221 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_220 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_220;

architecture SYN_full_adder_arch of FullAdder_220 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_219 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_219;

architecture SYN_full_adder_arch of FullAdder_219 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_218 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_218;

architecture SYN_full_adder_arch of FullAdder_218 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_217 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_217;

architecture SYN_full_adder_arch of FullAdder_217 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_216 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_216;

architecture SYN_full_adder_arch of FullAdder_216 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_215 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_215;

architecture SYN_full_adder_arch of FullAdder_215 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_214 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_214;

architecture SYN_full_adder_arch of FullAdder_214 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_213 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_213;

architecture SYN_full_adder_arch of FullAdder_213 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_212 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_212;

architecture SYN_full_adder_arch of FullAdder_212 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_211 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_211;

architecture SYN_full_adder_arch of FullAdder_211 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_210 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_210;

architecture SYN_full_adder_arch of FullAdder_210 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_209 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_209;

architecture SYN_full_adder_arch of FullAdder_209 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_208 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_208;

architecture SYN_full_adder_arch of FullAdder_208 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_207 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_207;

architecture SYN_full_adder_arch of FullAdder_207 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_206 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_206;

architecture SYN_full_adder_arch of FullAdder_206 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_205 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_205;

architecture SYN_full_adder_arch of FullAdder_205 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_204 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_204;

architecture SYN_full_adder_arch of FullAdder_204 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_203 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_203;

architecture SYN_full_adder_arch of FullAdder_203 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_202 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_202;

architecture SYN_full_adder_arch of FullAdder_202 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_201 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_201;

architecture SYN_full_adder_arch of FullAdder_201 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_200 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_200;

architecture SYN_full_adder_arch of FullAdder_200 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_199 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_199;

architecture SYN_full_adder_arch of FullAdder_199 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_198 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_198;

architecture SYN_full_adder_arch of FullAdder_198 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_197 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_197;

architecture SYN_full_adder_arch of FullAdder_197 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_196 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_196;

architecture SYN_full_adder_arch of FullAdder_196 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_195 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_195;

architecture SYN_full_adder_arch of FullAdder_195 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_194 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_194;

architecture SYN_full_adder_arch of FullAdder_194 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_193 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_193;

architecture SYN_full_adder_arch of FullAdder_193 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_192 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_192;

architecture SYN_full_adder_arch of FullAdder_192 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_191 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_191;

architecture SYN_full_adder_arch of FullAdder_191 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_190 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_190;

architecture SYN_full_adder_arch of FullAdder_190 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_189 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_189;

architecture SYN_full_adder_arch of FullAdder_189 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_188 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_188;

architecture SYN_full_adder_arch of FullAdder_188 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_187 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_187;

architecture SYN_full_adder_arch of FullAdder_187 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_186 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_186;

architecture SYN_full_adder_arch of FullAdder_186 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_185 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_185;

architecture SYN_full_adder_arch of FullAdder_185 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_184 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_184;

architecture SYN_full_adder_arch of FullAdder_184 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_183 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_183;

architecture SYN_full_adder_arch of FullAdder_183 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_182 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_182;

architecture SYN_full_adder_arch of FullAdder_182 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_181 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_181;

architecture SYN_full_adder_arch of FullAdder_181 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_180 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_180;

architecture SYN_full_adder_arch of FullAdder_180 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_179 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_179;

architecture SYN_full_adder_arch of FullAdder_179 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_178 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_178;

architecture SYN_full_adder_arch of FullAdder_178 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_177 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_177;

architecture SYN_full_adder_arch of FullAdder_177 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_176 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_176;

architecture SYN_full_adder_arch of FullAdder_176 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_175 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_175;

architecture SYN_full_adder_arch of FullAdder_175 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_174 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_174;

architecture SYN_full_adder_arch of FullAdder_174 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_173 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_173;

architecture SYN_full_adder_arch of FullAdder_173 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_172 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_172;

architecture SYN_full_adder_arch of FullAdder_172 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_171 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_171;

architecture SYN_full_adder_arch of FullAdder_171 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_170 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_170;

architecture SYN_full_adder_arch of FullAdder_170 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_169 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_169;

architecture SYN_full_adder_arch of FullAdder_169 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_168 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_168;

architecture SYN_full_adder_arch of FullAdder_168 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_167 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_167;

architecture SYN_full_adder_arch of FullAdder_167 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_166 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_166;

architecture SYN_full_adder_arch of FullAdder_166 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_165 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_165;

architecture SYN_full_adder_arch of FullAdder_165 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_164 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_164;

architecture SYN_full_adder_arch of FullAdder_164 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_163 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_163;

architecture SYN_full_adder_arch of FullAdder_163 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_162 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_162;

architecture SYN_full_adder_arch of FullAdder_162 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_161 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_161;

architecture SYN_full_adder_arch of FullAdder_161 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_160 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_160;

architecture SYN_full_adder_arch of FullAdder_160 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_159 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_159;

architecture SYN_full_adder_arch of FullAdder_159 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_158 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_158;

architecture SYN_full_adder_arch of FullAdder_158 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_157 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_157;

architecture SYN_full_adder_arch of FullAdder_157 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_156 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_156;

architecture SYN_full_adder_arch of FullAdder_156 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_155 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_155;

architecture SYN_full_adder_arch of FullAdder_155 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_154 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_154;

architecture SYN_full_adder_arch of FullAdder_154 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_153 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_153;

architecture SYN_full_adder_arch of FullAdder_153 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_152 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_152;

architecture SYN_full_adder_arch of FullAdder_152 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_151 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_151;

architecture SYN_full_adder_arch of FullAdder_151 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_150 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_150;

architecture SYN_full_adder_arch of FullAdder_150 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_149 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_149;

architecture SYN_full_adder_arch of FullAdder_149 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_148 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_148;

architecture SYN_full_adder_arch of FullAdder_148 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_147 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_147;

architecture SYN_full_adder_arch of FullAdder_147 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_146 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_146;

architecture SYN_full_adder_arch of FullAdder_146 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_145 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_145;

architecture SYN_full_adder_arch of FullAdder_145 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_144 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_144;

architecture SYN_full_adder_arch of FullAdder_144 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_143 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_143;

architecture SYN_full_adder_arch of FullAdder_143 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_142 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_142;

architecture SYN_full_adder_arch of FullAdder_142 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_141 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_141;

architecture SYN_full_adder_arch of FullAdder_141 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_140 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_140;

architecture SYN_full_adder_arch of FullAdder_140 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_139 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_139;

architecture SYN_full_adder_arch of FullAdder_139 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_138 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_138;

architecture SYN_full_adder_arch of FullAdder_138 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_137 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_137;

architecture SYN_full_adder_arch of FullAdder_137 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_136 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_136;

architecture SYN_full_adder_arch of FullAdder_136 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_135 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_135;

architecture SYN_full_adder_arch of FullAdder_135 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_134 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_134;

architecture SYN_full_adder_arch of FullAdder_134 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_133 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_133;

architecture SYN_full_adder_arch of FullAdder_133 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_132 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_132;

architecture SYN_full_adder_arch of FullAdder_132 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_131 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_131;

architecture SYN_full_adder_arch of FullAdder_131 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_130 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_130;

architecture SYN_full_adder_arch of FullAdder_130 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_129 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_129;

architecture SYN_full_adder_arch of FullAdder_129 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_128 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_128;

architecture SYN_full_adder_arch of FullAdder_128 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_127 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_127;

architecture SYN_full_adder_arch of FullAdder_127 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_126 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_126;

architecture SYN_full_adder_arch of FullAdder_126 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_125 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_125;

architecture SYN_full_adder_arch of FullAdder_125 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_124 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_124;

architecture SYN_full_adder_arch of FullAdder_124 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_123 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_123;

architecture SYN_full_adder_arch of FullAdder_123 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_122 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_122;

architecture SYN_full_adder_arch of FullAdder_122 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_121 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_121;

architecture SYN_full_adder_arch of FullAdder_121 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_120 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_120;

architecture SYN_full_adder_arch of FullAdder_120 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_119 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_119;

architecture SYN_full_adder_arch of FullAdder_119 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_118 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_118;

architecture SYN_full_adder_arch of FullAdder_118 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_117 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_117;

architecture SYN_full_adder_arch of FullAdder_117 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_116 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_116;

architecture SYN_full_adder_arch of FullAdder_116 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_115 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_115;

architecture SYN_full_adder_arch of FullAdder_115 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_114 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_114;

architecture SYN_full_adder_arch of FullAdder_114 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_113 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_113;

architecture SYN_full_adder_arch of FullAdder_113 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_112 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_112;

architecture SYN_full_adder_arch of FullAdder_112 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_111 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_111;

architecture SYN_full_adder_arch of FullAdder_111 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_110 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_110;

architecture SYN_full_adder_arch of FullAdder_110 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_109 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_109;

architecture SYN_full_adder_arch of FullAdder_109 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_108 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_108;

architecture SYN_full_adder_arch of FullAdder_108 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_107 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_107;

architecture SYN_full_adder_arch of FullAdder_107 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_106 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_106;

architecture SYN_full_adder_arch of FullAdder_106 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_105 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_105;

architecture SYN_full_adder_arch of FullAdder_105 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_104 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_104;

architecture SYN_full_adder_arch of FullAdder_104 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_103 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_103;

architecture SYN_full_adder_arch of FullAdder_103 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_102 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_102;

architecture SYN_full_adder_arch of FullAdder_102 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_101 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_101;

architecture SYN_full_adder_arch of FullAdder_101 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_100 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_100;

architecture SYN_full_adder_arch of FullAdder_100 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_99 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_99;

architecture SYN_full_adder_arch of FullAdder_99 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_98 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_98;

architecture SYN_full_adder_arch of FullAdder_98 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_97 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_97;

architecture SYN_full_adder_arch of FullAdder_97 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_96 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_96;

architecture SYN_full_adder_arch of FullAdder_96 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_95 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_95;

architecture SYN_full_adder_arch of FullAdder_95 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_94 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_94;

architecture SYN_full_adder_arch of FullAdder_94 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_93 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_93;

architecture SYN_full_adder_arch of FullAdder_93 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_92 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_92;

architecture SYN_full_adder_arch of FullAdder_92 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_91 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_91;

architecture SYN_full_adder_arch of FullAdder_91 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_90 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_90;

architecture SYN_full_adder_arch of FullAdder_90 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_89 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_89;

architecture SYN_full_adder_arch of FullAdder_89 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_88 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_88;

architecture SYN_full_adder_arch of FullAdder_88 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_87 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_87;

architecture SYN_full_adder_arch of FullAdder_87 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_86 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_86;

architecture SYN_full_adder_arch of FullAdder_86 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_85 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_85;

architecture SYN_full_adder_arch of FullAdder_85 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_84 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_84;

architecture SYN_full_adder_arch of FullAdder_84 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_83 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_83;

architecture SYN_full_adder_arch of FullAdder_83 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_82 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_82;

architecture SYN_full_adder_arch of FullAdder_82 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_81 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_81;

architecture SYN_full_adder_arch of FullAdder_81 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_80 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_80;

architecture SYN_full_adder_arch of FullAdder_80 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_79 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_79;

architecture SYN_full_adder_arch of FullAdder_79 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_78 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_78;

architecture SYN_full_adder_arch of FullAdder_78 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_77 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_77;

architecture SYN_full_adder_arch of FullAdder_77 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_76 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_76;

architecture SYN_full_adder_arch of FullAdder_76 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_75 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_75;

architecture SYN_full_adder_arch of FullAdder_75 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_74 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_74;

architecture SYN_full_adder_arch of FullAdder_74 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_73 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_73;

architecture SYN_full_adder_arch of FullAdder_73 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_72 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_72;

architecture SYN_full_adder_arch of FullAdder_72 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_71 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_71;

architecture SYN_full_adder_arch of FullAdder_71 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_70 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_70;

architecture SYN_full_adder_arch of FullAdder_70 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_69 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_69;

architecture SYN_full_adder_arch of FullAdder_69 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_68 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_68;

architecture SYN_full_adder_arch of FullAdder_68 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_67 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_67;

architecture SYN_full_adder_arch of FullAdder_67 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_66 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_66;

architecture SYN_full_adder_arch of FullAdder_66 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_65 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_65;

architecture SYN_full_adder_arch of FullAdder_65 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_64 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_64;

architecture SYN_full_adder_arch of FullAdder_64 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_63 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_63;

architecture SYN_full_adder_arch of FullAdder_63 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_62 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_62;

architecture SYN_full_adder_arch of FullAdder_62 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_61 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_61;

architecture SYN_full_adder_arch of FullAdder_61 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_60 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_60;

architecture SYN_full_adder_arch of FullAdder_60 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_59 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_59;

architecture SYN_full_adder_arch of FullAdder_59 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_58 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_58;

architecture SYN_full_adder_arch of FullAdder_58 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_57 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_57;

architecture SYN_full_adder_arch of FullAdder_57 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_56 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_56;

architecture SYN_full_adder_arch of FullAdder_56 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_55 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_55;

architecture SYN_full_adder_arch of FullAdder_55 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_54 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_54;

architecture SYN_full_adder_arch of FullAdder_54 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_53 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_53;

architecture SYN_full_adder_arch of FullAdder_53 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_52 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_52;

architecture SYN_full_adder_arch of FullAdder_52 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_51 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_51;

architecture SYN_full_adder_arch of FullAdder_51 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_50 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_50;

architecture SYN_full_adder_arch of FullAdder_50 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_49 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_49;

architecture SYN_full_adder_arch of FullAdder_49 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_48 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_48;

architecture SYN_full_adder_arch of FullAdder_48 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_47 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_47;

architecture SYN_full_adder_arch of FullAdder_47 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_46 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_46;

architecture SYN_full_adder_arch of FullAdder_46 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_45 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_45;

architecture SYN_full_adder_arch of FullAdder_45 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_44 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_44;

architecture SYN_full_adder_arch of FullAdder_44 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_43 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_43;

architecture SYN_full_adder_arch of FullAdder_43 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_42 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_42;

architecture SYN_full_adder_arch of FullAdder_42 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_41 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_41;

architecture SYN_full_adder_arch of FullAdder_41 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_40 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_40;

architecture SYN_full_adder_arch of FullAdder_40 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_39 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_39;

architecture SYN_full_adder_arch of FullAdder_39 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_38 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_38;

architecture SYN_full_adder_arch of FullAdder_38 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_37 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_37;

architecture SYN_full_adder_arch of FullAdder_37 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_36 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_36;

architecture SYN_full_adder_arch of FullAdder_36 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_35 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_35;

architecture SYN_full_adder_arch of FullAdder_35 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_34 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_34;

architecture SYN_full_adder_arch of FullAdder_34 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_33 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_33;

architecture SYN_full_adder_arch of FullAdder_33 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_32 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_32;

architecture SYN_full_adder_arch of FullAdder_32 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_31 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_31;

architecture SYN_full_adder_arch of FullAdder_31 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_30 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_30;

architecture SYN_full_adder_arch of FullAdder_30 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_29 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_29;

architecture SYN_full_adder_arch of FullAdder_29 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_28 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_28;

architecture SYN_full_adder_arch of FullAdder_28 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_27 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_27;

architecture SYN_full_adder_arch of FullAdder_27 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_26 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_26;

architecture SYN_full_adder_arch of FullAdder_26 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_25 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_25;

architecture SYN_full_adder_arch of FullAdder_25 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_24 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_24;

architecture SYN_full_adder_arch of FullAdder_24 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_23 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_23;

architecture SYN_full_adder_arch of FullAdder_23 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_22 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_22;

architecture SYN_full_adder_arch of FullAdder_22 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_21 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_21;

architecture SYN_full_adder_arch of FullAdder_21 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_20 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_20;

architecture SYN_full_adder_arch of FullAdder_20 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_19 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_19;

architecture SYN_full_adder_arch of FullAdder_19 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_18 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_18;

architecture SYN_full_adder_arch of FullAdder_18 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_17 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_17;

architecture SYN_full_adder_arch of FullAdder_17 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_16 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_16;

architecture SYN_full_adder_arch of FullAdder_16 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_15 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_15;

architecture SYN_full_adder_arch of FullAdder_15 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_14 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_14;

architecture SYN_full_adder_arch of FullAdder_14 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_13 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_13;

architecture SYN_full_adder_arch of FullAdder_13 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_12 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_12;

architecture SYN_full_adder_arch of FullAdder_12 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_11 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_11;

architecture SYN_full_adder_arch of FullAdder_11 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_10 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_10;

architecture SYN_full_adder_arch of FullAdder_10 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_9 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_9;

architecture SYN_full_adder_arch of FullAdder_9 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_8 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_8;

architecture SYN_full_adder_arch of FullAdder_8 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_7 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_7;

architecture SYN_full_adder_arch of FullAdder_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_6 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_6;

architecture SYN_full_adder_arch of FullAdder_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_5 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_5;

architecture SYN_full_adder_arch of FullAdder_5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_4 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_4;

architecture SYN_full_adder_arch of FullAdder_4 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_3 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_3;

architecture SYN_full_adder_arch of FullAdder_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_2 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_2;

architecture SYN_full_adder_arch of FullAdder_2 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_1 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_1;

architecture SYN_full_adder_arch of FullAdder_1 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n5, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n5);
   U1 : INV_X1 port map( A => n4, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n5, B2 => ci, ZN => n4);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_83 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_83;

architecture SYN_mux_arch of Mux_DATA_SIZE4_83 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => dout(0));
   U2 : INV_X1 port map( A => n5, ZN => dout(3));
   U3 : INV_X1 port map( A => n2, ZN => dout(1));
   U4 : INV_X1 port map( A => n3, ZN => dout(2));
   U5 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U6 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U7 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U8 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_82 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_82;

architecture SYN_mux_arch of Mux_DATA_SIZE4_82 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => dout(2));
   U2 : INV_X1 port map( A => n2, ZN => dout(1));
   U3 : INV_X1 port map( A => n1, ZN => dout(0));
   U4 : INV_X1 port map( A => n5, ZN => dout(3));
   U5 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U7 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U8 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_81 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_81;

architecture SYN_mux_arch of Mux_DATA_SIZE4_81 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => dout(2));
   U2 : INV_X1 port map( A => n2, ZN => dout(1));
   U3 : INV_X1 port map( A => n1, ZN => dout(0));
   U4 : INV_X1 port map( A => n5, ZN => dout(3));
   U5 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U7 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U8 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_80 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_80;

architecture SYN_mux_arch of Mux_DATA_SIZE4_80 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => dout(3));
   U2 : INV_X1 port map( A => n3, ZN => dout(2));
   U3 : INV_X1 port map( A => n2, ZN => dout(1));
   U4 : INV_X1 port map( A => n1, ZN => dout(0));
   U5 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U7 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U8 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_79 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_79;

architecture SYN_mux_arch of Mux_DATA_SIZE4_79 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => dout(3));
   U2 : INV_X1 port map( A => n1, ZN => dout(0));
   U3 : INV_X1 port map( A => n2, ZN => dout(1));
   U4 : INV_X1 port map( A => n3, ZN => dout(2));
   U5 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U6 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U7 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U8 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_78 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_78;

architecture SYN_mux_arch of Mux_DATA_SIZE4_78 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => dout(3));
   U2 : INV_X1 port map( A => n2, ZN => dout(1));
   U3 : INV_X1 port map( A => n1, ZN => dout(0));
   U4 : INV_X1 port map( A => n3, ZN => dout(2));
   U5 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U7 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U8 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_77 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_77;

architecture SYN_mux_arch of Mux_DATA_SIZE4_77 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n7 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => sel, Z => n1);
   U2 : INV_X1 port map( A => sel, ZN => n2);
   U3 : INV_X1 port map( A => n5, ZN => dout(2));
   U4 : INV_X1 port map( A => n7, ZN => dout(3));
   U5 : INV_X1 port map( A => n3, ZN => dout(0));
   U6 : AOI22_X1 port map( A1 => n2, A2 => din0(1), B1 => n1, B2 => din1(1), ZN
                           => n4);
   U7 : AOI22_X1 port map( A1 => n2, A2 => din0(2), B1 => n1, B2 => din1(2), ZN
                           => n5);
   U8 : AOI22_X1 port map( A1 => n2, A2 => din0(0), B1 => n1, B2 => din1(0), ZN
                           => n3);
   U9 : AOI22_X1 port map( A1 => din0(3), A2 => n2, B1 => n1, B2 => din1(3), ZN
                           => n7);
   U10 : INV_X1 port map( A => n4, ZN => dout(1));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_76 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_76;

architecture SYN_mux_arch of Mux_DATA_SIZE4_76 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => dout(3));
   U2 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U3 : INV_X1 port map( A => n3, ZN => dout(2));
   U4 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U5 : INV_X1 port map( A => n2, ZN => dout(1));
   U6 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U7 : INV_X1 port map( A => n1, ZN => dout(0));
   U8 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_75 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_75;

architecture SYN_mux_arch of Mux_DATA_SIZE4_75 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => dout(3));
   U2 : INV_X1 port map( A => n3, ZN => dout(2));
   U3 : INV_X1 port map( A => n2, ZN => dout(1));
   U4 : INV_X1 port map( A => n1, ZN => dout(0));
   U5 : INV_X1 port map( A => sel, ZN => n4);
   U6 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U7 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U8 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U9 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_74 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_74;

architecture SYN_mux_arch of Mux_DATA_SIZE4_74 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => dout(1));
   U2 : INV_X1 port map( A => n1, ZN => dout(0));
   U3 : INV_X1 port map( A => n3, ZN => dout(2));
   U4 : INV_X1 port map( A => n5, ZN => dout(3));
   U5 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U7 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U8 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_73 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_73;

architecture SYN_mux_arch of Mux_DATA_SIZE4_73 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => dout(0));
   U2 : INV_X1 port map( A => n5, ZN => dout(3));
   U3 : INV_X1 port map( A => n3, ZN => dout(2));
   U4 : INV_X1 port map( A => n2, ZN => dout(1));
   U5 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U6 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U7 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U8 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_72 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_72;

architecture SYN_mux_arch of Mux_DATA_SIZE4_72 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => sel, Z => n1);
   U2 : INV_X1 port map( A => n4, ZN => dout(2));
   U3 : INV_X1 port map( A => n3, ZN => dout(1));
   U4 : INV_X1 port map( A => n2, ZN => dout(0));
   U5 : INV_X1 port map( A => n7, ZN => dout(3));
   U6 : AOI22_X1 port map( A1 => din0(3), A2 => n5, B1 => n1, B2 => din1(3), ZN
                           => n7);
   U7 : AOI22_X1 port map( A1 => din0(2), A2 => n5, B1 => din1(2), B2 => n1, ZN
                           => n4);
   U8 : AOI22_X1 port map( A1 => din0(0), A2 => n5, B1 => din1(0), B2 => n1, ZN
                           => n2);
   U9 : AOI22_X1 port map( A1 => din0(1), A2 => n5, B1 => din1(1), B2 => sel, 
                           ZN => n3);
   U10 : INV_X1 port map( A => sel, ZN => n5);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_71 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_71;

architecture SYN_mux_arch of Mux_DATA_SIZE4_71 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => dout(1));
   U2 : INV_X1 port map( A => n1, ZN => dout(0));
   U3 : INV_X1 port map( A => n3, ZN => dout(2));
   U4 : INV_X1 port map( A => n5, ZN => dout(3));
   U5 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U7 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U8 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_70 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_70;

architecture SYN_mux_arch of Mux_DATA_SIZE4_70 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n8, n9 : std_logic;

begin
   
   U1 : INV_X1 port map( A => din1(0), ZN => n3);
   U2 : INV_X1 port map( A => din0(0), ZN => n2);
   U3 : OAI22_X1 port map( A1 => n2, A2 => sel, B1 => n3, B2 => n8, ZN => 
                           dout(0));
   U4 : INV_X1 port map( A => n4, ZN => dout(1));
   U5 : INV_X1 port map( A => n5, ZN => dout(2));
   U6 : INV_X1 port map( A => n9, ZN => dout(3));
   U7 : AOI22_X1 port map( A1 => din0(3), A2 => n8, B1 => sel, B2 => din1(3), 
                           ZN => n9);
   U8 : AOI22_X1 port map( A1 => din0(2), A2 => n8, B1 => din1(2), B2 => sel, 
                           ZN => n5);
   U9 : AOI22_X1 port map( A1 => din0(1), A2 => n8, B1 => din1(1), B2 => sel, 
                           ZN => n4);
   U10 : INV_X1 port map( A => sel, ZN => n8);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_69 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_69;

architecture SYN_mux_arch of Mux_DATA_SIZE4_69 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n3, n4, n5, n10, n11, n12, n13, n14, n15 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => sel, Z => n5);
   U2 : INV_X1 port map( A => din1(0), ZN => n4);
   U3 : INV_X1 port map( A => din0(0), ZN => n3);
   U4 : CLKBUF_X1 port map( A => n14, Z => n1);
   U5 : OAI22_X1 port map( A1 => n5, A2 => n3, B1 => n14, B2 => n4, ZN => 
                           dout(0));
   U6 : INV_X1 port map( A => n15, ZN => dout(3));
   U7 : CLKBUF_X1 port map( A => n1, Z => n10);
   U8 : INV_X1 port map( A => n13, ZN => dout(2));
   U9 : INV_X1 port map( A => n12, ZN => dout(1));
   U10 : INV_X1 port map( A => n10, ZN => n11);
   U11 : AOI22_X1 port map( A1 => din0(3), A2 => n10, B1 => n11, B2 => din1(3),
                           ZN => n15);
   U12 : AOI22_X1 port map( A1 => n1, A2 => din0(1), B1 => n5, B2 => din1(1), 
                           ZN => n12);
   U13 : AOI22_X1 port map( A1 => n1, A2 => din0(2), B1 => n5, B2 => din1(2), 
                           ZN => n13);
   U14 : INV_X1 port map( A => sel, ZN => n14);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_68 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_68;

architecture SYN_mux_arch of Mux_DATA_SIZE4_68 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => dout(3));
   U2 : INV_X1 port map( A => n4, ZN => dout(2));
   U3 : INV_X1 port map( A => n3, ZN => dout(1));
   U4 : INV_X1 port map( A => n2, ZN => dout(0));
   U5 : AOI22_X1 port map( A1 => din0(2), A2 => n1, B1 => din1(2), B2 => sel, 
                           ZN => n4);
   U6 : AOI22_X1 port map( A1 => din0(3), A2 => n1, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U7 : AOI22_X1 port map( A1 => din0(0), A2 => n1, B1 => din1(0), B2 => sel, 
                           ZN => n2);
   U8 : AOI22_X1 port map( A1 => din0(1), A2 => n1, B1 => din1(1), B2 => sel, 
                           ZN => n3);
   U9 : INV_X1 port map( A => sel, ZN => n1);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_67 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_67;

architecture SYN_mux_arch of Mux_DATA_SIZE4_67 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => dout(3));
   U2 : INV_X1 port map( A => n3, ZN => dout(2));
   U3 : INV_X1 port map( A => n2, ZN => dout(1));
   U4 : INV_X1 port map( A => n1, ZN => dout(0));
   U5 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U6 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U7 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U8 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_66 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_66;

architecture SYN_mux_arch of Mux_DATA_SIZE4_66 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => dout(3));
   U2 : INV_X1 port map( A => n3, ZN => dout(2));
   U3 : INV_X1 port map( A => n2, ZN => dout(1));
   U4 : INV_X1 port map( A => n1, ZN => dout(0));
   U5 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U6 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U7 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U8 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_65 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_65;

architecture SYN_mux_arch of Mux_DATA_SIZE4_65 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => dout(3));
   U2 : INV_X1 port map( A => n3, ZN => dout(2));
   U3 : INV_X1 port map( A => n2, ZN => dout(1));
   U4 : INV_X1 port map( A => n1, ZN => dout(0));
   U5 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U7 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U8 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_64 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_64;

architecture SYN_mux_arch of Mux_DATA_SIZE4_64 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => dout(3));
   U2 : INV_X1 port map( A => n2, ZN => dout(1));
   U3 : INV_X1 port map( A => n3, ZN => dout(2));
   U4 : INV_X1 port map( A => n1, ZN => dout(0));
   U5 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U7 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U8 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_63 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_63;

architecture SYN_mux_arch of Mux_DATA_SIZE4_63 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => dout(3));
   U2 : INV_X1 port map( A => n3, ZN => dout(2));
   U3 : INV_X1 port map( A => n2, ZN => dout(1));
   U4 : INV_X1 port map( A => n1, ZN => dout(0));
   U5 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U6 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U7 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U8 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_62 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_62;

architecture SYN_mux_arch of Mux_DATA_SIZE4_62 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => dout(3));
   U2 : INV_X1 port map( A => n3, ZN => dout(2));
   U3 : INV_X1 port map( A => n2, ZN => dout(1));
   U4 : INV_X1 port map( A => n1, ZN => dout(0));
   U5 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U6 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U7 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U8 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_61 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_61;

architecture SYN_mux_arch of Mux_DATA_SIZE4_61 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n8, n11, n12, n13, n14 : std_logic;

begin
   
   U1 : INV_X1 port map( A => din1(3), ZN => n11);
   U2 : INV_X1 port map( A => din1(2), ZN => n3);
   U3 : INV_X1 port map( A => din0(3), ZN => n8);
   U4 : INV_X1 port map( A => din0(2), ZN => n2);
   U5 : OAI22_X1 port map( A1 => sel, A2 => n8, B1 => n5, B2 => n11, ZN => 
                           dout(3));
   U6 : CLKBUF_X1 port map( A => sel, Z => n4);
   U7 : OAI22_X1 port map( A1 => n2, A2 => n4, B1 => n14, B2 => n3, ZN => 
                           dout(2));
   U8 : INV_X1 port map( A => sel, ZN => n5);
   U9 : INV_X1 port map( A => n12, ZN => dout(0));
   U10 : INV_X1 port map( A => n13, ZN => dout(1));
   U11 : AOI22_X1 port map( A1 => din0(0), A2 => n14, B1 => n4, B2 => din1(0), 
                           ZN => n12);
   U12 : AOI22_X1 port map( A1 => n14, A2 => din0(1), B1 => din1(1), B2 => sel,
                           ZN => n13);
   U13 : INV_X1 port map( A => sel, ZN => n14);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_60 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_60;

architecture SYN_mux_arch of Mux_DATA_SIZE4_60 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => dout(0));
   U2 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U3 : INV_X1 port map( A => n2, ZN => dout(1));
   U4 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U5 : INV_X1 port map( A => n3, ZN => dout(2));
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U7 : INV_X1 port map( A => n5, ZN => dout(3));
   U8 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_59 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_59;

architecture SYN_mux_arch of Mux_DATA_SIZE4_59 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => sel, ZN => n4);
   U2 : INV_X1 port map( A => n1, ZN => dout(0));
   U3 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U4 : INV_X1 port map( A => n2, ZN => dout(1));
   U5 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U6 : INV_X1 port map( A => n3, ZN => dout(2));
   U7 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U8 : INV_X1 port map( A => n5, ZN => dout(3));
   U9 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_58 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_58;

architecture SYN_mux_arch of Mux_DATA_SIZE4_58 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => sel, ZN => n4);
   U2 : INV_X1 port map( A => n1, ZN => dout(0));
   U3 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U4 : INV_X1 port map( A => n2, ZN => dout(1));
   U5 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U6 : INV_X1 port map( A => n3, ZN => dout(2));
   U7 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U8 : INV_X1 port map( A => n5, ZN => dout(3));
   U9 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_57 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_57;

architecture SYN_mux_arch of Mux_DATA_SIZE4_57 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => sel, ZN => n4);
   U2 : INV_X1 port map( A => n5, ZN => dout(3));
   U3 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U4 : INV_X1 port map( A => n1, ZN => dout(0));
   U5 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U6 : INV_X1 port map( A => n2, ZN => dout(1));
   U7 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U8 : INV_X1 port map( A => n3, ZN => dout(2));
   U9 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_56 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_56;

architecture SYN_mux_arch of Mux_DATA_SIZE4_56 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => dout(1));
   U2 : INV_X1 port map( A => n3, ZN => dout(2));
   U3 : INV_X1 port map( A => n5, ZN => dout(3));
   U4 : INV_X1 port map( A => n1, ZN => dout(0));
   U5 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U6 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U7 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U8 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_55 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_55;

architecture SYN_mux_arch of Mux_DATA_SIZE4_55 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U2 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U3 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U4 : INV_X1 port map( A => sel, ZN => n4);
   U5 : INV_X1 port map( A => n3, ZN => dout(2));
   U6 : INV_X1 port map( A => n5, ZN => dout(3));
   U7 : INV_X1 port map( A => n1, ZN => dout(0));
   U8 : INV_X1 port map( A => n2, ZN => dout(1));
   U9 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_54 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_54;

architecture SYN_mux_arch of Mux_DATA_SIZE4_54 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U2 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U3 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U4 : INV_X1 port map( A => sel, ZN => n4);
   U5 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U6 : INV_X1 port map( A => n1, ZN => dout(0));
   U7 : INV_X1 port map( A => n2, ZN => dout(1));
   U8 : INV_X1 port map( A => n3, ZN => dout(2));
   U9 : INV_X1 port map( A => n5, ZN => dout(3));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_53 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_53;

architecture SYN_mux_arch of Mux_DATA_SIZE4_53 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => sel, ZN => n4);
   U2 : INV_X1 port map( A => n5, ZN => dout(3));
   U3 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U4 : INV_X1 port map( A => n2, ZN => dout(1));
   U5 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U6 : INV_X1 port map( A => n3, ZN => dout(2));
   U7 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U8 : INV_X1 port map( A => n1, ZN => dout(0));
   U9 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_52 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_52;

architecture SYN_mux_arch of Mux_DATA_SIZE4_52 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => sel, ZN => n4);
   U2 : INV_X1 port map( A => n5, ZN => dout(3));
   U3 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U4 : INV_X1 port map( A => n2, ZN => dout(1));
   U5 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U6 : INV_X1 port map( A => n3, ZN => dout(2));
   U7 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U8 : INV_X1 port map( A => n1, ZN => dout(0));
   U9 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_51 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_51;

architecture SYN_mux_arch of Mux_DATA_SIZE4_51 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => sel, ZN => n4);
   U2 : INV_X1 port map( A => n2, ZN => dout(1));
   U3 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U4 : INV_X1 port map( A => n3, ZN => dout(2));
   U5 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U6 : INV_X1 port map( A => n5, ZN => dout(3));
   U7 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U8 : INV_X1 port map( A => n1, ZN => dout(0));
   U9 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_50 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_50;

architecture SYN_mux_arch of Mux_DATA_SIZE4_50 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => sel, ZN => n4);
   U2 : INV_X1 port map( A => n5, ZN => dout(3));
   U3 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U4 : INV_X1 port map( A => n2, ZN => dout(1));
   U5 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U6 : INV_X1 port map( A => n3, ZN => dout(2));
   U7 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U8 : INV_X1 port map( A => n1, ZN => dout(0));
   U9 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_49 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_49;

architecture SYN_mux_arch of Mux_DATA_SIZE4_49 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n4, n5, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : INV_X1 port map( A => sel, ZN => n1);
   U2 : INV_X1 port map( A => din1(1), ZN => n5);
   U3 : INV_X1 port map( A => din0(1), ZN => n4);
   U4 : CLKBUF_X1 port map( A => sel, Z => n2);
   U5 : OAI22_X1 port map( A1 => n4, A2 => n2, B1 => n5, B2 => n1, ZN => 
                           dout(1));
   U6 : INV_X1 port map( A => n12, ZN => dout(3));
   U7 : AOI22_X1 port map( A1 => din0(3), A2 => n1, B1 => sel, B2 => din1(3), 
                           ZN => n12);
   U8 : INV_X1 port map( A => n9, ZN => dout(0));
   U9 : AOI22_X1 port map( A1 => din0(0), A2 => n11, B1 => sel, B2 => din1(0), 
                           ZN => n9);
   U10 : AOI22_X1 port map( A1 => din0(2), A2 => n11, B1 => sel, B2 => din1(2),
                           ZN => n10);
   U11 : INV_X1 port map( A => sel, ZN => n11);
   U12 : INV_X1 port map( A => n10, ZN => dout(2));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_48 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_48;

architecture SYN_mux_arch of Mux_DATA_SIZE4_48 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => dout(3));
   U2 : AOI22_X1 port map( A1 => din0(3), A2 => n1, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U3 : INV_X1 port map( A => n4, ZN => dout(2));
   U4 : AOI22_X1 port map( A1 => din0(2), A2 => n1, B1 => din1(2), B2 => sel, 
                           ZN => n4);
   U5 : INV_X1 port map( A => n3, ZN => dout(1));
   U6 : AOI22_X1 port map( A1 => din0(1), A2 => n1, B1 => din1(1), B2 => sel, 
                           ZN => n3);
   U7 : INV_X1 port map( A => n2, ZN => dout(0));
   U8 : AOI22_X1 port map( A1 => din0(0), A2 => n1, B1 => din1(0), B2 => sel, 
                           ZN => n2);
   U9 : INV_X1 port map( A => sel, ZN => n1);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_47 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_47;

architecture SYN_mux_arch of Mux_DATA_SIZE4_47 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => dout(3));
   U2 : INV_X1 port map( A => n3, ZN => dout(2));
   U3 : INV_X1 port map( A => n2, ZN => dout(1));
   U4 : INV_X1 port map( A => n1, ZN => dout(0));
   U5 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U7 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U8 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_46 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_46;

architecture SYN_mux_arch of Mux_DATA_SIZE4_46 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => dout(3));
   U2 : INV_X1 port map( A => n3, ZN => dout(2));
   U3 : INV_X1 port map( A => n2, ZN => dout(1));
   U4 : INV_X1 port map( A => n1, ZN => dout(0));
   U5 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U7 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U8 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_45 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_45;

architecture SYN_mux_arch of Mux_DATA_SIZE4_45 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => dout(3));
   U2 : INV_X1 port map( A => n3, ZN => dout(2));
   U3 : INV_X1 port map( A => n2, ZN => dout(1));
   U4 : INV_X1 port map( A => n1, ZN => dout(0));
   U5 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U6 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U7 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U8 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_44 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_44;

architecture SYN_mux_arch of Mux_DATA_SIZE4_44 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => dout(3));
   U2 : INV_X1 port map( A => n3, ZN => dout(2));
   U3 : INV_X1 port map( A => n2, ZN => dout(1));
   U4 : INV_X1 port map( A => n1, ZN => dout(0));
   U5 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U7 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U8 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_43 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_43;

architecture SYN_mux_arch of Mux_DATA_SIZE4_43 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => dout(3));
   U2 : INV_X1 port map( A => n3, ZN => dout(2));
   U3 : INV_X1 port map( A => n2, ZN => dout(1));
   U4 : INV_X1 port map( A => n1, ZN => dout(0));
   U5 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U7 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U8 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_42 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_42;

architecture SYN_mux_arch of Mux_DATA_SIZE4_42 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => dout(3));
   U2 : INV_X1 port map( A => n3, ZN => dout(2));
   U3 : INV_X1 port map( A => n2, ZN => dout(1));
   U4 : INV_X1 port map( A => n1, ZN => dout(0));
   U5 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U7 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U8 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_41 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_41;

architecture SYN_mux_arch of Mux_DATA_SIZE4_41 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3, n5, n6, n7, n9, n10, n11, n13, n14 : std_logic;

begin
   
   U1 : INV_X1 port map( A => din1(3), ZN => n3);
   U2 : INV_X1 port map( A => din1(2), ZN => n14);
   U3 : INV_X1 port map( A => din1(1), ZN => n10);
   U4 : INV_X1 port map( A => din1(0), ZN => n6);
   U5 : INV_X1 port map( A => din0(3), ZN => n2);
   U6 : INV_X1 port map( A => din0(2), ZN => n13);
   U7 : INV_X1 port map( A => din0(1), ZN => n9);
   U8 : INV_X1 port map( A => din0(0), ZN => n5);
   U9 : BUF_X1 port map( A => sel, Z => n11);
   U10 : OAI22_X1 port map( A1 => n11, A2 => n2, B1 => n7, B2 => n3, ZN => 
                           dout(3));
   U11 : OAI22_X1 port map( A1 => n11, A2 => n5, B1 => n7, B2 => n6, ZN => 
                           dout(0));
   U12 : INV_X1 port map( A => sel, ZN => n7);
   U13 : OAI22_X1 port map( A1 => n11, A2 => n9, B1 => n7, B2 => n10, ZN => 
                           dout(1));
   U14 : OAI22_X1 port map( A1 => n13, A2 => n11, B1 => n7, B2 => n14, ZN => 
                           dout(2));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_40 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_40;

architecture SYN_mux_arch of Mux_DATA_SIZE4_40 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => dout(1));
   U2 : AOI22_X1 port map( A1 => din0(1), A2 => n1, B1 => din1(1), B2 => sel, 
                           ZN => n3);
   U3 : INV_X1 port map( A => n5, ZN => dout(3));
   U4 : AOI22_X1 port map( A1 => din0(3), A2 => n1, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U5 : INV_X1 port map( A => n4, ZN => dout(2));
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n1, B1 => din1(2), B2 => sel, 
                           ZN => n4);
   U7 : INV_X1 port map( A => n2, ZN => dout(0));
   U8 : AOI22_X1 port map( A1 => din0(0), A2 => n1, B1 => din1(0), B2 => sel, 
                           ZN => n2);
   U9 : INV_X1 port map( A => sel, ZN => n1);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_39 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_39;

architecture SYN_mux_arch of Mux_DATA_SIZE4_39 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => dout(3));
   U2 : INV_X1 port map( A => n3, ZN => dout(2));
   U3 : INV_X1 port map( A => n2, ZN => dout(1));
   U4 : INV_X1 port map( A => n1, ZN => dout(0));
   U5 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U7 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U8 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_38 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_38;

architecture SYN_mux_arch of Mux_DATA_SIZE4_38 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => dout(3));
   U2 : INV_X1 port map( A => n3, ZN => dout(2));
   U3 : INV_X1 port map( A => n2, ZN => dout(1));
   U4 : INV_X1 port map( A => n1, ZN => dout(0));
   U5 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U7 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U8 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_37 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_37;

architecture SYN_mux_arch of Mux_DATA_SIZE4_37 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => dout(3));
   U2 : INV_X1 port map( A => n3, ZN => dout(2));
   U3 : INV_X1 port map( A => n2, ZN => dout(1));
   U4 : INV_X1 port map( A => n1, ZN => dout(0));
   U5 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U7 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U8 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_36 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_36;

architecture SYN_mux_arch of Mux_DATA_SIZE4_36 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => dout(3));
   U2 : INV_X1 port map( A => n3, ZN => dout(2));
   U3 : INV_X1 port map( A => n2, ZN => dout(1));
   U4 : INV_X1 port map( A => n1, ZN => dout(0));
   U5 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U7 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U8 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_35 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_35;

architecture SYN_mux_arch of Mux_DATA_SIZE4_35 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => sel, ZN => n4);
   U2 : INV_X1 port map( A => n5, ZN => dout(3));
   U3 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U4 : INV_X1 port map( A => n3, ZN => dout(2));
   U5 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U6 : INV_X1 port map( A => n2, ZN => dout(1));
   U7 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U8 : INV_X1 port map( A => n1, ZN => dout(0));
   U9 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_34 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_34;

architecture SYN_mux_arch of Mux_DATA_SIZE4_34 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => dout(2));
   U2 : INV_X1 port map( A => n2, ZN => dout(1));
   U3 : INV_X1 port map( A => n1, ZN => dout(0));
   U4 : INV_X1 port map( A => n5, ZN => dout(3));
   U5 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U7 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U8 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_33 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_33;

architecture SYN_mux_arch of Mux_DATA_SIZE4_33 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n3, n4, n6, n7, n9, n10, n11, n13, n14 : std_logic;

begin
   
   U1 : INV_X1 port map( A => din0(3), ZN => n13);
   U2 : INV_X1 port map( A => din0(2), ZN => n9);
   U3 : INV_X1 port map( A => din1(0), ZN => n4);
   U4 : INV_X1 port map( A => din0(1), ZN => n6);
   U5 : INV_X1 port map( A => din1(1), ZN => n7);
   U6 : INV_X1 port map( A => din0(0), ZN => n3);
   U7 : INV_X1 port map( A => din1(2), ZN => n10);
   U8 : INV_X1 port map( A => din1(3), ZN => n14);
   U9 : BUF_X1 port map( A => sel, Z => n11);
   U10 : INV_X1 port map( A => sel, ZN => n1);
   U11 : OAI22_X1 port map( A1 => n11, A2 => n3, B1 => n1, B2 => n4, ZN => 
                           dout(0));
   U12 : OAI22_X1 port map( A1 => n6, A2 => n11, B1 => n7, B2 => n1, ZN => 
                           dout(1));
   U13 : OAI22_X1 port map( A1 => n9, A2 => n11, B1 => n1, B2 => n10, ZN => 
                           dout(2));
   U14 : OAI22_X1 port map( A1 => n13, A2 => n11, B1 => n14, B2 => n1, ZN => 
                           dout(3));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_32 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_32;

architecture SYN_mux_arch of Mux_DATA_SIZE4_32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n2, ZN => dout(0));
   U2 : AOI22_X1 port map( A1 => din0(0), A2 => n1, B1 => din1(0), B2 => sel, 
                           ZN => n2);
   U3 : INV_X1 port map( A => n3, ZN => dout(1));
   U4 : AOI22_X1 port map( A1 => din0(1), A2 => n1, B1 => din1(1), B2 => sel, 
                           ZN => n3);
   U5 : INV_X1 port map( A => n4, ZN => dout(2));
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n1, B1 => din1(2), B2 => sel, 
                           ZN => n4);
   U7 : INV_X1 port map( A => n5, ZN => dout(3));
   U8 : AOI22_X1 port map( A1 => din0(3), A2 => n1, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U9 : INV_X1 port map( A => sel, ZN => n1);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_31 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_31;

architecture SYN_mux_arch of Mux_DATA_SIZE4_31 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => sel, ZN => n4);
   U2 : INV_X1 port map( A => n5, ZN => dout(3));
   U3 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U4 : INV_X1 port map( A => n2, ZN => dout(1));
   U5 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U6 : INV_X1 port map( A => n1, ZN => dout(0));
   U7 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U8 : INV_X1 port map( A => n3, ZN => dout(2));
   U9 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_30 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_30;

architecture SYN_mux_arch of Mux_DATA_SIZE4_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => dout(3));
   U2 : INV_X1 port map( A => n1, ZN => dout(0));
   U3 : INV_X1 port map( A => n2, ZN => dout(1));
   U4 : INV_X1 port map( A => n3, ZN => dout(2));
   U5 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U6 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U7 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U8 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_29 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_29;

architecture SYN_mux_arch of Mux_DATA_SIZE4_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => dout(0));
   U2 : INV_X1 port map( A => n2, ZN => dout(1));
   U3 : INV_X1 port map( A => n3, ZN => dout(2));
   U4 : INV_X1 port map( A => n5, ZN => dout(3));
   U5 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U6 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U7 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U8 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_28 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_28;

architecture SYN_mux_arch of Mux_DATA_SIZE4_28 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => sel, ZN => n4);
   U2 : INV_X1 port map( A => n1, ZN => dout(0));
   U3 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U4 : INV_X1 port map( A => n2, ZN => dout(1));
   U5 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U6 : INV_X1 port map( A => n3, ZN => dout(2));
   U7 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U8 : INV_X1 port map( A => n5, ZN => dout(3));
   U9 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_27 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_27;

architecture SYN_mux_arch of Mux_DATA_SIZE4_27 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => sel, ZN => n4);
   U2 : INV_X1 port map( A => n1, ZN => dout(0));
   U3 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U4 : INV_X1 port map( A => n2, ZN => dout(1));
   U5 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U6 : INV_X1 port map( A => n3, ZN => dout(2));
   U7 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U8 : INV_X1 port map( A => n5, ZN => dout(3));
   U9 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_26 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_26;

architecture SYN_mux_arch of Mux_DATA_SIZE4_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => dout(0));
   U2 : INV_X1 port map( A => n2, ZN => dout(1));
   U3 : INV_X1 port map( A => n3, ZN => dout(2));
   U4 : INV_X1 port map( A => n5, ZN => dout(3));
   U5 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U7 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U8 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_25 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_25;

architecture SYN_mux_arch of Mux_DATA_SIZE4_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => dout(0));
   U2 : INV_X1 port map( A => n2, ZN => dout(1));
   U3 : INV_X1 port map( A => n3, ZN => dout(2));
   U4 : INV_X1 port map( A => n5, ZN => dout(3));
   U5 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U7 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U8 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_24 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_24;

architecture SYN_mux_arch of Mux_DATA_SIZE4_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => dout(0));
   U2 : INV_X1 port map( A => n2, ZN => dout(1));
   U3 : INV_X1 port map( A => n3, ZN => dout(2));
   U4 : INV_X1 port map( A => n5, ZN => dout(3));
   U5 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U7 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U8 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_23 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_23;

architecture SYN_mux_arch of Mux_DATA_SIZE4_23 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => sel, ZN => n4);
   U2 : INV_X1 port map( A => n1, ZN => dout(0));
   U3 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U4 : INV_X1 port map( A => n2, ZN => dout(1));
   U5 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U6 : INV_X1 port map( A => n3, ZN => dout(2));
   U7 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U8 : INV_X1 port map( A => n5, ZN => dout(3));
   U9 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_22 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_22;

architecture SYN_mux_arch of Mux_DATA_SIZE4_22 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => sel, ZN => n4);
   U2 : INV_X1 port map( A => n1, ZN => dout(0));
   U3 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U4 : INV_X1 port map( A => n2, ZN => dout(1));
   U5 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U6 : INV_X1 port map( A => n3, ZN => dout(2));
   U7 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U8 : INV_X1 port map( A => n5, ZN => dout(3));
   U9 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_21 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_21;

architecture SYN_mux_arch of Mux_DATA_SIZE4_21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => dout(0));
   U2 : INV_X1 port map( A => n2, ZN => dout(1));
   U3 : INV_X1 port map( A => n3, ZN => dout(2));
   U4 : INV_X1 port map( A => n5, ZN => dout(3));
   U5 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U7 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U8 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_20 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_20;

architecture SYN_mux_arch of Mux_DATA_SIZE4_20 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));
   U2 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U3 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U4 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_19 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_19;

architecture SYN_mux_arch of Mux_DATA_SIZE4_19 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));
   U2 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U3 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U4 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_18 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_18;

architecture SYN_mux_arch of Mux_DATA_SIZE4_18 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));
   U2 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U3 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U4 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_17 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_17;

architecture SYN_mux_arch of Mux_DATA_SIZE4_17 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));
   U2 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U3 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U4 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_16 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_16;

architecture SYN_mux_arch of Mux_DATA_SIZE4_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n5, ZN => dout(3));
   U2 : AOI22_X1 port map( A1 => din0(3), A2 => n1, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U3 : INV_X1 port map( A => n3, ZN => dout(1));
   U4 : AOI22_X1 port map( A1 => din0(1), A2 => n1, B1 => din1(1), B2 => sel, 
                           ZN => n3);
   U5 : INV_X1 port map( A => n4, ZN => dout(2));
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n1, B1 => din1(2), B2 => sel, 
                           ZN => n4);
   U7 : INV_X1 port map( A => n2, ZN => dout(0));
   U8 : AOI22_X1 port map( A1 => din0(0), A2 => n1, B1 => din1(0), B2 => sel, 
                           ZN => n2);
   U9 : INV_X1 port map( A => sel, ZN => n1);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_15 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_15;

architecture SYN_mux_arch of Mux_DATA_SIZE4_15 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => sel, ZN => n4);
   U2 : INV_X1 port map( A => n5, ZN => dout(3));
   U3 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U4 : INV_X1 port map( A => n2, ZN => dout(1));
   U5 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U6 : INV_X1 port map( A => n3, ZN => dout(2));
   U7 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U8 : INV_X1 port map( A => n1, ZN => dout(0));
   U9 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_14 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_14;

architecture SYN_mux_arch of Mux_DATA_SIZE4_14 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => sel, ZN => n4);
   U2 : INV_X1 port map( A => n5, ZN => dout(3));
   U3 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U4 : INV_X1 port map( A => n2, ZN => dout(1));
   U5 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U6 : INV_X1 port map( A => n3, ZN => dout(2));
   U7 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U8 : INV_X1 port map( A => n1, ZN => dout(0));
   U9 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_13 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_13;

architecture SYN_mux_arch of Mux_DATA_SIZE4_13 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => sel, ZN => n4);
   U2 : INV_X1 port map( A => n5, ZN => dout(3));
   U3 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U4 : INV_X1 port map( A => n2, ZN => dout(1));
   U5 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U6 : INV_X1 port map( A => n3, ZN => dout(2));
   U7 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U8 : INV_X1 port map( A => n1, ZN => dout(0));
   U9 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_12 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_12;

architecture SYN_mux_arch of Mux_DATA_SIZE4_12 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => sel, ZN => n4);
   U2 : INV_X1 port map( A => n5, ZN => dout(3));
   U3 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U4 : INV_X1 port map( A => n2, ZN => dout(1));
   U5 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U6 : INV_X1 port map( A => n3, ZN => dout(2));
   U7 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U8 : INV_X1 port map( A => n1, ZN => dout(0));
   U9 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_11 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_11;

architecture SYN_mux_arch of Mux_DATA_SIZE4_11 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => sel, ZN => n4);
   U2 : INV_X1 port map( A => n2, ZN => dout(1));
   U3 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U4 : INV_X1 port map( A => n3, ZN => dout(2));
   U5 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U6 : INV_X1 port map( A => n5, ZN => dout(3));
   U7 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U8 : INV_X1 port map( A => n1, ZN => dout(0));
   U9 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_10 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_10;

architecture SYN_mux_arch of Mux_DATA_SIZE4_10 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => sel, ZN => n4);
   U2 : INV_X1 port map( A => n5, ZN => dout(3));
   U3 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U4 : INV_X1 port map( A => n2, ZN => dout(1));
   U5 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U6 : INV_X1 port map( A => n3, ZN => dout(2));
   U7 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U8 : INV_X1 port map( A => n1, ZN => dout(0));
   U9 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_9 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_9;

architecture SYN_mux_arch of Mux_DATA_SIZE4_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n3, n4, n6, n8, n10, n11, n13, n14, n15 : std_logic;

begin
   
   U1 : INV_X1 port map( A => din0(0), ZN => n10);
   U2 : INV_X1 port map( A => din0(1), ZN => n3);
   U3 : INV_X1 port map( A => din0(2), ZN => n6);
   U4 : INV_X1 port map( A => din0(3), ZN => n13);
   U5 : INV_X1 port map( A => din1(0), ZN => n11);
   U6 : INV_X1 port map( A => din1(1), ZN => n4);
   U7 : INV_X1 port map( A => din1(2), ZN => n8);
   U8 : INV_X1 port map( A => din1(3), ZN => n14);
   U9 : BUF_X1 port map( A => sel, Z => n1);
   U10 : OAI22_X1 port map( A1 => n3, A2 => n1, B1 => n15, B2 => n4, ZN => 
                           dout(1));
   U11 : OAI22_X1 port map( A1 => n6, A2 => n1, B1 => n15, B2 => n8, ZN => 
                           dout(2));
   U12 : OAI22_X1 port map( A1 => n10, A2 => n1, B1 => n15, B2 => n11, ZN => 
                           dout(0));
   U13 : OAI22_X1 port map( A1 => n13, A2 => n1, B1 => n15, B2 => n14, ZN => 
                           dout(3));
   U14 : INV_X1 port map( A => sel, ZN => n15);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_8 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_8;

architecture SYN_mux_arch of Mux_DATA_SIZE4_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n3, ZN => dout(1));
   U2 : AOI22_X1 port map( A1 => din0(1), A2 => n1, B1 => din1(1), B2 => sel, 
                           ZN => n3);
   U3 : INV_X1 port map( A => n2, ZN => dout(0));
   U4 : AOI22_X1 port map( A1 => din0(0), A2 => n1, B1 => din1(0), B2 => sel, 
                           ZN => n2);
   U5 : INV_X1 port map( A => n5, ZN => dout(3));
   U6 : AOI22_X1 port map( A1 => din0(3), A2 => n1, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U7 : INV_X1 port map( A => n4, ZN => dout(2));
   U8 : AOI22_X1 port map( A1 => din0(2), A2 => n1, B1 => din1(2), B2 => sel, 
                           ZN => n4);
   U9 : INV_X1 port map( A => sel, ZN => n1);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_7 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_7;

architecture SYN_mux_arch of Mux_DATA_SIZE4_7 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => sel, ZN => n4);
   U2 : INV_X1 port map( A => n5, ZN => dout(3));
   U3 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U4 : INV_X1 port map( A => n1, ZN => dout(0));
   U5 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U6 : INV_X1 port map( A => n2, ZN => dout(1));
   U7 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U8 : INV_X1 port map( A => n3, ZN => dout(2));
   U9 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_6 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_6;

architecture SYN_mux_arch of Mux_DATA_SIZE4_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => dout(0));
   U2 : INV_X1 port map( A => n2, ZN => dout(1));
   U3 : INV_X1 port map( A => n3, ZN => dout(2));
   U4 : INV_X1 port map( A => n5, ZN => dout(3));
   U5 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U6 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U7 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U8 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_5 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_5;

architecture SYN_mux_arch of Mux_DATA_SIZE4_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => dout(0));
   U2 : INV_X1 port map( A => n2, ZN => dout(1));
   U3 : INV_X1 port map( A => n3, ZN => dout(2));
   U4 : INV_X1 port map( A => n5, ZN => dout(3));
   U5 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U6 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U7 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U8 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_4 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_4;

architecture SYN_mux_arch of Mux_DATA_SIZE4_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => dout(0));
   U2 : INV_X1 port map( A => n2, ZN => dout(1));
   U3 : INV_X1 port map( A => n5, ZN => dout(3));
   U4 : INV_X1 port map( A => n3, ZN => dout(2));
   U5 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U6 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U7 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U8 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_3 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_3;

architecture SYN_mux_arch of Mux_DATA_SIZE4_3 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => sel, ZN => n4);
   U2 : INV_X1 port map( A => n1, ZN => dout(0));
   U3 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U4 : INV_X1 port map( A => n2, ZN => dout(1));
   U5 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U6 : INV_X1 port map( A => n3, ZN => dout(2));
   U7 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U8 : INV_X1 port map( A => n5, ZN => dout(3));
   U9 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_2 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_2;

architecture SYN_mux_arch of Mux_DATA_SIZE4_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n1, ZN => dout(0));
   U2 : INV_X1 port map( A => n2, ZN => dout(1));
   U3 : INV_X1 port map( A => n5, ZN => dout(3));
   U4 : INV_X1 port map( A => n3, ZN => dout(2));
   U5 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => sel, B2 => din1(3), 
                           ZN => n5);
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => sel, 
                           ZN => n3);
   U7 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => sel, 
                           ZN => n2);
   U8 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => sel, 
                           ZN => n1);
   U9 : INV_X1 port map( A => sel, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_1 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_1;

architecture SYN_mux_arch of Mux_DATA_SIZE4_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n3, n4, n6, n8, n10, n11, n13, n14, n15 : std_logic;

begin
   
   U1 : INV_X1 port map( A => din0(0), ZN => n3);
   U2 : INV_X1 port map( A => din0(1), ZN => n10);
   U3 : INV_X1 port map( A => din0(2), ZN => n13);
   U4 : INV_X1 port map( A => din0(3), ZN => n6);
   U5 : INV_X1 port map( A => din1(0), ZN => n4);
   U6 : INV_X1 port map( A => din1(1), ZN => n11);
   U7 : INV_X1 port map( A => din1(2), ZN => n14);
   U8 : INV_X1 port map( A => din1(3), ZN => n8);
   U9 : BUF_X1 port map( A => sel, Z => n1);
   U10 : OAI22_X1 port map( A1 => n3, A2 => n1, B1 => n15, B2 => n4, ZN => 
                           dout(0));
   U11 : OAI22_X1 port map( A1 => n6, A2 => n1, B1 => n15, B2 => n8, ZN => 
                           dout(3));
   U12 : OAI22_X1 port map( A1 => n10, A2 => n1, B1 => n11, B2 => n15, ZN => 
                           dout(1));
   U13 : OAI22_X1 port map( A1 => n13, A2 => n1, B1 => n14, B2 => n15, ZN => 
                           dout(2));
   U14 : INV_X1 port map( A => sel, ZN => n15);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_167 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_167;

architecture SYN_rca_arch of Rca_DATA_SIZE4_167 is

   component FullAdder_665
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_666
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_667
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_668
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_668 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_667 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_666 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_665 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_166 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_166;

architecture SYN_rca_arch of Rca_DATA_SIZE4_166 is

   component FullAdder_661
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_662
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_663
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_664
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_664 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_663 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_662 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_661 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_165 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_165;

architecture SYN_rca_arch of Rca_DATA_SIZE4_165 is

   component FullAdder_657
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_658
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_659
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_660
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_660 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_659 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_658 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_657 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_164 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_164;

architecture SYN_rca_arch of Rca_DATA_SIZE4_164 is

   component FullAdder_653
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_654
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_655
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_656
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_656 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_655 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_654 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_653 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_163 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_163;

architecture SYN_rca_arch of Rca_DATA_SIZE4_163 is

   component FullAdder_649
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_650
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_651
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_652
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_652 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_651 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_650 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_649 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_162 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_162;

architecture SYN_rca_arch of Rca_DATA_SIZE4_162 is

   component FullAdder_645
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_646
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_647
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_648
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_648 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_647 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_646 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_645 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_161 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_161;

architecture SYN_rca_arch of Rca_DATA_SIZE4_161 is

   component FullAdder_641
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_642
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_643
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_644
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_644 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_643 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_642 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_641 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_160 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_160;

architecture SYN_rca_arch of Rca_DATA_SIZE4_160 is

   component FullAdder_637
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_638
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_639
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_640
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_640 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_639 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_638 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_637 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_159 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_159;

architecture SYN_rca_arch of Rca_DATA_SIZE4_159 is

   component FullAdder_633
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_634
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_635
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_636
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_636 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_635 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_634 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_633 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_158 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_158;

architecture SYN_rca_arch of Rca_DATA_SIZE4_158 is

   component FullAdder_629
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_630
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_631
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_632
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_632 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_631 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_630 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_629 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_157 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_157;

architecture SYN_rca_arch of Rca_DATA_SIZE4_157 is

   component FullAdder_625
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_626
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_627
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_628
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_628 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_627 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_626 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_625 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_156 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_156;

architecture SYN_rca_arch of Rca_DATA_SIZE4_156 is

   component FullAdder_621
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_622
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_623
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_624
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_624 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_623 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_622 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_621 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_155 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_155;

architecture SYN_rca_arch of Rca_DATA_SIZE4_155 is

   component FullAdder_617
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_618
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_619
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_620
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_620 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_619 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_618 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_617 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_154 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_154;

architecture SYN_rca_arch of Rca_DATA_SIZE4_154 is

   component FullAdder_613
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_614
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_615
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_616
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_616 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_615 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_614 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_613 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_153 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_153;

architecture SYN_rca_arch of Rca_DATA_SIZE4_153 is

   component FullAdder_609
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_610
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_611
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_612
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_612 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_611 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_610 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_609 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_152 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_152;

architecture SYN_rca_arch of Rca_DATA_SIZE4_152 is

   component FullAdder_605
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_606
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_607
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_608
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_608 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_607 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_606 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_605 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_151 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_151;

architecture SYN_rca_arch of Rca_DATA_SIZE4_151 is

   component FullAdder_601
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_602
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_603
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_604
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_604 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_603 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_602 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_601 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_150 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_150;

architecture SYN_rca_arch of Rca_DATA_SIZE4_150 is

   component FullAdder_597
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_598
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_599
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_600
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_600 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_599 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_598 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_597 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_149 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_149;

architecture SYN_rca_arch of Rca_DATA_SIZE4_149 is

   component FullAdder_593
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_594
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_595
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_596
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_596 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_595 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_594 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_593 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_148 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_148;

architecture SYN_rca_arch of Rca_DATA_SIZE4_148 is

   component FullAdder_589
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_590
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_591
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_592
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_592 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_591 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_590 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_589 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_147 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_147;

architecture SYN_rca_arch of Rca_DATA_SIZE4_147 is

   component FullAdder_585
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_586
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_587
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_588
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_588 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_587 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_586 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_585 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_146 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_146;

architecture SYN_rca_arch of Rca_DATA_SIZE4_146 is

   component FullAdder_581
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_582
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_583
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_584
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_584 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_583 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_582 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_581 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_145 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_145;

architecture SYN_rca_arch of Rca_DATA_SIZE4_145 is

   component FullAdder_577
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_578
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_579
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_580
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_580 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_579 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_578 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_577 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_144 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_144;

architecture SYN_rca_arch of Rca_DATA_SIZE4_144 is

   component FullAdder_573
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_574
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_575
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_576
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_576 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_575 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_574 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_573 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_143 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_143;

architecture SYN_rca_arch of Rca_DATA_SIZE4_143 is

   component FullAdder_569
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_570
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_571
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_572
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_572 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_571 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_570 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_569 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_142 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_142;

architecture SYN_rca_arch of Rca_DATA_SIZE4_142 is

   component FullAdder_565
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_566
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_567
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_568
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_568 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_567 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_566 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_565 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_141 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_141;

architecture SYN_rca_arch of Rca_DATA_SIZE4_141 is

   component FullAdder_561
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_562
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_563
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_564
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_564 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_563 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_562 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_561 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_140 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_140;

architecture SYN_rca_arch of Rca_DATA_SIZE4_140 is

   component FullAdder_557
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_558
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_559
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_560
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_560 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_559 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_558 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_557 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_139 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_139;

architecture SYN_rca_arch of Rca_DATA_SIZE4_139 is

   component FullAdder_553
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_554
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_555
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_556
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_556 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_555 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_554 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_553 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_138 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_138;

architecture SYN_rca_arch of Rca_DATA_SIZE4_138 is

   component FullAdder_549
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_550
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_551
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_552
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_552 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_551 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_550 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_549 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_137 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_137;

architecture SYN_rca_arch of Rca_DATA_SIZE4_137 is

   component FullAdder_545
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_546
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_547
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_548
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_548 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_547 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_546 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_545 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_136 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_136;

architecture SYN_rca_arch of Rca_DATA_SIZE4_136 is

   component FullAdder_541
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_542
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_543
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_544
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_544 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_543 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_542 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_541 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_135 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_135;

architecture SYN_rca_arch of Rca_DATA_SIZE4_135 is

   component FullAdder_537
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_538
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_539
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_540
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_540 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_539 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_538 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_537 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_134 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_134;

architecture SYN_rca_arch of Rca_DATA_SIZE4_134 is

   component FullAdder_533
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_534
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_535
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_536
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_536 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_535 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_534 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_533 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_133 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_133;

architecture SYN_rca_arch of Rca_DATA_SIZE4_133 is

   component FullAdder_529
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_530
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_531
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_532
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_532 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_531 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_530 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_529 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_132 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_132;

architecture SYN_rca_arch of Rca_DATA_SIZE4_132 is

   component FullAdder_525
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_526
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_527
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_528
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_528 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_527 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_526 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_525 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_131 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_131;

architecture SYN_rca_arch of Rca_DATA_SIZE4_131 is

   component FullAdder_521
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_522
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_523
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_524
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_524 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_523 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_522 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_521 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_130 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_130;

architecture SYN_rca_arch of Rca_DATA_SIZE4_130 is

   component FullAdder_517
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_518
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_519
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_520
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_520 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_519 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_518 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_517 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_129 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_129;

architecture SYN_rca_arch of Rca_DATA_SIZE4_129 is

   component FullAdder_513
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_514
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_515
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_516
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_516 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_515 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_514 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_513 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_128 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_128;

architecture SYN_rca_arch of Rca_DATA_SIZE4_128 is

   component FullAdder_509
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_510
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_511
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_512
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_512 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_511 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_510 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_509 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_127 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_127;

architecture SYN_rca_arch of Rca_DATA_SIZE4_127 is

   component FullAdder_505
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_506
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_507
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_508
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_508 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_507 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_506 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_505 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_126 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_126;

architecture SYN_rca_arch of Rca_DATA_SIZE4_126 is

   component FullAdder_501
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_502
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_503
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_504
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_504 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_503 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_502 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_501 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_125 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_125;

architecture SYN_rca_arch of Rca_DATA_SIZE4_125 is

   component FullAdder_497
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_498
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_499
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_500
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_500 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_499 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_498 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_497 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_124 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_124;

architecture SYN_rca_arch of Rca_DATA_SIZE4_124 is

   component FullAdder_493
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_494
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_495
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_496
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_496 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_495 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_494 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_493 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_123 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_123;

architecture SYN_rca_arch of Rca_DATA_SIZE4_123 is

   component FullAdder_489
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_490
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_491
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_492
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_492 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_491 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_490 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_489 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_122 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_122;

architecture SYN_rca_arch of Rca_DATA_SIZE4_122 is

   component FullAdder_485
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_486
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_487
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_488
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_488 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_487 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_486 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_485 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_121 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_121;

architecture SYN_rca_arch of Rca_DATA_SIZE4_121 is

   component FullAdder_481
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_482
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_483
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_484
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_484 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_483 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_482 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_481 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_120 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_120;

architecture SYN_rca_arch of Rca_DATA_SIZE4_120 is

   component FullAdder_477
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_478
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_479
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_480
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_480 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_479 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_478 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_477 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_119 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_119;

architecture SYN_rca_arch of Rca_DATA_SIZE4_119 is

   component FullAdder_473
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_474
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_475
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_476
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_476 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_475 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_474 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_473 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_118 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_118;

architecture SYN_rca_arch of Rca_DATA_SIZE4_118 is

   component FullAdder_469
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_470
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_471
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_472
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_472 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_471 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_470 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_469 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_117 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_117;

architecture SYN_rca_arch of Rca_DATA_SIZE4_117 is

   component FullAdder_465
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_466
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_467
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_468
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_468 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_467 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_466 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_465 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_116 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_116;

architecture SYN_rca_arch of Rca_DATA_SIZE4_116 is

   component FullAdder_461
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_462
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_463
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_464
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_464 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_463 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_462 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_461 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_115 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_115;

architecture SYN_rca_arch of Rca_DATA_SIZE4_115 is

   component FullAdder_457
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_458
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_459
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_460
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_460 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_459 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_458 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_457 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_114 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_114;

architecture SYN_rca_arch of Rca_DATA_SIZE4_114 is

   component FullAdder_453
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_454
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_455
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_456
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_456 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_455 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_454 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_453 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_113 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_113;

architecture SYN_rca_arch of Rca_DATA_SIZE4_113 is

   component FullAdder_449
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_450
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_451
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_452
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_452 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_451 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_450 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_449 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_112 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_112;

architecture SYN_rca_arch of Rca_DATA_SIZE4_112 is

   component FullAdder_445
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_446
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_447
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_448
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_448 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_447 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_446 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_445 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_111 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_111;

architecture SYN_rca_arch of Rca_DATA_SIZE4_111 is

   component FullAdder_441
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_442
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_443
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_444
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_444 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_443 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_442 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_441 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_110 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_110;

architecture SYN_rca_arch of Rca_DATA_SIZE4_110 is

   component FullAdder_437
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_438
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_439
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_440
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_440 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_439 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_438 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_437 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_109 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_109;

architecture SYN_rca_arch of Rca_DATA_SIZE4_109 is

   component FullAdder_433
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_434
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_435
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_436
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_436 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_435 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_434 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_433 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_108 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_108;

architecture SYN_rca_arch of Rca_DATA_SIZE4_108 is

   component FullAdder_429
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_430
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_431
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_432
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_432 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_431 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_430 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_429 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_107 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_107;

architecture SYN_rca_arch of Rca_DATA_SIZE4_107 is

   component FullAdder_425
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_426
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_427
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_428
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_428 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_427 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_426 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_425 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_106 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_106;

architecture SYN_rca_arch of Rca_DATA_SIZE4_106 is

   component FullAdder_421
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_422
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_423
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_424
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_424 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_423 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_422 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_421 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_105 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_105;

architecture SYN_rca_arch of Rca_DATA_SIZE4_105 is

   component FullAdder_417
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_418
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_419
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_420
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_420 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_419 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_418 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_417 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_104 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_104;

architecture SYN_rca_arch of Rca_DATA_SIZE4_104 is

   component FullAdder_413
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_414
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_415
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_416
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_416 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_415 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_414 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_413 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_103 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_103;

architecture SYN_rca_arch of Rca_DATA_SIZE4_103 is

   component FullAdder_409
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_410
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_411
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_412
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_412 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_411 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_410 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_409 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_102 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_102;

architecture SYN_rca_arch of Rca_DATA_SIZE4_102 is

   component FullAdder_405
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_406
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_407
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_408
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_408 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_407 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_406 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_405 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_101 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_101;

architecture SYN_rca_arch of Rca_DATA_SIZE4_101 is

   component FullAdder_401
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_402
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_403
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_404
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_404 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_403 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_402 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_401 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_100 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_100;

architecture SYN_rca_arch of Rca_DATA_SIZE4_100 is

   component FullAdder_397
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_398
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_399
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_400
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_400 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_399 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_398 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_397 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_99 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_99;

architecture SYN_rca_arch of Rca_DATA_SIZE4_99 is

   component FullAdder_393
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_394
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_395
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_396
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_396 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_395 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_394 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_393 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_98 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_98;

architecture SYN_rca_arch of Rca_DATA_SIZE4_98 is

   component FullAdder_389
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_390
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_391
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_392
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_392 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_391 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_390 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_389 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_97 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_97;

architecture SYN_rca_arch of Rca_DATA_SIZE4_97 is

   component FullAdder_385
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_386
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_387
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_388
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_388 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_387 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_386 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_385 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_96 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_96;

architecture SYN_rca_arch of Rca_DATA_SIZE4_96 is

   component FullAdder_381
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_382
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_383
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_384
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_384 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_383 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_382 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_381 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_95 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_95;

architecture SYN_rca_arch of Rca_DATA_SIZE4_95 is

   component FullAdder_377
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_378
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_379
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_380
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_380 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_379 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_378 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_377 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_94 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_94;

architecture SYN_rca_arch of Rca_DATA_SIZE4_94 is

   component FullAdder_373
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_374
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_375
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_376
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_376 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_375 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_374 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_373 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_93 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_93;

architecture SYN_rca_arch of Rca_DATA_SIZE4_93 is

   component FullAdder_369
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_370
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_371
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_372
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_372 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_371 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_370 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_369 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_92 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_92;

architecture SYN_rca_arch of Rca_DATA_SIZE4_92 is

   component FullAdder_365
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_366
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_367
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_368
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_368 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_367 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_366 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_365 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_91 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_91;

architecture SYN_rca_arch of Rca_DATA_SIZE4_91 is

   component FullAdder_361
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_362
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_363
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_364
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_364 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_363 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_362 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_361 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_90 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_90;

architecture SYN_rca_arch of Rca_DATA_SIZE4_90 is

   component FullAdder_357
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_358
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_359
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_360
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_360 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_359 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_358 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_357 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_89 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_89;

architecture SYN_rca_arch of Rca_DATA_SIZE4_89 is

   component FullAdder_353
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_354
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_355
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_356
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_356 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_355 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_354 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_353 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_88 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_88;

architecture SYN_rca_arch of Rca_DATA_SIZE4_88 is

   component FullAdder_349
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_350
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_351
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_352
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_352 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_351 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_350 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_349 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_87 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_87;

architecture SYN_rca_arch of Rca_DATA_SIZE4_87 is

   component FullAdder_345
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_346
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_347
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_348
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_348 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_347 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_346 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_345 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_86 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_86;

architecture SYN_rca_arch of Rca_DATA_SIZE4_86 is

   component FullAdder_341
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_342
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_343
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_344
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_344 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_343 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_342 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_341 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_85 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_85;

architecture SYN_rca_arch of Rca_DATA_SIZE4_85 is

   component FullAdder_337
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_338
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_339
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_340
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_340 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_339 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_338 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_337 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_84 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_84;

architecture SYN_rca_arch of Rca_DATA_SIZE4_84 is

   component FullAdder_333
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_334
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_335
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_336
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_336 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_335 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_334 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_333 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_83 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_83;

architecture SYN_rca_arch of Rca_DATA_SIZE4_83 is

   component FullAdder_329
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_330
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_331
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_332
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_332 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_331 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_330 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_329 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_82 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_82;

architecture SYN_rca_arch of Rca_DATA_SIZE4_82 is

   component FullAdder_325
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_326
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_327
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_328
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_328 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_327 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_326 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_325 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_81 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_81;

architecture SYN_rca_arch of Rca_DATA_SIZE4_81 is

   component FullAdder_321
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_322
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_323
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_324
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_324 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_323 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_322 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_321 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_80 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_80;

architecture SYN_rca_arch of Rca_DATA_SIZE4_80 is

   component FullAdder_317
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_318
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_319
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_320
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_320 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_319 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_318 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_317 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_79 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_79;

architecture SYN_rca_arch of Rca_DATA_SIZE4_79 is

   component FullAdder_313
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_314
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_315
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_316
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_316 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_315 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_314 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_313 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_78 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_78;

architecture SYN_rca_arch of Rca_DATA_SIZE4_78 is

   component FullAdder_309
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_310
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_311
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_312
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_312 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_311 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_310 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_309 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_77 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_77;

architecture SYN_rca_arch of Rca_DATA_SIZE4_77 is

   component FullAdder_305
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_306
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_307
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_308
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_308 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_307 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_306 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_305 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_76 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_76;

architecture SYN_rca_arch of Rca_DATA_SIZE4_76 is

   component FullAdder_301
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_302
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_303
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_304
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_304 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_303 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_302 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_301 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_75 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_75;

architecture SYN_rca_arch of Rca_DATA_SIZE4_75 is

   component FullAdder_297
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_298
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_299
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_300
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_300 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_299 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_298 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_297 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_74 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_74;

architecture SYN_rca_arch of Rca_DATA_SIZE4_74 is

   component FullAdder_293
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_294
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_295
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_296
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_296 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_295 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_294 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_293 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_73 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_73;

architecture SYN_rca_arch of Rca_DATA_SIZE4_73 is

   component FullAdder_289
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_290
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_291
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_292
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_292 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_291 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_290 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_289 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_72 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_72;

architecture SYN_rca_arch of Rca_DATA_SIZE4_72 is

   component FullAdder_285
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_286
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_287
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_288
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_288 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_287 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_286 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_285 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_71 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_71;

architecture SYN_rca_arch of Rca_DATA_SIZE4_71 is

   component FullAdder_281
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_282
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_283
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_284
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_284 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_283 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_282 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_281 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_70 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_70;

architecture SYN_rca_arch of Rca_DATA_SIZE4_70 is

   component FullAdder_277
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_278
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_279
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_280
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_280 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_279 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_278 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_277 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_69 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_69;

architecture SYN_rca_arch of Rca_DATA_SIZE4_69 is

   component FullAdder_273
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_274
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_275
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_276
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_276 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_275 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_274 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_273 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_68 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_68;

architecture SYN_rca_arch of Rca_DATA_SIZE4_68 is

   component FullAdder_269
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_270
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_271
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_272
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_272 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_271 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_270 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_269 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_67 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_67;

architecture SYN_rca_arch of Rca_DATA_SIZE4_67 is

   component FullAdder_265
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_266
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_267
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_268
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_268 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_267 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_266 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_265 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_66 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_66;

architecture SYN_rca_arch of Rca_DATA_SIZE4_66 is

   component FullAdder_261
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_262
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_263
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_264
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_264 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_263 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_262 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_261 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_65 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_65;

architecture SYN_rca_arch of Rca_DATA_SIZE4_65 is

   component FullAdder_257
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_258
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_259
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_260
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_260 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_259 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_258 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_257 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_64 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_64;

architecture SYN_rca_arch of Rca_DATA_SIZE4_64 is

   component FullAdder_253
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_254
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_255
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_256
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_256 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_255 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_254 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_253 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_63 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_63;

architecture SYN_rca_arch of Rca_DATA_SIZE4_63 is

   component FullAdder_249
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_250
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_251
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_252
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_252 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_251 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_250 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_249 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_62 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_62;

architecture SYN_rca_arch of Rca_DATA_SIZE4_62 is

   component FullAdder_245
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_246
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_247
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_248
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_248 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_247 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_246 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_245 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_61 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_61;

architecture SYN_rca_arch of Rca_DATA_SIZE4_61 is

   component FullAdder_241
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_242
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_243
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_244
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_244 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_243 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_242 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_241 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_60 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_60;

architecture SYN_rca_arch of Rca_DATA_SIZE4_60 is

   component FullAdder_237
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_238
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_239
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_240
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_240 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_239 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_238 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_237 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_59 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_59;

architecture SYN_rca_arch of Rca_DATA_SIZE4_59 is

   component FullAdder_233
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_234
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_235
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_236
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_236 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_235 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_234 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_233 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_58 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_58;

architecture SYN_rca_arch of Rca_DATA_SIZE4_58 is

   component FullAdder_229
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_230
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_231
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_232
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_232 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_231 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_230 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_229 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_57 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_57;

architecture SYN_rca_arch of Rca_DATA_SIZE4_57 is

   component FullAdder_225
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_226
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_227
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_228
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_228 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_227 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_226 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_225 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_56 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_56;

architecture SYN_rca_arch of Rca_DATA_SIZE4_56 is

   component FullAdder_221
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_222
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_223
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_224
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_224 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_223 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_222 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_221 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_55 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_55;

architecture SYN_rca_arch of Rca_DATA_SIZE4_55 is

   component FullAdder_217
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_218
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_219
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_220
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_220 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_219 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_218 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_217 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_54 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_54;

architecture SYN_rca_arch of Rca_DATA_SIZE4_54 is

   component FullAdder_213
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_214
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_215
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_216
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_216 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_215 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_214 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_213 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_53 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_53;

architecture SYN_rca_arch of Rca_DATA_SIZE4_53 is

   component FullAdder_209
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_210
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_211
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_212
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_212 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_211 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_210 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_209 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_52 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_52;

architecture SYN_rca_arch of Rca_DATA_SIZE4_52 is

   component FullAdder_205
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_206
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_207
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_208
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_208 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_207 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_206 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_205 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_51 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_51;

architecture SYN_rca_arch of Rca_DATA_SIZE4_51 is

   component FullAdder_201
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_202
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_203
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_204
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_204 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_203 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_202 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_201 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_50 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_50;

architecture SYN_rca_arch of Rca_DATA_SIZE4_50 is

   component FullAdder_197
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_198
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_199
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_200
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_200 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_199 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_198 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_197 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_49 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_49;

architecture SYN_rca_arch of Rca_DATA_SIZE4_49 is

   component FullAdder_193
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_194
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_195
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_196
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_196 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_195 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_194 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_193 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_48 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_48;

architecture SYN_rca_arch of Rca_DATA_SIZE4_48 is

   component FullAdder_189
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_190
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_191
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_192
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_192 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_191 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_190 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_189 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_47 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_47;

architecture SYN_rca_arch of Rca_DATA_SIZE4_47 is

   component FullAdder_185
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_186
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_187
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_188
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_188 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_187 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_186 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_185 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_46 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_46;

architecture SYN_rca_arch of Rca_DATA_SIZE4_46 is

   component FullAdder_181
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_182
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_183
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_184
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_184 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_183 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_182 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_181 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_45 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_45;

architecture SYN_rca_arch of Rca_DATA_SIZE4_45 is

   component FullAdder_177
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_178
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_179
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_180
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_180 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_179 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_178 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_177 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_44 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_44;

architecture SYN_rca_arch of Rca_DATA_SIZE4_44 is

   component FullAdder_173
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_174
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_175
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_176
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_176 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_175 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_174 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_173 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_43 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_43;

architecture SYN_rca_arch of Rca_DATA_SIZE4_43 is

   component FullAdder_169
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_170
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_171
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_172
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_172 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_171 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_170 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_169 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_42 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_42;

architecture SYN_rca_arch of Rca_DATA_SIZE4_42 is

   component FullAdder_165
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_166
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_167
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_168
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_168 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_167 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_166 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_165 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_41 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_41;

architecture SYN_rca_arch of Rca_DATA_SIZE4_41 is

   component FullAdder_161
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_162
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_163
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_164
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_164 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_163 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_162 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_161 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_40 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_40;

architecture SYN_rca_arch of Rca_DATA_SIZE4_40 is

   component FullAdder_157
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_158
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_159
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_160
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_160 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_159 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_158 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_157 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_39 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_39;

architecture SYN_rca_arch of Rca_DATA_SIZE4_39 is

   component FullAdder_153
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_154
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_155
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_156
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_156 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_155 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_154 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_153 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_38 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_38;

architecture SYN_rca_arch of Rca_DATA_SIZE4_38 is

   component FullAdder_149
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_150
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_151
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_152
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_152 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_151 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_150 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_149 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_37 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_37;

architecture SYN_rca_arch of Rca_DATA_SIZE4_37 is

   component FullAdder_145
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_146
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_147
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_148
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_148 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_147 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_146 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_145 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_36 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_36;

architecture SYN_rca_arch of Rca_DATA_SIZE4_36 is

   component FullAdder_141
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_142
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_143
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_144
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_144 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_143 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_142 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_141 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_35 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_35;

architecture SYN_rca_arch of Rca_DATA_SIZE4_35 is

   component FullAdder_137
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_138
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_139
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_140
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_140 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_139 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_138 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_137 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_34 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_34;

architecture SYN_rca_arch of Rca_DATA_SIZE4_34 is

   component FullAdder_133
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_134
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_135
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_136
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_136 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_135 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_134 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_133 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_33 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_33;

architecture SYN_rca_arch of Rca_DATA_SIZE4_33 is

   component FullAdder_129
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_130
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_131
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_132
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_132 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_131 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_130 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_129 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_32 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_32;

architecture SYN_rca_arch of Rca_DATA_SIZE4_32 is

   component FullAdder_125
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_126
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_127
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_128
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_128 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_127 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_126 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_125 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_31 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_31;

architecture SYN_rca_arch of Rca_DATA_SIZE4_31 is

   component FullAdder_121
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_122
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_123
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_124
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_124 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_123 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_122 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_121 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_30 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_30;

architecture SYN_rca_arch of Rca_DATA_SIZE4_30 is

   component FullAdder_117
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_118
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_119
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_120
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_120 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_119 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_118 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_117 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_29 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_29;

architecture SYN_rca_arch of Rca_DATA_SIZE4_29 is

   component FullAdder_113
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_114
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_115
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_116
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_116 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_115 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_114 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_113 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_28 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_28;

architecture SYN_rca_arch of Rca_DATA_SIZE4_28 is

   component FullAdder_109
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_110
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_111
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_112
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_112 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_111 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_110 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_109 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_27 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_27;

architecture SYN_rca_arch of Rca_DATA_SIZE4_27 is

   component FullAdder_105
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_106
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_107
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_108
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_108 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_107 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_106 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_105 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_26 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_26;

architecture SYN_rca_arch of Rca_DATA_SIZE4_26 is

   component FullAdder_101
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_102
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_103
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_104
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_104 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_103 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_102 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_101 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_25 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_25;

architecture SYN_rca_arch of Rca_DATA_SIZE4_25 is

   component FullAdder_97
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_98
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_99
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_100
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_100 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_99 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_98 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_97 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_24 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_24;

architecture SYN_rca_arch of Rca_DATA_SIZE4_24 is

   component FullAdder_93
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_94
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_95
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_96
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_96 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_95 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_94 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_93 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_23 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_23;

architecture SYN_rca_arch of Rca_DATA_SIZE4_23 is

   component FullAdder_89
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_90
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_91
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_92
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_92 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_91 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_90 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_89 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_22 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_22;

architecture SYN_rca_arch of Rca_DATA_SIZE4_22 is

   component FullAdder_85
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_86
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_87
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_88
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_88 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_87 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_86 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_85 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_21 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_21;

architecture SYN_rca_arch of Rca_DATA_SIZE4_21 is

   component FullAdder_81
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_82
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_83
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_84
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_84 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_83 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_82 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_81 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_20 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_20;

architecture SYN_rca_arch of Rca_DATA_SIZE4_20 is

   component FullAdder_77
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_78
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_79
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_80
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_80 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_79 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_78 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_77 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_19 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_19;

architecture SYN_rca_arch of Rca_DATA_SIZE4_19 is

   component FullAdder_73
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_74
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_75
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_76
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_76 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_75 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_74 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_73 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_18 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_18;

architecture SYN_rca_arch of Rca_DATA_SIZE4_18 is

   component FullAdder_69
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_70
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_71
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_72
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_72 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_71 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_70 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_69 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_17 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_17;

architecture SYN_rca_arch of Rca_DATA_SIZE4_17 is

   component FullAdder_65
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_66
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_67
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_68
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_68 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_67 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_66 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_65 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_16 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_16;

architecture SYN_rca_arch of Rca_DATA_SIZE4_16 is

   component FullAdder_61
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_62
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_63
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_64
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_64 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_63 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_62 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_61 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_15 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_15;

architecture SYN_rca_arch of Rca_DATA_SIZE4_15 is

   component FullAdder_57
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_58
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_59
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_60
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_60 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_59 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_58 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_57 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_14 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_14;

architecture SYN_rca_arch of Rca_DATA_SIZE4_14 is

   component FullAdder_53
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_54
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_55
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_56
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_56 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_55 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_54 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_53 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_13 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_13;

architecture SYN_rca_arch of Rca_DATA_SIZE4_13 is

   component FullAdder_49
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_50
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_51
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_52
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_52 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_51 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_50 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_49 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_12 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_12;

architecture SYN_rca_arch of Rca_DATA_SIZE4_12 is

   component FullAdder_45
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_46
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_47
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_48
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_48 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_47 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_46 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_45 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_11 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_11;

architecture SYN_rca_arch of Rca_DATA_SIZE4_11 is

   component FullAdder_41
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_42
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_43
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_44
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_44 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_43 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_42 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_41 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_10 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_10;

architecture SYN_rca_arch of Rca_DATA_SIZE4_10 is

   component FullAdder_37
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_38
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_39
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_40
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_40 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_39 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_38 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_37 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_9 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_9;

architecture SYN_rca_arch of Rca_DATA_SIZE4_9 is

   component FullAdder_33
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_34
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_35
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_36
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_36 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_35 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_34 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_33 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_8 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_8;

architecture SYN_rca_arch of Rca_DATA_SIZE4_8 is

   component FullAdder_29
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_30
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_31
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_32
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_32 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_31 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_30 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_29 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_7 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_7;

architecture SYN_rca_arch of Rca_DATA_SIZE4_7 is

   component FullAdder_25
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_26
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_27
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_28
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_28 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_27 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_26 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_25 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_6 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_6;

architecture SYN_rca_arch of Rca_DATA_SIZE4_6 is

   component FullAdder_21
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_22
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_23
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_24
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_24 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_23 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_22 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_21 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_5 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_5;

architecture SYN_rca_arch of Rca_DATA_SIZE4_5 is

   component FullAdder_17
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_18
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_19
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_20
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_20 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_19 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_18 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_17 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_4 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_4;

architecture SYN_rca_arch of Rca_DATA_SIZE4_4 is

   component FullAdder_13
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_14
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_15
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_16
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_16 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_15 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_14 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_13 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_3 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_3;

architecture SYN_rca_arch of Rca_DATA_SIZE4_3 is

   component FullAdder_9
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_10
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_11
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_12
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_12 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_11 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_10 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_9 port map( ci => carry_3_port, a => a(3), b => b(3), s =>
                           s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_2 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_2;

architecture SYN_rca_arch of Rca_DATA_SIZE4_2 is

   component FullAdder_5
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_6
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_7
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_8
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_8 port map( ci => ci, a => a(0), b => b(0), s => s(0), co 
                           => carry_1_port);
   FA3_1 : FullAdder_7 port map( ci => carry_1_port, a => a(1), b => b(1), s =>
                           s(1), co => carry_2_port);
   FA3_2 : FullAdder_6 port map( ci => carry_2_port, a => a(2), b => b(2), s =>
                           s(2), co => carry_3_port);
   FA3_3 : FullAdder_5 port map( ci => carry_3_port, a => a(3), b => b(3), s =>
                           s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_1 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_1;

architecture SYN_rca_arch of Rca_DATA_SIZE4_1 is

   component FullAdder_1
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_2
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_3
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_4
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_4 port map( ci => ci, a => a(0), b => b(0), s => s(0), co 
                           => carry_1_port);
   FA3_1 : FullAdder_3 port map( ci => carry_1_port, a => a(1), b => b(1), s =>
                           s(1), co => carry_2_port);
   FA3_2 : FullAdder_2 port map( ci => carry_2_port, a => a(2), b => b(2), s =>
                           s(2), co => carry_3_port);
   FA3_3 : FullAdder_1 port map( ci => carry_3_port, a => a(3), b => b(3), s =>
                           s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_83 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_83;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_83 is

   component Mux_DATA_SIZE4_83
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_165
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_166
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_166 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_165 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_83 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_82 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_82;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_82 is

   component Mux_DATA_SIZE4_82
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_163
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_164
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_164 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_163 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_82 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_81 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_81;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_81 is

   component Mux_DATA_SIZE4_81
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_161
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_162
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_162 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_161 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_81 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_80 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_80;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_80 is

   component Mux_DATA_SIZE4_80
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_159
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_160
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_160 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_159 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_80 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_79 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_79;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_79 is

   component Mux_DATA_SIZE4_79
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_157
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_158
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_158 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_157 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_79 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_78 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_78;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_78 is

   component Mux_DATA_SIZE4_78
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_155
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_156
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_156 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_155 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_78 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_77 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_77;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_77 is

   component Mux_DATA_SIZE4_77
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_153
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_154
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_154 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_153 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_77 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_76 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_76;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_76 is

   component Mux_DATA_SIZE4_76
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_151
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_152
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_152 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_151 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_76 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_75 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_75;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_75 is

   component Mux_DATA_SIZE4_75
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_149
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_150
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_150 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_149 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_75 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_74 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_74;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_74 is

   component Mux_DATA_SIZE4_74
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_147
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_148
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_148 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_147 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_74 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_73 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_73;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_73 is

   component Mux_DATA_SIZE4_73
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_145
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_146
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_146 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_145 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_73 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_72 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_72;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_72 is

   component Mux_DATA_SIZE4_72
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_143
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_144
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_144 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_143 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_72 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_71 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_71;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_71 is

   component Mux_DATA_SIZE4_71
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_141
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_142
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_142 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_141 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_71 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_70 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_70;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_70 is

   component Mux_DATA_SIZE4_70
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_139
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_140
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_140 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_139 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_70 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_69 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_69;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_69 is

   component Mux_DATA_SIZE4_69
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_137
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_138
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_138 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_137 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_69 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_68 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_68;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_68 is

   component Mux_DATA_SIZE4_68
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_135
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_136
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_136 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_135 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_68 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_67 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_67;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_67 is

   component Mux_DATA_SIZE4_67
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_133
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_134
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_134 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_133 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_67 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_66 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_66;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_66 is

   component Mux_DATA_SIZE4_66
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_131
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_132
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_132 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_131 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_66 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_65 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_65;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_65 is

   component Mux_DATA_SIZE4_65
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_129
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_130
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_130 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_129 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_65 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_64 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_64;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_64 is

   component Mux_DATA_SIZE4_64
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_127
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_128
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_128 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_127 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_64 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_63 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_63;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_63 is

   component Mux_DATA_SIZE4_63
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_125
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_126
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_126 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_125 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_63 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_62 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_62;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_62 is

   component Mux_DATA_SIZE4_62
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_123
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_124
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_124 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_123 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_62 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_61 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_61;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_61 is

   component Mux_DATA_SIZE4_61
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_121
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_122
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_122 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_121 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_61 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_60 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_60;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_60 is

   component Mux_DATA_SIZE4_60
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_119
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_120
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_120 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_119 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_60 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_59 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_59;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_59 is

   component Mux_DATA_SIZE4_59
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_117
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_118
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_118 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_117 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_59 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_58 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_58;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_58 is

   component Mux_DATA_SIZE4_58
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_115
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_116
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_116 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_115 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_58 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_57 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_57;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_57 is

   component Mux_DATA_SIZE4_57
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_113
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_114
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_114 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_113 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_57 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_56 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_56;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_56 is

   component Mux_DATA_SIZE4_56
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_111
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_112
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_112 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_111 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_56 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_55 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_55;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_55 is

   component Mux_DATA_SIZE4_55
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_109
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_110
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_110 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_109 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_55 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_54 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_54;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_54 is

   component Mux_DATA_SIZE4_54
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_107
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_108
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_108 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_107 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_54 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_53 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_53;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_53 is

   component Mux_DATA_SIZE4_53
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_105
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_106
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_106 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_105 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_53 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_52 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_52;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_52 is

   component Mux_DATA_SIZE4_52
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_103
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_104
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_104 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_103 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_52 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_51 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_51;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_51 is

   component Mux_DATA_SIZE4_51
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_101
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_102
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_102 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_101 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_51 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_50 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_50;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_50 is

   component Mux_DATA_SIZE4_50
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_99
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_100
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_100 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_99 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_50 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_49 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_49;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_49 is

   component Mux_DATA_SIZE4_49
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_97
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_98
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_98 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_97 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_49 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_48 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_48;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_48 is

   component Mux_DATA_SIZE4_48
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_95
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_96
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_96 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_95 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_48 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_47 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_47;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_47 is

   component Mux_DATA_SIZE4_47
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_93
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_94
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_94 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_93 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_47 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_46 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_46;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_46 is

   component Mux_DATA_SIZE4_46
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_91
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_92
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_92 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_91 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_46 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_45 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_45;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_45 is

   component Mux_DATA_SIZE4_45
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_89
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_90
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_90 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_89 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_45 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_44 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_44;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_44 is

   component Mux_DATA_SIZE4_44
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_87
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_88
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_88 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_87 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_44 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_43 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_43;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_43 is

   component Mux_DATA_SIZE4_43
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_85
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_86
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_86 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_85 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_43 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_42 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_42;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_42 is

   component Mux_DATA_SIZE4_42
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_83
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_84
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_84 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_83 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_42 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_41 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_41;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_41 is

   component Mux_DATA_SIZE4_41
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_81
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_82
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_82 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_81 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_41 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_40 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_40;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_40 is

   component Mux_DATA_SIZE4_40
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_79
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_80
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_80 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_79 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_40 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_39 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_39;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_39 is

   component Mux_DATA_SIZE4_39
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_77
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_78
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_78 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_77 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_39 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_38 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_38;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_38 is

   component Mux_DATA_SIZE4_38
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_75
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_76
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_76 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_75 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_38 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_37 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_37;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_37 is

   component Mux_DATA_SIZE4_37
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_73
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_74
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_74 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_73 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_37 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_36 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_36;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_36 is

   component Mux_DATA_SIZE4_36
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_71
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_72
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_72 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_71 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_36 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_35 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_35;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_35 is

   component Mux_DATA_SIZE4_35
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_69
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_70
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_70 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_69 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_35 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_34 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_34;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_34 is

   component Mux_DATA_SIZE4_34
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_67
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_68
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_68 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_67 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_34 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_33 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_33;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_33 is

   component Mux_DATA_SIZE4_33
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_65
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_66
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_66 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_65 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_33 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_32 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_32;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_32 is

   component Mux_DATA_SIZE4_32
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_63
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_64
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_64 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_63 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_32 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_31 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_31;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_31 is

   component Mux_DATA_SIZE4_31
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_61
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_62
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_62 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_61 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_31 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_30 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_30;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_30 is

   component Mux_DATA_SIZE4_30
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_59
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_60
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_60 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_59 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_30 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_29 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_29;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_29 is

   component Mux_DATA_SIZE4_29
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_57
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_58
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_58 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_57 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_29 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_28 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_28;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_28 is

   component Mux_DATA_SIZE4_28
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_55
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_56
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_56 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_55 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_28 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_27 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_27;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_27 is

   component Mux_DATA_SIZE4_27
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_53
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_54
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_54 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_53 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_27 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_26 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_26;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_26 is

   component Mux_DATA_SIZE4_26
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_51
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_52
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_52 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_51 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_26 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_25 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_25;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_25 is

   component Mux_DATA_SIZE4_25
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_49
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_50
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_50 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_49 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_25 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_24 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_24;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_24 is

   component Mux_DATA_SIZE4_24
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_47
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_48
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_48 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_47 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_24 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_23 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_23;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_23 is

   component Mux_DATA_SIZE4_23
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_45
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_46
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_46 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_45 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_23 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_22 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_22;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_22 is

   component Mux_DATA_SIZE4_22
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_43
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_44
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_44 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_43 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_22 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_21 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_21;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_21 is

   component Mux_DATA_SIZE4_21
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_41
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_42
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_42 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_41 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_21 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_20 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_20;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_20 is

   component Mux_DATA_SIZE4_20
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_39
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_40
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_40 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_39 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_20 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_19 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_19;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_19 is

   component Mux_DATA_SIZE4_19
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_37
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_38
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_38 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_37 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_19 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_18 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_18;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_18 is

   component Mux_DATA_SIZE4_18
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_35
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_36
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_36 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_35 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_18 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_17 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_17;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_17 is

   component Mux_DATA_SIZE4_17
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_33
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_34
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_34 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_33 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_17 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_16 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_16;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_16 is

   component Mux_DATA_SIZE4_16
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_31
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_32
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_32 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_31 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_16 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_15 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_15;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_15 is

   component Mux_DATA_SIZE4_15
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_29
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_30
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_30 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_29 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_15 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_14 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_14;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_14 is

   component Mux_DATA_SIZE4_14
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_27
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_28
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_28 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_27 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_14 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_13 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_13;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_13 is

   component Mux_DATA_SIZE4_13
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_25
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_26
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_26 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_25 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_13 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_12 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_12;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_12 is

   component Mux_DATA_SIZE4_12
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_23
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_24
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_24 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_23 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_12 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_11 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_11;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_11 is

   component Mux_DATA_SIZE4_11
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_21
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_22
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_22 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_21 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_11 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_10 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_10;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_10 is

   component Mux_DATA_SIZE4_10
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_19
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_20
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_20 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_19 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_10 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_9 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_9;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_9 is

   component Mux_DATA_SIZE4_9
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_17
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_18
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_18 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_17 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_9 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_8 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_8;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_8 is

   component Mux_DATA_SIZE4_8
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_15
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_16
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_16 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_15 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_8 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_7 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_7;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_7 is

   component Mux_DATA_SIZE4_7
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_13
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_14
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_14 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_13 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_7 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_6 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_6;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_6 is

   component Mux_DATA_SIZE4_6
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_11
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_12
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_12 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_11 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_6 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_5 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_5;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_5 is

   component Mux_DATA_SIZE4_5
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_9
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_10
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_10 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_9 port map( ci => X_Logic1_port, a(3) => a(3), a(2) =>
                           a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2)
                           => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_5 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_4 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_4;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_4 is

   component Mux_DATA_SIZE4_4
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_7
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_8
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_8 port map( ci => X_Logic0_port, a(3) => a(3), a(2) =>
                           a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2)
                           => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_7 port map( ci => X_Logic1_port, a(3) => a(3), a(2) =>
                           a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2)
                           => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_4 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_3 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_3;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_3 is

   component Mux_DATA_SIZE4_3
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_5
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_6
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_6 port map( ci => X_Logic0_port, a(3) => a(3), a(2) =>
                           a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2)
                           => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_5 port map( ci => X_Logic1_port, a(3) => a(3), a(2) =>
                           a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2)
                           => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_3 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_2 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_2;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_2 is

   component Mux_DATA_SIZE4_2
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_3
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_4
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_4 port map( ci => X_Logic0_port, a(3) => a(3), a(2) =>
                           a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2)
                           => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_3 port map( ci => X_Logic1_port, a(3) => a(3), a(2) =>
                           a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2)
                           => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_2 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_1 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_1;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_1 is

   component Mux_DATA_SIZE4_1
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_1
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_2
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_2 port map( ci => X_Logic0_port, a(3) => a(3), a(2) =>
                           a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2)
                           => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_1 port map( ci => X_Logic1_port, a(3) => a(3), a(2) =>
                           a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2)
                           => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_1 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderSumGenerator_DATA_SIZE32_SPARSITY4_7 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic_vector 
         (7 downto 0);  sum : out std_logic_vector (31 downto 0));

end AdderSumGenerator_DATA_SIZE32_SPARSITY4_7;

architecture SYN_adder_sum_generator_arch of 
   AdderSumGenerator_DATA_SIZE32_SPARSITY4_7 is

   component AdderCarrySelect_DATA_SIZE4_69
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_70
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_71
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_72
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_73
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_74
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_75
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_76
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;

begin
   
   ACSi_0 : AdderCarrySelect_DATA_SIZE4_76 port map( a(3) => a(3), a(2) => a(2)
                           , a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), sel => cin(0), 
                           sum(3) => sum(3), sum(2) => sum(2), sum(1) => sum(1)
                           , sum(0) => sum(0));
   ACSi_1 : AdderCarrySelect_DATA_SIZE4_75 port map( a(3) => a(7), a(2) => a(6)
                           , a(1) => a(5), a(0) => a(4), b(3) => b(7), b(2) => 
                           b(6), b(1) => b(5), b(0) => b(4), sel => cin(1), 
                           sum(3) => sum(7), sum(2) => sum(6), sum(1) => sum(5)
                           , sum(0) => sum(4));
   ACSi_2 : AdderCarrySelect_DATA_SIZE4_74 port map( a(3) => a(11), a(2) => 
                           a(10), a(1) => a(9), a(0) => a(8), b(3) => b(11), 
                           b(2) => b(10), b(1) => b(9), b(0) => b(8), sel => 
                           cin(2), sum(3) => sum(11), sum(2) => sum(10), sum(1)
                           => sum(9), sum(0) => sum(8));
   ACSi_3 : AdderCarrySelect_DATA_SIZE4_73 port map( a(3) => a(15), a(2) => 
                           a(14), a(1) => a(13), a(0) => a(12), b(3) => b(15), 
                           b(2) => b(14), b(1) => b(13), b(0) => b(12), sel => 
                           cin(3), sum(3) => sum(15), sum(2) => sum(14), sum(1)
                           => sum(13), sum(0) => sum(12));
   ACSi_4 : AdderCarrySelect_DATA_SIZE4_72 port map( a(3) => a(19), a(2) => 
                           a(18), a(1) => a(17), a(0) => a(16), b(3) => b(19), 
                           b(2) => b(18), b(1) => b(17), b(0) => b(16), sel => 
                           cin(4), sum(3) => sum(19), sum(2) => sum(18), sum(1)
                           => sum(17), sum(0) => sum(16));
   ACSi_5 : AdderCarrySelect_DATA_SIZE4_71 port map( a(3) => a(23), a(2) => 
                           a(22), a(1) => a(21), a(0) => a(20), b(3) => b(23), 
                           b(2) => b(22), b(1) => b(21), b(0) => b(20), sel => 
                           cin(5), sum(3) => sum(23), sum(2) => sum(22), sum(1)
                           => sum(21), sum(0) => sum(20));
   ACSi_6 : AdderCarrySelect_DATA_SIZE4_70 port map( a(3) => a(27), a(2) => 
                           a(26), a(1) => a(25), a(0) => a(24), b(3) => b(27), 
                           b(2) => b(26), b(1) => b(25), b(0) => b(24), sel => 
                           cin(6), sum(3) => sum(27), sum(2) => sum(26), sum(1)
                           => sum(25), sum(0) => sum(24));
   ACSi_7 : AdderCarrySelect_DATA_SIZE4_69 port map( a(3) => a(31), a(2) => 
                           a(30), a(1) => a(29), a(0) => a(28), b(3) => b(31), 
                           b(2) => b(30), b(1) => b(29), b(0) => b(28), sel => 
                           cin(7), sum(3) => sum(31), sum(2) => sum(30), sum(1)
                           => sum(29), sum(0) => sum(28));

end SYN_adder_sum_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderSumGenerator_DATA_SIZE32_SPARSITY4_6 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic_vector 
         (7 downto 0);  sum : out std_logic_vector (31 downto 0));

end AdderSumGenerator_DATA_SIZE32_SPARSITY4_6;

architecture SYN_adder_sum_generator_arch of 
   AdderSumGenerator_DATA_SIZE32_SPARSITY4_6 is

   component AdderCarrySelect_DATA_SIZE4_61
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_62
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_63
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_64
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_65
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_66
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_67
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_68
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;

begin
   
   ACSi_0 : AdderCarrySelect_DATA_SIZE4_68 port map( a(3) => a(3), a(2) => a(2)
                           , a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), sel => cin(0), 
                           sum(3) => sum(3), sum(2) => sum(2), sum(1) => sum(1)
                           , sum(0) => sum(0));
   ACSi_1 : AdderCarrySelect_DATA_SIZE4_67 port map( a(3) => a(7), a(2) => a(6)
                           , a(1) => a(5), a(0) => a(4), b(3) => b(7), b(2) => 
                           b(6), b(1) => b(5), b(0) => b(4), sel => cin(1), 
                           sum(3) => sum(7), sum(2) => sum(6), sum(1) => sum(5)
                           , sum(0) => sum(4));
   ACSi_2 : AdderCarrySelect_DATA_SIZE4_66 port map( a(3) => a(11), a(2) => 
                           a(10), a(1) => a(9), a(0) => a(8), b(3) => b(11), 
                           b(2) => b(10), b(1) => b(9), b(0) => b(8), sel => 
                           cin(2), sum(3) => sum(11), sum(2) => sum(10), sum(1)
                           => sum(9), sum(0) => sum(8));
   ACSi_3 : AdderCarrySelect_DATA_SIZE4_65 port map( a(3) => a(15), a(2) => 
                           a(14), a(1) => a(13), a(0) => a(12), b(3) => b(15), 
                           b(2) => b(14), b(1) => b(13), b(0) => b(12), sel => 
                           cin(3), sum(3) => sum(15), sum(2) => sum(14), sum(1)
                           => sum(13), sum(0) => sum(12));
   ACSi_4 : AdderCarrySelect_DATA_SIZE4_64 port map( a(3) => a(19), a(2) => 
                           a(18), a(1) => a(17), a(0) => a(16), b(3) => b(19), 
                           b(2) => b(18), b(1) => b(17), b(0) => b(16), sel => 
                           cin(4), sum(3) => sum(19), sum(2) => sum(18), sum(1)
                           => sum(17), sum(0) => sum(16));
   ACSi_5 : AdderCarrySelect_DATA_SIZE4_63 port map( a(3) => a(23), a(2) => 
                           a(22), a(1) => a(21), a(0) => a(20), b(3) => b(23), 
                           b(2) => b(22), b(1) => b(21), b(0) => b(20), sel => 
                           cin(5), sum(3) => sum(23), sum(2) => sum(22), sum(1)
                           => sum(21), sum(0) => sum(20));
   ACSi_6 : AdderCarrySelect_DATA_SIZE4_62 port map( a(3) => a(27), a(2) => 
                           a(26), a(1) => a(25), a(0) => a(24), b(3) => b(27), 
                           b(2) => b(26), b(1) => b(25), b(0) => b(24), sel => 
                           cin(6), sum(3) => sum(27), sum(2) => sum(26), sum(1)
                           => sum(25), sum(0) => sum(24));
   ACSi_7 : AdderCarrySelect_DATA_SIZE4_61 port map( a(3) => a(31), a(2) => 
                           a(30), a(1) => a(29), a(0) => a(28), b(3) => b(31), 
                           b(2) => b(30), b(1) => b(29), b(0) => b(28), sel => 
                           cin(7), sum(3) => sum(31), sum(2) => sum(30), sum(1)
                           => sum(29), sum(0) => sum(28));

end SYN_adder_sum_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderSumGenerator_DATA_SIZE32_SPARSITY4_5 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic_vector 
         (7 downto 0);  sum : out std_logic_vector (31 downto 0));

end AdderSumGenerator_DATA_SIZE32_SPARSITY4_5;

architecture SYN_adder_sum_generator_arch of 
   AdderSumGenerator_DATA_SIZE32_SPARSITY4_5 is

   component AdderCarrySelect_DATA_SIZE4_49
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_50
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_51
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_52
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_53
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_54
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_55
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_56
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;

begin
   
   ACSi_0 : AdderCarrySelect_DATA_SIZE4_56 port map( a(3) => a(3), a(2) => a(2)
                           , a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), sel => cin(0), 
                           sum(3) => sum(3), sum(2) => sum(2), sum(1) => sum(1)
                           , sum(0) => sum(0));
   ACSi_1 : AdderCarrySelect_DATA_SIZE4_55 port map( a(3) => a(7), a(2) => a(6)
                           , a(1) => a(5), a(0) => a(4), b(3) => b(7), b(2) => 
                           b(6), b(1) => b(5), b(0) => b(4), sel => cin(1), 
                           sum(3) => sum(7), sum(2) => sum(6), sum(1) => sum(5)
                           , sum(0) => sum(4));
   ACSi_2 : AdderCarrySelect_DATA_SIZE4_54 port map( a(3) => a(11), a(2) => 
                           a(10), a(1) => a(9), a(0) => a(8), b(3) => b(11), 
                           b(2) => b(10), b(1) => b(9), b(0) => b(8), sel => 
                           cin(2), sum(3) => sum(11), sum(2) => sum(10), sum(1)
                           => sum(9), sum(0) => sum(8));
   ACSi_3 : AdderCarrySelect_DATA_SIZE4_53 port map( a(3) => a(15), a(2) => 
                           a(14), a(1) => a(13), a(0) => a(12), b(3) => b(15), 
                           b(2) => b(14), b(1) => b(13), b(0) => b(12), sel => 
                           cin(3), sum(3) => sum(15), sum(2) => sum(14), sum(1)
                           => sum(13), sum(0) => sum(12));
   ACSi_4 : AdderCarrySelect_DATA_SIZE4_52 port map( a(3) => a(19), a(2) => 
                           a(18), a(1) => a(17), a(0) => a(16), b(3) => b(19), 
                           b(2) => b(18), b(1) => b(17), b(0) => b(16), sel => 
                           cin(4), sum(3) => sum(19), sum(2) => sum(18), sum(1)
                           => sum(17), sum(0) => sum(16));
   ACSi_5 : AdderCarrySelect_DATA_SIZE4_51 port map( a(3) => a(23), a(2) => 
                           a(22), a(1) => a(21), a(0) => a(20), b(3) => b(23), 
                           b(2) => b(22), b(1) => b(21), b(0) => b(20), sel => 
                           cin(5), sum(3) => sum(23), sum(2) => sum(22), sum(1)
                           => sum(21), sum(0) => sum(20));
   ACSi_6 : AdderCarrySelect_DATA_SIZE4_50 port map( a(3) => a(27), a(2) => 
                           a(26), a(1) => a(25), a(0) => a(24), b(3) => b(27), 
                           b(2) => b(26), b(1) => b(25), b(0) => b(24), sel => 
                           cin(6), sum(3) => sum(27), sum(2) => sum(26), sum(1)
                           => sum(25), sum(0) => sum(24));
   ACSi_7 : AdderCarrySelect_DATA_SIZE4_49 port map( a(3) => a(31), a(2) => 
                           a(30), a(1) => a(29), a(0) => a(28), b(3) => b(31), 
                           b(2) => b(30), b(1) => b(29), b(0) => b(28), sel => 
                           cin(7), sum(3) => sum(31), sum(2) => sum(30), sum(1)
                           => sum(29), sum(0) => sum(28));

end SYN_adder_sum_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderSumGenerator_DATA_SIZE32_SPARSITY4_4 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic_vector 
         (7 downto 0);  sum : out std_logic_vector (31 downto 0));

end AdderSumGenerator_DATA_SIZE32_SPARSITY4_4;

architecture SYN_adder_sum_generator_arch of 
   AdderSumGenerator_DATA_SIZE32_SPARSITY4_4 is

   component AdderCarrySelect_DATA_SIZE4_41
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_42
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_43
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_44
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_45
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_46
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_47
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_48
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;

begin
   
   ACSi_0 : AdderCarrySelect_DATA_SIZE4_48 port map( a(3) => a(3), a(2) => a(2)
                           , a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), sel => cin(0), 
                           sum(3) => sum(3), sum(2) => sum(2), sum(1) => sum(1)
                           , sum(0) => sum(0));
   ACSi_1 : AdderCarrySelect_DATA_SIZE4_47 port map( a(3) => a(7), a(2) => a(6)
                           , a(1) => a(5), a(0) => a(4), b(3) => b(7), b(2) => 
                           b(6), b(1) => b(5), b(0) => b(4), sel => cin(1), 
                           sum(3) => sum(7), sum(2) => sum(6), sum(1) => sum(5)
                           , sum(0) => sum(4));
   ACSi_2 : AdderCarrySelect_DATA_SIZE4_46 port map( a(3) => a(11), a(2) => 
                           a(10), a(1) => a(9), a(0) => a(8), b(3) => b(11), 
                           b(2) => b(10), b(1) => b(9), b(0) => b(8), sel => 
                           cin(2), sum(3) => sum(11), sum(2) => sum(10), sum(1)
                           => sum(9), sum(0) => sum(8));
   ACSi_3 : AdderCarrySelect_DATA_SIZE4_45 port map( a(3) => a(15), a(2) => 
                           a(14), a(1) => a(13), a(0) => a(12), b(3) => b(15), 
                           b(2) => b(14), b(1) => b(13), b(0) => b(12), sel => 
                           cin(3), sum(3) => sum(15), sum(2) => sum(14), sum(1)
                           => sum(13), sum(0) => sum(12));
   ACSi_4 : AdderCarrySelect_DATA_SIZE4_44 port map( a(3) => a(19), a(2) => 
                           a(18), a(1) => a(17), a(0) => a(16), b(3) => b(19), 
                           b(2) => b(18), b(1) => b(17), b(0) => b(16), sel => 
                           cin(4), sum(3) => sum(19), sum(2) => sum(18), sum(1)
                           => sum(17), sum(0) => sum(16));
   ACSi_5 : AdderCarrySelect_DATA_SIZE4_43 port map( a(3) => a(23), a(2) => 
                           a(22), a(1) => a(21), a(0) => a(20), b(3) => b(23), 
                           b(2) => b(22), b(1) => b(21), b(0) => b(20), sel => 
                           cin(5), sum(3) => sum(23), sum(2) => sum(22), sum(1)
                           => sum(21), sum(0) => sum(20));
   ACSi_6 : AdderCarrySelect_DATA_SIZE4_42 port map( a(3) => a(27), a(2) => 
                           a(26), a(1) => a(25), a(0) => a(24), b(3) => b(27), 
                           b(2) => b(26), b(1) => b(25), b(0) => b(24), sel => 
                           cin(6), sum(3) => sum(27), sum(2) => sum(26), sum(1)
                           => sum(25), sum(0) => sum(24));
   ACSi_7 : AdderCarrySelect_DATA_SIZE4_41 port map( a(3) => a(31), a(2) => 
                           a(30), a(1) => a(29), a(0) => a(28), b(3) => b(31), 
                           b(2) => b(30), b(1) => b(29), b(0) => b(28), sel => 
                           cin(7), sum(3) => sum(31), sum(2) => sum(30), sum(1)
                           => sum(29), sum(0) => sum(28));

end SYN_adder_sum_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderSumGenerator_DATA_SIZE32_SPARSITY4_3 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic_vector 
         (7 downto 0);  sum : out std_logic_vector (31 downto 0));

end AdderSumGenerator_DATA_SIZE32_SPARSITY4_3;

architecture SYN_adder_sum_generator_arch of 
   AdderSumGenerator_DATA_SIZE32_SPARSITY4_3 is

   component AdderCarrySelect_DATA_SIZE4_33
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_34
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_35
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_36
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_37
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_38
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_39
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_40
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;

begin
   
   ACSi_0 : AdderCarrySelect_DATA_SIZE4_40 port map( a(3) => a(3), a(2) => a(2)
                           , a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), sel => cin(0), 
                           sum(3) => sum(3), sum(2) => sum(2), sum(1) => sum(1)
                           , sum(0) => sum(0));
   ACSi_1 : AdderCarrySelect_DATA_SIZE4_39 port map( a(3) => a(7), a(2) => a(6)
                           , a(1) => a(5), a(0) => a(4), b(3) => b(7), b(2) => 
                           b(6), b(1) => b(5), b(0) => b(4), sel => cin(1), 
                           sum(3) => sum(7), sum(2) => sum(6), sum(1) => sum(5)
                           , sum(0) => sum(4));
   ACSi_2 : AdderCarrySelect_DATA_SIZE4_38 port map( a(3) => a(11), a(2) => 
                           a(10), a(1) => a(9), a(0) => a(8), b(3) => b(11), 
                           b(2) => b(10), b(1) => b(9), b(0) => b(8), sel => 
                           cin(2), sum(3) => sum(11), sum(2) => sum(10), sum(1)
                           => sum(9), sum(0) => sum(8));
   ACSi_3 : AdderCarrySelect_DATA_SIZE4_37 port map( a(3) => a(15), a(2) => 
                           a(14), a(1) => a(13), a(0) => a(12), b(3) => b(15), 
                           b(2) => b(14), b(1) => b(13), b(0) => b(12), sel => 
                           cin(3), sum(3) => sum(15), sum(2) => sum(14), sum(1)
                           => sum(13), sum(0) => sum(12));
   ACSi_4 : AdderCarrySelect_DATA_SIZE4_36 port map( a(3) => a(19), a(2) => 
                           a(18), a(1) => a(17), a(0) => a(16), b(3) => b(19), 
                           b(2) => b(18), b(1) => b(17), b(0) => b(16), sel => 
                           cin(4), sum(3) => sum(19), sum(2) => sum(18), sum(1)
                           => sum(17), sum(0) => sum(16));
   ACSi_5 : AdderCarrySelect_DATA_SIZE4_35 port map( a(3) => a(23), a(2) => 
                           a(22), a(1) => a(21), a(0) => a(20), b(3) => b(23), 
                           b(2) => b(22), b(1) => b(21), b(0) => b(20), sel => 
                           cin(5), sum(3) => sum(23), sum(2) => sum(22), sum(1)
                           => sum(21), sum(0) => sum(20));
   ACSi_6 : AdderCarrySelect_DATA_SIZE4_34 port map( a(3) => a(27), a(2) => 
                           a(26), a(1) => a(25), a(0) => a(24), b(3) => b(27), 
                           b(2) => b(26), b(1) => b(25), b(0) => b(24), sel => 
                           cin(6), sum(3) => sum(27), sum(2) => sum(26), sum(1)
                           => sum(25), sum(0) => sum(24));
   ACSi_7 : AdderCarrySelect_DATA_SIZE4_33 port map( a(3) => a(31), a(2) => 
                           a(30), a(1) => a(29), a(0) => a(28), b(3) => b(31), 
                           b(2) => b(30), b(1) => b(29), b(0) => b(28), sel => 
                           cin(7), sum(3) => sum(31), sum(2) => sum(30), sum(1)
                           => sum(29), sum(0) => sum(28));

end SYN_adder_sum_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderSumGenerator_DATA_SIZE32_SPARSITY4_2 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic_vector 
         (7 downto 0);  sum : out std_logic_vector (31 downto 0));

end AdderSumGenerator_DATA_SIZE32_SPARSITY4_2;

architecture SYN_adder_sum_generator_arch of 
   AdderSumGenerator_DATA_SIZE32_SPARSITY4_2 is

   component AdderCarrySelect_DATA_SIZE4_9
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_10
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_11
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_12
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_13
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_14
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_15
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_16
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;

begin
   
   ACSi_0 : AdderCarrySelect_DATA_SIZE4_16 port map( a(3) => a(3), a(2) => a(2)
                           , a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), sel => cin(0), 
                           sum(3) => sum(3), sum(2) => sum(2), sum(1) => sum(1)
                           , sum(0) => sum(0));
   ACSi_1 : AdderCarrySelect_DATA_SIZE4_15 port map( a(3) => a(7), a(2) => a(6)
                           , a(1) => a(5), a(0) => a(4), b(3) => b(7), b(2) => 
                           b(6), b(1) => b(5), b(0) => b(4), sel => cin(1), 
                           sum(3) => sum(7), sum(2) => sum(6), sum(1) => sum(5)
                           , sum(0) => sum(4));
   ACSi_2 : AdderCarrySelect_DATA_SIZE4_14 port map( a(3) => a(11), a(2) => 
                           a(10), a(1) => a(9), a(0) => a(8), b(3) => b(11), 
                           b(2) => b(10), b(1) => b(9), b(0) => b(8), sel => 
                           cin(2), sum(3) => sum(11), sum(2) => sum(10), sum(1)
                           => sum(9), sum(0) => sum(8));
   ACSi_3 : AdderCarrySelect_DATA_SIZE4_13 port map( a(3) => a(15), a(2) => 
                           a(14), a(1) => a(13), a(0) => a(12), b(3) => b(15), 
                           b(2) => b(14), b(1) => b(13), b(0) => b(12), sel => 
                           cin(3), sum(3) => sum(15), sum(2) => sum(14), sum(1)
                           => sum(13), sum(0) => sum(12));
   ACSi_4 : AdderCarrySelect_DATA_SIZE4_12 port map( a(3) => a(19), a(2) => 
                           a(18), a(1) => a(17), a(0) => a(16), b(3) => b(19), 
                           b(2) => b(18), b(1) => b(17), b(0) => b(16), sel => 
                           cin(4), sum(3) => sum(19), sum(2) => sum(18), sum(1)
                           => sum(17), sum(0) => sum(16));
   ACSi_5 : AdderCarrySelect_DATA_SIZE4_11 port map( a(3) => a(23), a(2) => 
                           a(22), a(1) => a(21), a(0) => a(20), b(3) => b(23), 
                           b(2) => b(22), b(1) => b(21), b(0) => b(20), sel => 
                           cin(5), sum(3) => sum(23), sum(2) => sum(22), sum(1)
                           => sum(21), sum(0) => sum(20));
   ACSi_6 : AdderCarrySelect_DATA_SIZE4_10 port map( a(3) => a(27), a(2) => 
                           a(26), a(1) => a(25), a(0) => a(24), b(3) => b(27), 
                           b(2) => b(26), b(1) => b(25), b(0) => b(24), sel => 
                           cin(6), sum(3) => sum(27), sum(2) => sum(26), sum(1)
                           => sum(25), sum(0) => sum(24));
   ACSi_7 : AdderCarrySelect_DATA_SIZE4_9 port map( a(3) => a(31), a(2) => 
                           a(30), a(1) => a(29), a(0) => a(28), b(3) => b(31), 
                           b(2) => b(30), b(1) => b(29), b(0) => b(28), sel => 
                           cin(7), sum(3) => sum(31), sum(2) => sum(30), sum(1)
                           => sum(29), sum(0) => sum(28));

end SYN_adder_sum_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderSumGenerator_DATA_SIZE32_SPARSITY4_1 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic_vector 
         (7 downto 0);  sum : out std_logic_vector (31 downto 0));

end AdderSumGenerator_DATA_SIZE32_SPARSITY4_1;

architecture SYN_adder_sum_generator_arch of 
   AdderSumGenerator_DATA_SIZE32_SPARSITY4_1 is

   component AdderCarrySelect_DATA_SIZE4_1
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_2
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_3
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_4
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_5
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_6
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_7
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_8
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;

begin
   
   ACSi_0 : AdderCarrySelect_DATA_SIZE4_8 port map( a(3) => a(3), a(2) => a(2),
                           a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), sel => cin(0), 
                           sum(3) => sum(3), sum(2) => sum(2), sum(1) => sum(1)
                           , sum(0) => sum(0));
   ACSi_1 : AdderCarrySelect_DATA_SIZE4_7 port map( a(3) => a(7), a(2) => a(6),
                           a(1) => a(5), a(0) => a(4), b(3) => b(7), b(2) => 
                           b(6), b(1) => b(5), b(0) => b(4), sel => cin(1), 
                           sum(3) => sum(7), sum(2) => sum(6), sum(1) => sum(5)
                           , sum(0) => sum(4));
   ACSi_2 : AdderCarrySelect_DATA_SIZE4_6 port map( a(3) => a(11), a(2) => 
                           a(10), a(1) => a(9), a(0) => a(8), b(3) => b(11), 
                           b(2) => b(10), b(1) => b(9), b(0) => b(8), sel => 
                           cin(2), sum(3) => sum(11), sum(2) => sum(10), sum(1)
                           => sum(9), sum(0) => sum(8));
   ACSi_3 : AdderCarrySelect_DATA_SIZE4_5 port map( a(3) => a(15), a(2) => 
                           a(14), a(1) => a(13), a(0) => a(12), b(3) => b(15), 
                           b(2) => b(14), b(1) => b(13), b(0) => b(12), sel => 
                           cin(3), sum(3) => sum(15), sum(2) => sum(14), sum(1)
                           => sum(13), sum(0) => sum(12));
   ACSi_4 : AdderCarrySelect_DATA_SIZE4_4 port map( a(3) => a(19), a(2) => 
                           a(18), a(1) => a(17), a(0) => a(16), b(3) => b(19), 
                           b(2) => b(18), b(1) => b(17), b(0) => b(16), sel => 
                           cin(4), sum(3) => sum(19), sum(2) => sum(18), sum(1)
                           => sum(17), sum(0) => sum(16));
   ACSi_5 : AdderCarrySelect_DATA_SIZE4_3 port map( a(3) => a(23), a(2) => 
                           a(22), a(1) => a(21), a(0) => a(20), b(3) => b(23), 
                           b(2) => b(22), b(1) => b(21), b(0) => b(20), sel => 
                           cin(5), sum(3) => sum(23), sum(2) => sum(22), sum(1)
                           => sum(21), sum(0) => sum(20));
   ACSi_6 : AdderCarrySelect_DATA_SIZE4_2 port map( a(3) => a(27), a(2) => 
                           a(26), a(1) => a(25), a(0) => a(24), b(3) => b(27), 
                           b(2) => b(26), b(1) => b(25), b(0) => b(24), sel => 
                           cin(6), sum(3) => sum(27), sum(2) => sum(26), sum(1)
                           => sum(25), sum(0) => sum(24));
   ACSi_7 : AdderCarrySelect_DATA_SIZE4_1 port map( a(3) => a(31), a(2) => 
                           a(30), a(1) => a(29), a(0) => a(28), b(3) => b(31), 
                           b(2) => b(30), b(1) => b(29), b(0) => b(28), sel => 
                           cin(7), sum(3) => sum(31), sum(2) => sum(30), sum(1)
                           => sum(29), sum(0) => sum(28));

end SYN_adder_sum_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4CarryGenerator_DATA_SIZE32_SPARSITY4_7 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  cout :
         out std_logic_vector (7 downto 0));

end P4CarryGenerator_DATA_SIZE32_SPARSITY4_7;

architecture SYN_p4_carry_generator_arch of 
   P4CarryGenerator_DATA_SIZE32_SPARSITY4_7 is

   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal cout_7_port, n250, n251, n252, cout_0_port, n61, n63, n64, n102, n103
      , n111, n121, net138600, net138780, net138777, net138989, net139124, 
      net139150, net139158, net150681, net151348, net151510, net151886, 
      net153886, n104, n105, n106, n107, n108, n109, n110, n113, n114, n115, 
      n116, n117, n118, n119, n120, n123, n124, n125, n126, n127, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, 
      n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, 
      n190, n191, n192, n193, cout_2_port, cout_5_port, n196, cout_6_port, n198
      , n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      cout_3_port, n211, n212, cout_1_port, n214, n215, n216, n217, n218, n219,
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n245, n246, n247, n248, n249 : std_logic;

begin
   cout <= ( cout_7_port, cout_6_port, cout_5_port, net151348, cout_3_port, 
      cout_2_port, cout_1_port, cout_0_port );
   
   syn264 : NAND3_X1 port map( A1 => n179, A2 => n174, A3 => n180, ZN => n184);
   syn249 : NAND3_X1 port map( A1 => n110, A2 => a(15), A3 => n131, ZN => n150)
                           ;
   U1 : INV_X1 port map( A => a(3), ZN => n165);
   U2 : NAND2_X1 port map( A1 => net150681, A2 => n169, ZN => n186);
   U3 : INV_X1 port map( A => a(6), ZN => n169);
   U4 : NAND2_X1 port map( A1 => net150681, A2 => n168, ZN => n185);
   U5 : INV_X1 port map( A => b(6), ZN => n168);
   U6 : NAND2_X1 port map( A1 => n133, A2 => n153, ZN => n152);
   U7 : INV_X1 port map( A => a(20), ZN => n133);
   U8 : INV_X1 port map( A => b(20), ZN => n143);
   U9 : NOR2_X1 port map( A1 => a(21), A2 => b(21), ZN => n134);
   U10 : INV_X1 port map( A => b(21), ZN => n64);
   U11 : NAND2_X1 port map( A1 => n124, A2 => n123, ZN => n138);
   U12 : INV_X1 port map( A => a(17), ZN => n123);
   U13 : INV_X1 port map( A => b(17), ZN => n124);
   U14 : OAI21_X1 port map( B1 => n115, B2 => n116, A => n117, ZN => n114);
   U15 : NAND2_X1 port map( A1 => b(16), A2 => a(16), ZN => n116);
   U16 : NAND2_X1 port map( A1 => b(17), A2 => a(17), ZN => n117);
   U17 : INV_X1 port map( A => n138, ZN => n115);
   U18 : NAND2_X1 port map( A1 => n136, A2 => n138, ZN => n137);
   U19 : NOR2_X1 port map( A1 => n129, A2 => n128, ZN => n136);
   U20 : NOR2_X1 port map( A1 => a(18), A2 => b(18), ZN => n128);
   U21 : NOR2_X1 port map( A1 => a(19), A2 => b(19), ZN => n129);
   U22 : INV_X1 port map( A => b(15), ZN => n146);
   U23 : INV_X1 port map( A => b(16), ZN => n125);
   U24 : INV_X1 port map( A => a(16), ZN => n126);
   U25 : NOR2_X1 port map( A1 => n114, A2 => a(18), ZN => n127);
   U26 : NOR2_X1 port map( A1 => b(19), A2 => a(19), ZN => n132);
   U27 : NAND2_X1 port map( A1 => n114, A2 => a(18), ZN => n148);
   U28 : INV_X1 port map( A => b(18), ZN => n147);
   U29 : NAND2_X1 port map( A1 => n160, A2 => net138600, ZN => n181);
   U30 : NOR2_X1 port map( A1 => n160, A2 => net138600, ZN => n172);
   U31 : INV_X1 port map( A => a(7), ZN => n102);
   U32 : NAND2_X1 port map( A1 => a(6), A2 => b(6), ZN => n187);
   U33 : NAND2_X1 port map( A1 => n186, A2 => n185, ZN => n171);
   U34 : NAND2_X1 port map( A1 => n185, A2 => n186, ZN => n163);
   U35 : INV_X1 port map( A => a(21), ZN => n63);
   U36 : INV_X1 port map( A => a(1), ZN => n173);
   U37 : INV_X1 port map( A => a(2), ZN => n178);
   U38 : INV_X1 port map( A => b(5), ZN => n160);
   U39 : NAND2_X1 port map( A1 => n176, A2 => n178, ZN => n180);
   U40 : NAND2_X1 port map( A1 => n125, A2 => n126, ZN => n151);
   U41 : NAND2_X1 port map( A1 => n148, A2 => n147, ZN => n140);
   U42 : NOR2_X1 port map( A1 => n132, A2 => n127, ZN => n135);
   U43 : NAND2_X1 port map( A1 => n145, A2 => n144, ZN => n131);
   U44 : INV_X1 port map( A => a(14), ZN => n145);
   U45 : INV_X1 port map( A => b(14), ZN => n144);
   U46 : NAND2_X1 port map( A1 => n161, A2 => n162, ZN => net138780);
   U47 : INV_X1 port map( A => n170, ZN => n162);
   U48 : CLKBUF_X1 port map( A => n184, Z => n104);
   U49 : CLKBUF_X1 port map( A => n164, Z => n105);
   U50 : AND2_X1 port map( A1 => net139124, A2 => n131, ZN => n106);
   U51 : AND2_X1 port map( A1 => n170, A2 => net150681, ZN => n107);
   U52 : AND2_X1 port map( A1 => a(19), A2 => b(19), ZN => n108);
   U53 : INV_X1 port map( A => b(27), ZN => n199);
   U54 : INV_X1 port map( A => a(27), ZN => n198);
   U55 : OAI222_X1 port map( A1 => n206, A2 => a(12), B1 => n227, B2 => b(12), 
                           C1 => b(13), C2 => a(13), ZN => n109);
   U56 : NAND2_X1 port map( A1 => n228, A2 => n203, ZN => n110);
   U57 : NAND2_X1 port map( A1 => n120, A2 => net138989, ZN => n61);
   U58 : NAND3_X1 port map( A1 => n139, A2 => n149, A3 => n151, ZN => n113);
   U59 : NAND2_X1 port map( A1 => n150, A2 => n146, ZN => n149);
   U60 : NAND2_X1 port map( A1 => a(15), A2 => n106, ZN => net153886);
   U61 : NAND2_X1 port map( A1 => n118, A2 => a(20), ZN => n142);
   U62 : AOI21_X1 port map( B1 => n110, B2 => n131, A => a(15), ZN => n130);
   U63 : NOR2_X1 port map( A1 => n130, A2 => n137, ZN => n139);
   U64 : NAND2_X1 port map( A1 => n113, A2 => n119, ZN => n118);
   U65 : INV_X1 port map( A => n153, ZN => net151348);
   U66 : AOI21_X1 port map( B1 => n135, B2 => n140, A => n108, ZN => n119);
   U67 : AND2_X2 port map( A1 => n113, A2 => n119, ZN => n153);
   U68 : AOI21_X1 port map( B1 => n142, B2 => n143, A => n134, ZN => n141);
   U69 : NAND2_X1 port map( A1 => n141, A2 => n152, ZN => n120);
   U70 : BUF_X1 port map( A => b(0), Z => n208);
   U71 : AND2_X1 port map( A1 => b(0), A2 => a(0), ZN => n154);
   U72 : OAI22_X1 port map( A1 => a(7), A2 => b(7), B1 => a(6), B2 => b(6), ZN 
                           => n170);
   U73 : INV_X1 port map( A => b(7), ZN => n103);
   U74 : OAI211_X1 port map( C1 => a(1), C2 => b(1), A => n182, B => n183, ZN 
                           => n155);
   U75 : AND4_X1 port map( A1 => n174, A2 => n179, A3 => n180, A4 => a(3), ZN 
                           => n158);
   U76 : INV_X1 port map( A => b(2), ZN => n176);
   U77 : OAI22_X1 port map( A1 => n208, A2 => a(0), B1 => n214, B2 => cin, ZN 
                           => n156);
   U78 : AND2_X1 port map( A1 => net138777, A2 => net139158, ZN => n157);
   U79 : NOR2_X1 port map( A1 => n166, A2 => n157, ZN => n167);
   U80 : OAI21_X1 port map( B1 => n158, B2 => b(3), A => n159, ZN => net138777)
                           ;
   U81 : OAI21_X1 port map( B1 => n167, B2 => n172, A => n181, ZN => n164);
   U82 : NAND2_X1 port map( A1 => n156, A2 => n173, ZN => n182);
   U83 : INV_X1 port map( A => b(1), ZN => n177);
   U84 : NAND2_X1 port map( A1 => n184, A2 => n165, ZN => n159);
   U85 : INV_X1 port map( A => n104, ZN => net151886);
   U86 : NAND2_X1 port map( A1 => n175, A2 => n178, ZN => n179);
   U87 : NOR2_X1 port map( A1 => n111, A2 => b(4), ZN => n166);
   U88 : NAND2_X1 port map( A1 => n155, A2 => n176, ZN => n174);
   U89 : OAI211_X1 port map( C1 => a(1), C2 => b(1), A => n183, B => n182, ZN 
                           => n175);
   U90 : NAND2_X1 port map( A1 => n121, A2 => n177, ZN => n183);
   U91 : NAND2_X1 port map( A1 => n187, A2 => n105, ZN => n161);
   U92 : AOI21_X1 port map( B1 => n164, B2 => n171, A => n107, ZN => n252);
   U93 : AOI21_X1 port map( B1 => n164, B2 => n163, A => n107, ZN => n188);
   U94 : BUF_X1 port map( A => n250, Z => cout_5_port);
   U95 : OAI21_X1 port map( B1 => a(23), B2 => n230, A => b(23), ZN => n189);
   U96 : NOR2_X1 port map( A1 => n190, A2 => a(24), ZN => n193);
   U97 : NOR2_X1 port map( A1 => n191, A2 => n231, ZN => n190);
   U98 : OAI22_X1 port map( A1 => a(22), A2 => net139150, B1 => b(22), B2 => 
                           n229, ZN => n191);
   U99 : OR2_X1 port map( A1 => n191, A2 => n231, ZN => n192);
   U100 : CLKBUF_X1 port map( A => n206, Z => cout_2_port);
   U101 : NAND2_X1 port map( A1 => n209, A2 => n192, ZN => n250);
   U102 : CLKBUF_X1 port map( A => n158, Z => net151510);
   U103 : OAI22_X1 port map( A1 => n198, A2 => n199, B1 => n239, B2 => n200, ZN
                           => cout_6_port);
   U104 : OR2_X1 port map( A1 => a(11), A2 => b(11), ZN => n196);
   U105 : NAND2_X1 port map( A1 => n225, A2 => n196, ZN => n226);
   U106 : NOR2_X1 port map( A1 => a(27), A2 => b(27), ZN => n200);
   U107 : AND2_X1 port map( A1 => b(9), A2 => a(9), ZN => n201);
   U108 : NOR2_X1 port map( A1 => n220, A2 => n201, ZN => n224);
   U109 : OAI22_X1 port map( A1 => a(22), A2 => net139150, B1 => n229, B2 => 
                           b(22), ZN => n202);
   U110 : OR2_X1 port map( A1 => n102, A2 => n103, ZN => net150681);
   U111 : INV_X1 port map( A => b(25), ZN => n233);
   U112 : OAI21_X1 port map( B1 => n249, B2 => n248, A => n247, ZN => 
                           cout_7_port);
   U113 : INV_X1 port map( A => b(29), ZN => n242);
   U114 : INV_X1 port map( A => a(10), ZN => n222);
   U115 : INV_X1 port map( A => b(10), ZN => n221);
   U116 : INV_X1 port map( A => a(5), ZN => net138600);
   U117 : OR2_X1 port map( A1 => a(26), A2 => b(26), ZN => n238);
   U118 : INV_X1 port map( A => a(25), ZN => n234);
   U119 : INV_X1 port map( A => a(9), ZN => n217);
   U120 : INV_X1 port map( A => b(9), ZN => n216);
   U121 : AND2_X1 port map( A1 => n205, A2 => n204, ZN => n203);
   U122 : NOR2_X1 port map( A1 => b(10), A2 => a(10), ZN => n223);
   U123 : NOR2_X1 port map( A1 => b(25), A2 => a(25), ZN => n235);
   U124 : NAND2_X1 port map( A1 => a(11), A2 => b(11), ZN => n212);
   U125 : NAND2_X1 port map( A1 => a(14), A2 => b(14), ZN => n204);
   U126 : NAND2_X1 port map( A1 => a(13), A2 => b(13), ZN => n205);
   U127 : OAI22_X1 port map( A1 => a(30), A2 => n245, B1 => b(30), B2 => n244, 
                           ZN => n249);
   U128 : AND2_X1 port map( A1 => n245, A2 => a(30), ZN => n244);
   U129 : OAI21_X1 port map( B1 => n243, B2 => n242, A => n241, ZN => n245);
   U130 : OAI222_X1 port map( A1 => a(28), A2 => n211, B1 => b(28), B2 => n240,
                           C1 => b(29), C2 => a(29), ZN => n241);
   U131 : OAI21_X1 port map( B1 => n246, B2 => a(31), A => b(31), ZN => n247);
   U132 : INV_X1 port map( A => n249, ZN => n246);
   U133 : INV_X1 port map( A => a(31), ZN => n248);
   U134 : INV_X1 port map( A => a(29), ZN => n243);
   U135 : INV_X1 port map( A => a(4), ZN => net139158);
   U136 : NOR2_X1 port map( A1 => net138777, A2 => net139158, ZN => n111);
   U137 : CLKBUF_X1 port map( A => n61, Z => net139150);
   U138 : NAND2_X1 port map( A1 => n109, A2 => n203, ZN => net139124);
   U139 : NAND2_X1 port map( A1 => n226, A2 => n212, ZN => n206);
   U140 : NAND2_X1 port map( A1 => n226, A2 => n212, ZN => n251);
   U141 : OR2_X1 port map( A1 => n63, A2 => n64, ZN => net138989);
   U142 : OAI21_X1 port map( B1 => a(15), B2 => n106, A => b(15), ZN => n207);
   U143 : OAI21_X1 port map( B1 => n230, B2 => a(23), A => b(23), ZN => n209);
   U144 : NAND2_X1 port map( A1 => net153886, A2 => n207, ZN => cout_3_port);
   U145 : NAND2_X1 port map( A1 => n193, A2 => n189, ZN => n232);
   U146 : OAI22_X1 port map( A1 => n224, A2 => n223, B1 => n222, B2 => n221, ZN
                           => n225);
   U147 : AOI22_X1 port map( A1 => n218, A2 => n219, B1 => n217, B2 => n216, ZN
                           => n220);
   U148 : AND2_X1 port map( A1 => n61, A2 => a(22), ZN => n229);
   U149 : INV_X1 port map( A => n202, ZN => n230);
   U150 : CLKBUF_X1 port map( A => cout_6_port, Z => n211);
   U151 : OAI21_X1 port map( B1 => n102, B2 => n103, A => net138780, ZN => 
                           cout_1_port);
   U152 : OAI222_X1 port map( A1 => n206, A2 => a(12), B1 => n227, B2 => b(12),
                           C1 => b(13), C2 => a(13), ZN => n228);
   U153 : OAI22_X1 port map( A1 => n208, A2 => a(0), B1 => n154, B2 => cin, ZN 
                           => n121);
   U154 : AND2_X1 port map( A1 => b(0), A2 => a(0), ZN => n214);
   U155 : INV_X1 port map( A => a(23), ZN => n231);
   U156 : AND2_X1 port map( A1 => n211, A2 => a(28), ZN => n240);
   U157 : AOI22_X1 port map( A1 => b(26), A2 => a(26), B1 => n237, B2 => n238, 
                           ZN => n239);
   U158 : NAND2_X1 port map( A1 => n188, A2 => a(8), ZN => n219);
   U159 : OAI22_X1 port map( A1 => n236, A2 => n235, B1 => n234, B2 => n233, ZN
                           => n237);
   U160 : AND2_X1 port map( A1 => n251, A2 => a(12), ZN => n227);
   U161 : OAI21_X1 port map( B1 => n252, B2 => a(8), A => b(8), ZN => n218);
   U162 : AOI22_X1 port map( A1 => n232, A2 => b(24), B1 => n250, B2 => a(24), 
                           ZN => n236);
   U163 : INV_X1 port map( A => n215, ZN => cout_0_port);
   U164 : OAI22_X1 port map( A1 => a(3), A2 => net151886, B1 => b(3), B2 => 
                           net151510, ZN => n215);

end SYN_p4_carry_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4CarryGenerator_DATA_SIZE32_SPARSITY4_6 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  cout :
         out std_logic_vector (7 downto 0));

end P4CarryGenerator_DATA_SIZE32_SPARSITY4_6;

architecture SYN_p4_carry_generator_arch of 
   P4CarryGenerator_DATA_SIZE32_SPARSITY4_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal cout_7_port, n246, n247, cout_2_port, n248, cout_0_port, n40, n42, 
      n43, n59, n69, n78, n79, n80, n103, net134390, net150386, net150417, 
      net150559, net151260, net151344, net151394, net151393, net151449, 
      net151838, net152641, net152651, net153832, n102, n104, n105, n106, n107,
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, 
      n120, n121, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205, n206, cout_5_port, n208, n209, n210, n211, n212, n213, n214, n215, 
      n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
      n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, 
      n240, n241, n242, n243, n244, n245 : std_logic;

begin
   cout <= ( cout_7_port, net151260, cout_5_port, net151394, net150417, 
      cout_2_port, net150386, cout_0_port );
   
   syn164 : NAND3_X1 port map( A1 => n247, A2 => n136, A3 => n133, ZN => n118);
   net154186 : NAND3_X1 port map( A1 => a(16), A2 => n79, A3 => b(16), ZN => 
                           n78);
   U1 : NAND2_X1 port map( A1 => n129, A2 => n130, ZN => n135);
   U2 : INV_X1 port map( A => a(21), ZN => n129);
   U3 : NOR2_X1 port map( A1 => a(7), A2 => b(7), ZN => n184);
   U4 : NAND2_X1 port map( A1 => n176, A2 => n177, ZN => n174);
   U5 : INV_X1 port map( A => b(6), ZN => n189);
   U6 : INV_X1 port map( A => b(16), ZN => n131);
   U7 : INV_X1 port map( A => n79, ZN => n126);
   U8 : INV_X1 port map( A => b(3), ZN => n188);
   U9 : INV_X1 port map( A => b(21), ZN => n130);
   U10 : NAND2_X1 port map( A1 => a(5), A2 => b(5), ZN => n185);
   U11 : INV_X1 port map( A => b(4), ZN => n182);
   U12 : INV_X1 port map( A => a(4), ZN => n181);
   U13 : INV_X1 port map( A => b(5), ZN => n176);
   U14 : INV_X1 port map( A => a(5), ZN => n177);
   U15 : NAND2_X1 port map( A1 => b(21), A2 => a(21), ZN => n123);
   U16 : INV_X1 port map( A => b(2), ZN => n187);
   U17 : INV_X1 port map( A => a(16), ZN => n132);
   U18 : INV_X1 port map( A => a(6), ZN => n183);
   U19 : INV_X1 port map( A => a(7), ZN => net134390);
   U20 : INV_X1 port map( A => b(7), ZN => n103);
   U21 : NOR2_X1 port map( A1 => n126, A2 => n134, ZN => n133);
   U22 : NAND2_X1 port map( A1 => n131, A2 => n132, ZN => n136);
   U23 : OAI22_X1 port map( A1 => b(19), A2 => a(19), B1 => b(18), B2 => a(18),
                           ZN => n134);
   U24 : NOR2_X1 port map( A1 => n128, A2 => n109, ZN => n117);
   U25 : NOR2_X1 port map( A1 => n69, A2 => n127, ZN => n128);
   U26 : NOR2_X1 port map( A1 => a(19), A2 => b(19), ZN => n127);
   U27 : INV_X1 port map( A => a(3), ZN => n180);
   U28 : CLKBUF_X1 port map( A => n105, Z => n102);
   U29 : AOI22_X1 port map( A1 => n146, A2 => b(24), B1 => n246, B2 => a(24), 
                           ZN => n104);
   U30 : NAND2_X1 port map( A1 => n117, A2 => n118, ZN => n105);
   U31 : AOI21_X1 port map( B1 => n105, B2 => a(20), A => b(20), ZN => n120);
   U32 : AOI22_X1 port map( A1 => n146, A2 => b(24), B1 => n246, B2 => a(24), 
                           ZN => n106);
   U33 : OAI22_X1 port map( A1 => n208, A2 => a(0), B1 => n225, B2 => cin, ZN 
                           => n107);
   U34 : OR2_X1 port map( A1 => n108, A2 => b(1), ZN => n160);
   U35 : NOR2_X1 port map( A1 => n107, A2 => n178, ZN => n108);
   U36 : AND2_X1 port map( A1 => b(19), A2 => a(19), ZN => n109);
   U37 : AND2_X1 port map( A1 => n196, A2 => n197, ZN => n110);
   U38 : NOR2_X1 port map( A1 => a(27), A2 => b(27), ZN => n111);
   U39 : INV_X1 port map( A => a(2), ZN => n179);
   U40 : INV_X1 port map( A => a(1), ZN => n178);
   U41 : INV_X1 port map( A => a(15), ZN => n138);
   U42 : AND2_X1 port map( A1 => n138, A2 => n112, ZN => n114);
   U43 : NAND2_X1 port map( A1 => n215, A2 => n211, ZN => n112);
   U44 : OR2_X1 port map( A1 => n114, A2 => n115, ZN => n113);
   U45 : NAND2_X1 port map( A1 => n113, A2 => n116, ZN => n247);
   U46 : INV_X1 port map( A => b(15), ZN => n115);
   U47 : OR2_X1 port map( A1 => n138, A2 => n80, ZN => n116);
   U48 : OAI21_X1 port map( B1 => net152641, B2 => a(20), A => n135, ZN => n121
                           );
   U49 : OAI21_X1 port map( B1 => n120, B2 => n121, A => n123, ZN => n119);
   U50 : OAI21_X1 port map( B1 => n120, B2 => n121, A => n123, ZN => n137);
   U51 : NAND2_X1 port map( A1 => n117, A2 => n118, ZN => net152641);
   U52 : OAI21_X1 port map( B1 => n119, B2 => a(22), A => b(22), ZN => n125);
   U53 : NAND2_X1 port map( A1 => n137, A2 => a(22), ZN => n124);
   U54 : NAND2_X1 port map( A1 => n125, A2 => n124, ZN => net153832);
   U55 : AND2_X1 port map( A1 => n125, A2 => n124, ZN => net151838);
   U56 : OAI222_X1 port map( A1 => net151260, A2 => a(28), B1 => b(28), B2 => 
                           n140, C1 => b(29), C2 => a(29), ZN => n139);
   U57 : NAND2_X1 port map( A1 => n139, A2 => net150559, ZN => n40);
   U58 : NAND2_X1 port map( A1 => n154, A2 => n155, ZN => n140);
   U59 : NAND2_X1 port map( A1 => a(28), A2 => n150, ZN => n155);
   U60 : INV_X1 port map( A => a(28), ZN => n153);
   U61 : OR2_X1 port map( A1 => n111, A2 => n153, ZN => n152);
   U62 : OR2_X1 port map( A1 => n152, A2 => n156, ZN => n154);
   U63 : AOI22_X1 port map( A1 => b(26), A2 => a(26), B1 => n158, B2 => n142, 
                           ZN => n156);
   U64 : OAI22_X1 port map( A1 => n144, A2 => n104, B1 => n147, B2 => n145, ZN 
                           => n158);
   U65 : INV_X1 port map( A => b(25), ZN => n145);
   U66 : OAI22_X1 port map( A1 => n106, A2 => n144, B1 => n147, B2 => n145, ZN 
                           => n143);
   U67 : INV_X1 port map( A => a(25), ZN => n147);
   U68 : NOR2_X1 port map( A1 => n141, A2 => n111, ZN => n151);
   U69 : OR2_X2 port map( A1 => n151, A2 => n150, ZN => net151260);
   U70 : AOI22_X1 port map( A1 => b(26), A2 => a(26), B1 => n142, B2 => n143, 
                           ZN => n141);
   U71 : INV_X1 port map( A => b(29), ZN => n43);
   U72 : INV_X1 port map( A => a(29), ZN => n42);
   U73 : NOR2_X1 port map( A1 => n148, A2 => n149, ZN => n150);
   U74 : INV_X1 port map( A => b(27), ZN => n149);
   U75 : INV_X1 port map( A => a(27), ZN => n148);
   U76 : OR2_X1 port map( A1 => a(26), A2 => b(26), ZN => n142);
   U77 : NOR2_X1 port map( A1 => b(25), A2 => a(25), ZN => n144);
   U78 : NAND2_X1 port map( A1 => n157, A2 => n59, ZN => n146);
   U79 : NOR2_X1 port map( A1 => net152651, A2 => a(24), ZN => n157);
   U80 : NAND2_X1 port map( A1 => n160, A2 => n159, ZN => n190);
   U81 : AND2_X1 port map( A1 => n164, A2 => a(2), ZN => n159);
   U82 : NAND2_X1 port map( A1 => n107, A2 => n178, ZN => n164);
   U83 : NAND2_X1 port map( A1 => n160, A2 => n164, ZN => n163);
   U84 : NAND2_X1 port map( A1 => n163, A2 => n179, ZN => n166);
   U85 : CLKBUF_X1 port map( A => n168, Z => n161);
   U86 : NAND2_X1 port map( A1 => n165, A2 => n180, ZN => n169);
   U87 : NAND2_X1 port map( A1 => n175, A2 => net151449, ZN => n162);
   U88 : INV_X1 port map( A => n161, ZN => cout_0_port);
   U89 : NAND2_X1 port map( A1 => n170, A2 => n169, ZN => n168);
   U90 : OAI21_X1 port map( B1 => n165, B2 => n180, A => n188, ZN => n170);
   U91 : NAND2_X1 port map( A1 => n166, A2 => n167, ZN => n165);
   U92 : NAND2_X1 port map( A1 => n175, A2 => net151449, ZN => n248);
   U93 : NAND2_X1 port map( A1 => n190, A2 => n187, ZN => n167);
   U94 : NAND2_X1 port map( A1 => n191, A2 => n186, ZN => n175);
   U95 : OAI21_X1 port map( B1 => n172, B2 => n173, A => n174, ZN => n171);
   U96 : OAI21_X1 port map( B1 => n171, B2 => n183, A => n189, ZN => n191);
   U97 : AOI21_X1 port map( B1 => n171, B2 => n183, A => n184, ZN => n186);
   U98 : OAI21_X1 port map( B1 => n168, B2 => n181, A => n185, ZN => n173);
   U99 : AOI21_X1 port map( B1 => n168, B2 => n181, A => n182, ZN => n172);
   U100 : NOR2_X1 port map( A1 => net151838, A2 => n223, ZN => net152651);
   U101 : OR2_X1 port map( A1 => net151838, A2 => n223, ZN => n192);
   U102 : OAI21_X1 port map( B1 => net153832, B2 => a(23), A => b(23), ZN => 
                           n193);
   U103 : AND2_X1 port map( A1 => n59, A2 => n192, ZN => n194);
   U104 : NAND2_X1 port map( A1 => n236, A2 => n110, ZN => n215);
   U105 : OAI22_X1 port map( A1 => a(30), A2 => net151344, B1 => n242, B2 => 
                           b(30), ZN => n195);
   U106 : OR2_X1 port map( A1 => net134390, A2 => n103, ZN => net151449);
   U107 : NAND2_X1 port map( A1 => n193, A2 => n192, ZN => n246);
   U108 : OR2_X1 port map( A1 => n216, A2 => n217, ZN => n196);
   U109 : OR2_X1 port map( A1 => n218, A2 => n219, ZN => n197);
   U110 : INV_X1 port map( A => n102, ZN => net151393);
   U111 : INV_X1 port map( A => net151393, ZN => net151394);
   U112 : CLKBUF_X1 port map( A => n40, Z => net151344);
   U113 : CLKBUF_X1 port map( A => n234, Z => n198);
   U114 : NAND2_X1 port map( A1 => n234, A2 => n201, ZN => n199);
   U115 : AND2_X1 port map( A1 => n199, A2 => n200, ZN => n213);
   U116 : OR2_X1 port map( A1 => b(12), A2 => a(12), ZN => n200);
   U117 : AND2_X1 port map( A1 => n206, A2 => n210, ZN => n201);
   U118 : NAND2_X1 port map( A1 => n202, A2 => n206, ZN => n212);
   U119 : AND2_X1 port map( A1 => n234, A2 => n203, ZN => n202);
   U120 : INV_X1 port map( A => a(12), ZN => n203);
   U121 : OR2_X1 port map( A1 => a(11), A2 => b(11), ZN => n204);
   U122 : NAND2_X1 port map( A1 => n233, A2 => n204, ZN => n234);
   U123 : OR2_X1 port map( A1 => n42, A2 => n43, ZN => net150559);
   U124 : OR2_X1 port map( A1 => n245, A2 => n224, ZN => n205);
   U125 : NAND2_X1 port map( A1 => n244, A2 => n205, ZN => cout_7_port);
   U126 : OR2_X1 port map( A1 => n222, A2 => n235, ZN => n206);
   U127 : NAND2_X1 port map( A1 => n206, A2 => n198, ZN => cout_2_port);
   U128 : CLKBUF_X1 port map( A => n247, Z => net150417);
   U129 : INV_X1 port map( A => n194, ZN => cout_5_port);
   U130 : CLKBUF_X1 port map( A => n162, Z => net150386);
   U131 : INV_X1 port map( A => b(14), ZN => n217);
   U132 : INV_X1 port map( A => b(12), ZN => n210);
   U133 : INV_X1 port map( A => b(10), ZN => n230);
   U134 : NOR2_X1 port map( A1 => b(10), A2 => a(10), ZN => n231);
   U135 : INV_X1 port map( A => b(17), ZN => n237);
   U136 : INV_X1 port map( A => a(14), ZN => n216);
   U137 : INV_X1 port map( A => a(13), ZN => n218);
   U138 : INV_X1 port map( A => b(13), ZN => n219);
   U139 : INV_X1 port map( A => b(11), ZN => n235);
   U140 : NAND2_X1 port map( A1 => n237, A2 => n238, ZN => n79);
   U141 : OAI21_X1 port map( B1 => a(18), B2 => n241, A => n240, ZN => n69);
   U142 : INV_X1 port map( A => n239, ZN => n240);
   U143 : AOI21_X1 port map( B1 => n241, B2 => a(18), A => b(18), ZN => n239);
   U144 : OAI21_X1 port map( B1 => n238, B2 => n237, A => n78, ZN => n241);
   U145 : INV_X1 port map( A => a(17), ZN => n238);
   U146 : CLKBUF_X1 port map( A => b(0), Z => n208);
   U147 : AND2_X1 port map( A1 => b(9), A2 => a(9), ZN => n209);
   U148 : NOR2_X1 port map( A1 => n229, A2 => n209, ZN => n232);
   U149 : INV_X1 port map( A => b(9), ZN => n226);
   U150 : OAI22_X1 port map( A1 => n232, A2 => n231, B1 => n221, B2 => n230, ZN
                           => n233);
   U151 : OR2_X1 port map( A1 => b(14), A2 => a(14), ZN => n211);
   U152 : NAND2_X1 port map( A1 => n215, A2 => n211, ZN => n80);
   U153 : OR2_X1 port map( A1 => b(13), A2 => a(13), ZN => n214);
   U154 : NAND3_X1 port map( A1 => n212, A2 => n213, A3 => n214, ZN => n236);
   U155 : AOI22_X1 port map( A1 => n228, A2 => n227, B1 => n220, B2 => n226, ZN
                           => n229);
   U156 : OAI21_X1 port map( B1 => n243, B2 => a(31), A => b(31), ZN => n244);
   U157 : NAND2_X1 port map( A1 => n162, A2 => a(8), ZN => n228);
   U158 : OAI22_X1 port map( A1 => a(30), A2 => net151344, B1 => b(30), B2 => 
                           n242, ZN => n245);
   U159 : OAI21_X1 port map( B1 => net153832, B2 => a(23), A => b(23), ZN => 
                           n59);
   U160 : AND2_X1 port map( A1 => n40, A2 => a(30), ZN => n242);
   U161 : INV_X1 port map( A => n195, ZN => n243);
   U162 : AND2_X1 port map( A1 => b(0), A2 => a(0), ZN => n225);
   U163 : OAI21_X1 port map( B1 => n248, B2 => a(8), A => b(8), ZN => n227);
   U164 : INV_X1 port map( A => a(9), ZN => n220);
   U165 : INV_X1 port map( A => a(10), ZN => n221);
   U166 : INV_X1 port map( A => a(11), ZN => n222);
   U167 : INV_X1 port map( A => a(23), ZN => n223);
   U168 : INV_X1 port map( A => a(31), ZN => n224);

end SYN_p4_carry_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4CarryGenerator_DATA_SIZE32_SPARSITY4_5 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  cout :
         out std_logic_vector (7 downto 0));

end P4CarryGenerator_DATA_SIZE32_SPARSITY4_5;

architecture SYN_p4_carry_generator_arch of 
   P4CarryGenerator_DATA_SIZE32_SPARSITY4_5 is

   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI221_X4
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal cout_7_port, n232, cout_4_port, n233, cout_2_port, n234, n235, 
      cout_5_port, cout_1_port, n125, cout_3_port, cout_0_port, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, cout_6_port, 
      n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, 
      n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, 
      n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, 
      n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, 
      n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, 
      n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, 
      n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, 
      n225, n226, n227, n228, n229, n230, n231 : std_logic;

begin
   cout <= ( cout_7_port, cout_6_port, cout_5_port, cout_4_port, cout_3_port, 
      cout_2_port, cout_1_port, cout_0_port );
   
   U95 : NAND3_X1 port map( A1 => a(16), A2 => n191, A3 => b(16), ZN => n192);
   U1 : OR2_X1 port map( A1 => n147, A2 => n148, ZN => n143);
   U2 : OR2_X1 port map( A1 => n149, A2 => n150, ZN => n144);
   U3 : OAI222_X1 port map( A1 => a(28), A2 => n125, B1 => b(28), B2 => n222, 
                           C1 => b(29), C2 => a(29), ZN => n223);
   U4 : CLKBUF_X1 port map( A => n232, Z => cout_5_port);
   U5 : CLKBUF_X1 port map( A => n234, Z => cout_1_port);
   U6 : CLKBUF_X1 port map( A => cout_6_port, Z => n125);
   U7 : OAI22_X1 port map( A1 => n141, A2 => n142, B1 => n132, B2 => n221, ZN 
                           => cout_6_port);
   U8 : CLKBUF_X1 port map( A => n233, Z => cout_3_port);
   U9 : CLKBUF_X1 port map( A => n235, Z => cout_0_port);
   U10 : NAND2_X1 port map( A1 => n136, A2 => n128, ZN => n214);
   U11 : AND2_X1 port map( A1 => n211, A2 => n129, ZN => n128);
   U12 : INV_X1 port map( A => a(24), ZN => n129);
   U13 : OR2_X1 port map( A1 => a(11), A2 => b(11), ZN => n130);
   U14 : NAND2_X1 port map( A1 => n130, A2 => n181, ZN => n182);
   U15 : NAND2_X1 port map( A1 => n145, A2 => n182, ZN => cout_2_port);
   U16 : OR2_X1 port map( A1 => n171, A2 => n170, ZN => n131);
   U17 : NAND2_X1 port map( A1 => n131, A2 => n169, ZN => n234);
   U18 : OAI221_X4 port map( B1 => n203, B2 => n202, C1 => n201, C2 => n200, A 
                           => n199, ZN => cout_4_port);
   U19 : NOR2_X1 port map( A1 => a(27), A2 => b(27), ZN => n132);
   U20 : INV_X1 port map( A => b(27), ZN => n142);
   U21 : INV_X1 port map( A => a(27), ZN => n141);
   U22 : CLKBUF_X1 port map( A => n168, Z => n133);
   U23 : CLKBUF_X1 port map( A => a(0), Z => n134);
   U24 : AND2_X1 port map( A1 => b(9), A2 => a(9), ZN => n135);
   U25 : NOR2_X1 port map( A1 => n176, A2 => n135, ZN => n180);
   U26 : OR2_X1 port map( A1 => n213, A2 => n212, ZN => n136);
   U27 : NAND2_X1 port map( A1 => n136, A2 => n211, ZN => n232);
   U28 : OR2_X1 port map( A1 => n190, A2 => n189, ZN => n137);
   U29 : NAND2_X1 port map( A1 => n137, A2 => n188, ZN => n233);
   U30 : OR2_X1 port map( A1 => b(14), A2 => a(14), ZN => n138);
   U31 : NAND2_X1 port map( A1 => n146, A2 => n138, ZN => n190);
   U32 : OR2_X1 port map( A1 => n207, A2 => n206, ZN => n139);
   U33 : NAND2_X1 port map( A1 => n139, A2 => n205, ZN => n209);
   U34 : NAND3_X1 port map( A1 => n186, A2 => n144, A3 => n143, ZN => n146);
   U35 : OR2_X1 port map( A1 => n184, A2 => n183, ZN => n145);
   U36 : INV_X1 port map( A => a(14), ZN => n147);
   U37 : INV_X1 port map( A => b(14), ZN => n148);
   U38 : INV_X1 port map( A => a(13), ZN => n149);
   U39 : INV_X1 port map( A => b(13), ZN => n150);
   U40 : OAI222_X1 port map( A1 => a(12), A2 => cout_2_port, B1 => b(12), B2 =>
                           n185, C1 => b(13), C2 => a(13), ZN => n186);
   U41 : INV_X1 port map( A => n201, ZN => n198);
   U42 : NAND2_X1 port map( A1 => n193, A2 => n194, ZN => n191);
   U43 : OAI21_X1 port map( B1 => n231, B2 => n230, A => n229, ZN => 
                           cout_7_port);
   U44 : INV_X1 port map( A => b(7), ZN => n170);
   U45 : INV_X1 port map( A => a(7), ZN => n171);
   U46 : INV_X1 port map( A => a(23), ZN => n212);
   U47 : INV_X1 port map( A => n213, ZN => n210);
   U48 : INV_X1 port map( A => a(15), ZN => n189);
   U49 : INV_X1 port map( A => n190, ZN => n187);
   U50 : OAI22_X1 port map( A1 => a(4), A2 => n235, B1 => b(4), B2 => n162, ZN 
                           => n163);
   U51 : AND2_X1 port map( A1 => n235, A2 => a(4), ZN => n162);
   U52 : OAI22_X1 port map( A1 => a(2), A2 => n157, B1 => b(2), B2 => n156, ZN 
                           => n158);
   U53 : AND2_X1 port map( A1 => n157, A2 => a(2), ZN => n156);
   U54 : INV_X1 port map( A => n155, ZN => n157);
   U55 : OAI22_X1 port map( A1 => a(1), A2 => n154, B1 => b(1), B2 => n153, ZN 
                           => n155);
   U56 : INV_X1 port map( A => b(11), ZN => n183);
   U57 : INV_X1 port map( A => a(11), ZN => n184);
   U58 : OAI21_X1 port map( B1 => a(18), B2 => n197, A => n196, ZN => n201);
   U59 : INV_X1 port map( A => n195, ZN => n196);
   U60 : AOI21_X1 port map( B1 => n197, B2 => a(18), A => b(18), ZN => n195);
   U61 : OAI21_X1 port map( B1 => n194, B2 => n193, A => n192, ZN => n197);
   U62 : AOI22_X1 port map( A1 => b(26), A2 => a(26), B1 => n219, B2 => n220, 
                           ZN => n221);
   U63 : OR2_X1 port map( A1 => a(26), A2 => b(26), ZN => n220);
   U64 : INV_X1 port map( A => b(25), ZN => n215);
   U65 : OAI22_X1 port map( A1 => n180, A2 => n179, B1 => n178, B2 => n177, ZN 
                           => n181);
   U66 : INV_X1 port map( A => b(10), ZN => n177);
   U67 : INV_X1 port map( A => a(10), ZN => n178);
   U68 : NOR2_X1 port map( A1 => b(10), A2 => a(10), ZN => n179);
   U69 : AOI22_X1 port map( A1 => n174, A2 => n175, B1 => n173, B2 => n172, ZN 
                           => n176);
   U70 : INV_X1 port map( A => b(9), ZN => n172);
   U71 : INV_X1 port map( A => a(9), ZN => n173);
   U72 : OAI22_X1 port map( A1 => a(22), A2 => n209, B1 => b(22), B2 => n208, 
                           ZN => n213);
   U73 : AND2_X1 port map( A1 => n209, A2 => a(22), ZN => n208);
   U74 : INV_X1 port map( A => b(21), ZN => n206);
   U75 : OAI21_X1 port map( B1 => n234, B2 => a(8), A => b(8), ZN => n174);
   U76 : NAND2_X1 port map( A1 => a(8), A2 => n234, ZN => n175);
   U77 : INV_X1 port map( A => a(17), ZN => n194);
   U78 : INV_X1 port map( A => a(19), ZN => n200);
   U79 : OAI22_X1 port map( A1 => b(19), A2 => a(19), B1 => b(18), B2 => a(18),
                           ZN => n202);
   U80 : OAI21_X1 port map( B1 => n198, B2 => a(19), A => b(19), ZN => n199);
   U81 : INV_X1 port map( A => b(17), ZN => n193);
   U82 : INV_X1 port map( A => n166, ZN => n168);
   U83 : OAI22_X1 port map( A1 => a(5), A2 => n165, B1 => b(5), B2 => n164, ZN 
                           => n166);
   U84 : AND2_X1 port map( A1 => n165, A2 => a(5), ZN => n164);
   U85 : INV_X1 port map( A => n163, ZN => n165);
   U86 : INV_X1 port map( A => n152, ZN => n154);
   U87 : OAI22_X1 port map( A1 => b(0), A2 => n134, B1 => cin, B2 => n151, ZN 
                           => n152);
   U88 : AND2_X1 port map( A1 => a(0), A2 => b(0), ZN => n151);
   U89 : AND2_X1 port map( A1 => n154, A2 => a(1), ZN => n153);
   U90 : OAI222_X1 port map( A1 => a(20), A2 => cout_4_port, B1 => b(20), B2 =>
                           n204, C1 => b(21), C2 => a(21), ZN => n205);
   U91 : AND2_X1 port map( A1 => cout_4_port, A2 => a(20), ZN => n204);
   U92 : INV_X1 port map( A => n161, ZN => n235);
   U93 : AND2_X1 port map( A1 => n160, A2 => a(3), ZN => n159);
   U94 : INV_X1 port map( A => n158, ZN => n160);
   U96 : NOR2_X1 port map( A1 => b(25), A2 => a(25), ZN => n217);
   U97 : INV_X1 port map( A => a(21), ZN => n207);
   U98 : INV_X1 port map( A => a(25), ZN => n216);
   U99 : AND2_X1 port map( A1 => n125, A2 => a(28), ZN => n222);
   U100 : OAI22_X1 port map( A1 => a(30), A2 => n227, B1 => b(30), B2 => n226, 
                           ZN => n231);
   U101 : AND2_X1 port map( A1 => n227, A2 => a(30), ZN => n226);
   U102 : OAI21_X1 port map( B1 => n225, B2 => n224, A => n223, ZN => n227);
   U103 : INV_X1 port map( A => a(29), ZN => n225);
   U104 : OAI21_X1 port map( B1 => n228, B2 => a(31), A => b(31), ZN => n229);
   U105 : INV_X1 port map( A => n231, ZN => n228);
   U106 : INV_X1 port map( A => b(29), ZN => n224);
   U107 : INV_X1 port map( A => a(31), ZN => n230);
   U108 : OAI22_X1 port map( A1 => n218, A2 => n217, B1 => n216, B2 => n215, ZN
                           => n219);
   U109 : AOI22_X1 port map( A1 => b(24), A2 => n214, B1 => a(24), B2 => n232, 
                           ZN => n218);
   U110 : OAI22_X1 port map( A1 => a(3), A2 => n160, B1 => b(3), B2 => n159, ZN
                           => n161);
   U111 : OAI222_X1 port map( A1 => a(6), A2 => n133, B1 => b(6), B2 => n167, 
                           C1 => b(7), C2 => a(7), ZN => n169);
   U112 : AND2_X1 port map( A1 => n168, A2 => a(6), ZN => n167);
   U113 : AND2_X1 port map( A1 => cout_2_port, A2 => a(12), ZN => n185);
   U114 : OAI21_X1 port map( B1 => n187, B2 => a(15), A => b(15), ZN => n188);
   U115 : OAI21_X1 port map( B1 => n210, B2 => a(23), A => b(23), ZN => n211);
   U116 : OAI211_X1 port map( C1 => b(16), C2 => a(16), A => n233, B => n191, 
                           ZN => n203);

end SYN_p4_carry_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4CarryGenerator_DATA_SIZE32_SPARSITY4_4 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  cout :
         out std_logic_vector (7 downto 0));

end P4CarryGenerator_DATA_SIZE32_SPARSITY4_4;

architecture SYN_p4_carry_generator_arch of 
   P4CarryGenerator_DATA_SIZE32_SPARSITY4_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal cout_7_port, cout_5_port, n250, n251, n252, n253, n123, n124, n125, 
      n126, cout_2_port, n128, n129, n130, n131, n132, n133, cout_4_port, n135,
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, cout_6_port, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, cout_0_port, cout_1_port, 
      cout_3_port, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, 
      n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, 
      n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, 
      n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, 
      n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, 
      n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, 
      n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249 : 
      std_logic;

begin
   cout <= ( cout_7_port, cout_6_port, cout_5_port, cout_4_port, cout_3_port, 
      cout_2_port, cout_1_port, cout_0_port );
   
   U95 : NAND3_X1 port map( A1 => a(16), A2 => n209, A3 => b(16), ZN => n210);
   U1 : INV_X1 port map( A => a(27), ZN => n157);
   U2 : AND2_X1 port map( A1 => n145, A2 => a(12), ZN => n133);
   U3 : INV_X1 port map( A => a(5), ZN => n139);
   U4 : OAI222_X1 port map( A1 => a(28), A2 => n153, B1 => b(28), B2 => n240, 
                           C1 => b(29), C2 => a(29), ZN => n241);
   U5 : AND2_X1 port map( A1 => n150, A2 => n151, ZN => n123);
   U6 : INV_X1 port map( A => b(27), ZN => n158);
   U7 : CLKBUF_X1 port map( A => n250, Z => n129);
   U8 : CLKBUF_X1 port map( A => n176, Z => n124);
   U9 : NAND2_X1 port map( A1 => n169, A2 => n125, ZN => n232);
   U10 : AND2_X1 port map( A1 => n229, A2 => n126, ZN => n125);
   U11 : INV_X1 port map( A => a(24), ZN => n126);
   U12 : CLKBUF_X1 port map( A => n152, Z => cout_2_port);
   U13 : OAI21_X1 port map( B1 => n203, B2 => n202, A => n201, ZN => n152);
   U14 : OAI22_X1 port map( A1 => n157, A2 => n158, B1 => n239, B2 => n159, ZN 
                           => cout_6_port);
   U15 : OAI22_X1 port map( A1 => n154, A2 => a(4), B1 => b(4), B2 => n181, ZN 
                           => n128);
   U16 : NAND2_X1 port map( A1 => n200, A2 => n133, ZN => n130);
   U17 : NAND2_X1 port map( A1 => n130, A2 => n131, ZN => n204);
   U18 : OR2_X1 port map( A1 => n132, A2 => n144, ZN => n131);
   U19 : INV_X1 port map( A => a(12), ZN => n132);
   U20 : CLKBUF_X1 port map( A => n129, Z => cout_4_port);
   U21 : OAI221_X1 port map( B1 => n221, B2 => n220, C1 => n219, C2 => n218, A 
                           => n217, ZN => n250);
   U22 : OR2_X1 port map( A1 => n190, A2 => n189, ZN => n135);
   U23 : NAND2_X1 port map( A1 => n188, A2 => n135, ZN => n252);
   U24 : CLKBUF_X1 port map( A => b(0), Z => n136);
   U25 : AND2_X1 port map( A1 => n161, A2 => n155, ZN => n137);
   U26 : NAND2_X1 port map( A1 => n205, A2 => n123, ZN => n161);
   U27 : OR2_X1 port map( A1 => n190, A2 => n189, ZN => n138);
   U28 : NAND2_X1 port map( A1 => n138, A2 => n147, ZN => n146);
   U29 : NOR2_X1 port map( A1 => n182, A2 => n139, ZN => n183);
   U30 : CLKBUF_X1 port map( A => n179, Z => n140);
   U31 : CLKBUF_X1 port map( A => n227, Z => n141);
   U32 : AND2_X1 port map( A1 => b(9), A2 => a(9), ZN => n142);
   U33 : NOR2_X1 port map( A1 => n195, A2 => n142, ZN => n199);
   U34 : CLKBUF_X1 port map( A => n187, Z => n143);
   U35 : OR2_X1 port map( A1 => n203, A2 => n202, ZN => n144);
   U36 : OR2_X1 port map( A1 => a(11), A2 => b(11), ZN => n145);
   U37 : NAND2_X1 port map( A1 => n200, A2 => n145, ZN => n201);
   U38 : OAI222_X1 port map( A1 => a(6), A2 => n143, B1 => n186, B2 => b(6), C1
                           => b(7), C2 => a(7), ZN => n147);
   U39 : OR2_X1 port map( A1 => n208, A2 => n207, ZN => n148);
   U40 : NAND2_X1 port map( A1 => n206, A2 => n148, ZN => n251);
   U41 : OR2_X1 port map( A1 => n225, A2 => n224, ZN => n149);
   U42 : NAND2_X1 port map( A1 => n149, A2 => n223, ZN => n227);
   U43 : OR2_X1 port map( A1 => n162, A2 => n163, ZN => n150);
   U44 : OR2_X1 port map( A1 => n164, A2 => n165, ZN => n151);
   U45 : INV_X1 port map( A => a(14), ZN => n162);
   U46 : INV_X1 port map( A => b(14), ZN => n163);
   U47 : INV_X1 port map( A => a(13), ZN => n164);
   U48 : INV_X1 port map( A => b(13), ZN => n165);
   U49 : CLKBUF_X1 port map( A => cout_6_port, Z => n153);
   U50 : NAND2_X2 port map( A1 => n169, A2 => n229, ZN => cout_5_port);
   U51 : CLKBUF_X1 port map( A => n253, Z => n154);
   U52 : OR2_X1 port map( A1 => b(14), A2 => a(14), ZN => n155);
   U53 : NAND2_X1 port map( A1 => n161, A2 => n155, ZN => n208);
   U54 : NOR2_X1 port map( A1 => a(27), A2 => b(27), ZN => n159);
   U55 : INV_X1 port map( A => n228, ZN => n160);
   U56 : CLKBUF_X1 port map( A => n154, Z => cout_0_port);
   U57 : CLKBUF_X1 port map( A => n252, Z => cout_1_port);
   U58 : CLKBUF_X1 port map( A => n251, Z => cout_3_port);
   U59 : OR2_X1 port map( A1 => n160, A2 => n230, ZN => n169);
   U60 : INV_X1 port map( A => b(17), ZN => n211);
   U61 : INV_X1 port map( A => b(21), ZN => n224);
   U62 : NAND2_X1 port map( A1 => n211, A2 => n212, ZN => n209);
   U63 : INV_X1 port map( A => n219, ZN => n216);
   U64 : INV_X1 port map( A => b(25), ZN => n233);
   U65 : INV_X1 port map( A => b(29), ZN => n242);
   U66 : OAI21_X1 port map( B1 => n249, B2 => n248, A => n247, ZN => 
                           cout_7_port);
   U67 : INV_X1 port map( A => a(7), ZN => n190);
   U68 : INV_X1 port map( A => b(7), ZN => n189);
   U69 : INV_X1 port map( A => a(11), ZN => n203);
   U70 : INV_X1 port map( A => b(11), ZN => n202);
   U71 : OAI22_X1 port map( A1 => a(2), A2 => n124, B1 => b(2), B2 => n175, ZN 
                           => n177);
   U72 : AND2_X1 port map( A1 => n176, A2 => a(2), ZN => n175);
   U73 : OAI22_X1 port map( A1 => a(1), A2 => n173, B1 => b(1), B2 => n172, ZN 
                           => n174);
   U74 : OR2_X1 port map( A1 => a(26), A2 => b(26), ZN => n238);
   U75 : INV_X1 port map( A => a(25), ZN => n234);
   U76 : OAI22_X1 port map( A1 => n199, A2 => n198, B1 => n197, B2 => n196, ZN 
                           => n200);
   U77 : INV_X1 port map( A => a(10), ZN => n197);
   U78 : NOR2_X1 port map( A1 => b(10), A2 => a(10), ZN => n198);
   U79 : INV_X1 port map( A => b(10), ZN => n196);
   U80 : AOI22_X1 port map( A1 => n193, A2 => n194, B1 => n192, B2 => n191, ZN 
                           => n195);
   U81 : INV_X1 port map( A => a(9), ZN => n192);
   U82 : INV_X1 port map( A => b(9), ZN => n191);
   U83 : OAI22_X1 port map( A1 => a(22), A2 => n141, B1 => b(22), B2 => n226, 
                           ZN => n231);
   U84 : AND2_X1 port map( A1 => n227, A2 => a(22), ZN => n226);
   U85 : INV_X1 port map( A => a(21), ZN => n225);
   U86 : OAI21_X1 port map( B1 => a(18), B2 => n215, A => n214, ZN => n219);
   U87 : INV_X1 port map( A => n213, ZN => n214);
   U88 : AOI21_X1 port map( B1 => n215, B2 => a(18), A => b(18), ZN => n213);
   U89 : OAI21_X1 port map( B1 => n212, B2 => n211, A => n210, ZN => n215);
   U90 : INV_X1 port map( A => a(15), ZN => n207);
   U91 : INV_X1 port map( A => a(23), ZN => n230);
   U92 : AND2_X1 port map( A1 => n179, A2 => a(3), ZN => n178);
   U93 : INV_X1 port map( A => a(19), ZN => n218);
   U94 : OAI22_X1 port map( A1 => b(19), A2 => a(19), B1 => b(18), B2 => a(18),
                           ZN => n220);
   U96 : OAI21_X1 port map( B1 => n216, B2 => a(19), A => b(19), ZN => n217);
   U97 : INV_X1 port map( A => n185, ZN => n187);
   U98 : AND2_X1 port map( A1 => n173, A2 => a(1), ZN => n172);
   U99 : OAI222_X1 port map( A1 => a(20), A2 => n129, B1 => n222, B2 => b(20), 
                           C1 => b(21), C2 => a(21), ZN => n223);
   U100 : NOR2_X1 port map( A1 => b(25), A2 => a(25), ZN => n235);
   U101 : OAI22_X1 port map( A1 => a(30), A2 => n245, B1 => b(30), B2 => n244, 
                           ZN => n249);
   U102 : AND2_X1 port map( A1 => n245, A2 => a(30), ZN => n244);
   U103 : OAI21_X1 port map( B1 => n243, B2 => n242, A => n241, ZN => n245);
   U104 : INV_X1 port map( A => a(29), ZN => n243);
   U105 : OAI21_X1 port map( B1 => n246, B2 => a(31), A => b(31), ZN => n247);
   U106 : INV_X1 port map( A => n249, ZN => n246);
   U107 : INV_X1 port map( A => a(17), ZN => n212);
   U108 : INV_X1 port map( A => a(31), ZN => n248);
   U109 : OAI222_X1 port map( A1 => n152, A2 => a(12), B1 => b(12), B2 => n204,
                           C1 => b(13), C2 => a(13), ZN => n205);
   U110 : INV_X1 port map( A => n231, ZN => n228);
   U111 : OAI22_X1 port map( A1 => a(3), A2 => n140, B1 => b(3), B2 => n178, ZN
                           => n180);
   U112 : OAI21_X1 port map( B1 => n137, B2 => a(15), A => b(15), ZN => n206);
   U113 : OAI21_X1 port map( B1 => n228, B2 => a(23), A => b(23), ZN => n229);
   U114 : OAI222_X1 port map( A1 => a(6), A2 => n143, B1 => b(6), B2 => n186, 
                           C1 => b(7), C2 => a(7), ZN => n188);
   U115 : AND2_X1 port map( A1 => n187, A2 => a(6), ZN => n186);
   U116 : OAI22_X1 port map( A1 => n236, A2 => n235, B1 => n234, B2 => n233, ZN
                           => n237);
   U117 : OAI22_X1 port map( A1 => n154, A2 => a(4), B1 => b(4), B2 => n181, ZN
                           => n182);
   U118 : AND2_X1 port map( A1 => n253, A2 => a(4), ZN => n181);
   U119 : INV_X1 port map( A => n180, ZN => n253);
   U120 : INV_X1 port map( A => n171, ZN => n173);
   U121 : OAI22_X1 port map( A1 => a(5), A2 => n184, B1 => b(5), B2 => n183, ZN
                           => n185);
   U122 : INV_X1 port map( A => n128, ZN => n184);
   U123 : OAI22_X1 port map( A1 => n136, A2 => a(0), B1 => cin, B2 => n170, ZN 
                           => n171);
   U124 : AND2_X1 port map( A1 => b(0), A2 => a(0), ZN => n170);
   U125 : AND2_X1 port map( A1 => n153, A2 => a(28), ZN => n240);
   U126 : AOI22_X1 port map( A1 => b(26), A2 => a(26), B1 => n237, B2 => n238, 
                           ZN => n239);
   U127 : AOI22_X1 port map( A1 => n232, A2 => b(24), B1 => a(24), B2 => 
                           cout_5_port, ZN => n236);
   U128 : AND2_X1 port map( A1 => n250, A2 => a(20), ZN => n222);
   U129 : OAI211_X1 port map( C1 => b(16), C2 => a(16), A => n251, B => n209, 
                           ZN => n221);
   U130 : NAND2_X1 port map( A1 => n252, A2 => a(8), ZN => n194);
   U131 : OAI21_X1 port map( B1 => n146, B2 => a(8), A => b(8), ZN => n193);
   U132 : INV_X1 port map( A => n177, ZN => n179);
   U133 : INV_X1 port map( A => n174, ZN => n176);

end SYN_p4_carry_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4CarryGenerator_DATA_SIZE32_SPARSITY4_3 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  cout :
         out std_logic_vector (7 downto 0));

end P4CarryGenerator_DATA_SIZE32_SPARSITY4_3;

architecture SYN_p4_carry_generator_arch of 
   P4CarryGenerator_DATA_SIZE32_SPARSITY4_3 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X4
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal cout_7_port, n258, n259, n260, n261, n262, n263, n105, n123, n124, 
      n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, cout_4_port, 
      n136, n137, n138, n139, n140, n141, n142, n143, cout_5_port, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, cout_2_port, n165, n166, n167, n168, n169, 
      n170, cout_6_port, n172, n173, cout_0_port, n175, cout_3_port, n177, 
      cout_1_port, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, 
      n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, 
      n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, 
      n213, n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, 
      n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, 
      n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, 
      n249, n250, n251, n252, n253, n254, n255, n256, n257 : std_logic;

begin
   cout <= ( cout_7_port, cout_6_port, cout_5_port, cout_4_port, cout_3_port, 
      cout_2_port, cout_1_port, cout_0_port );
   
   U95 : NAND3_X1 port map( A1 => a(16), A2 => n217, A3 => b(16), ZN => n218);
   U1 : INV_X1 port map( A => a(27), ZN => n172);
   U2 : INV_X1 port map( A => a(6), ZN => n139);
   U3 : INV_X1 port map( A => a(6), ZN => n138);
   U4 : OAI222_X1 port map( A1 => a(28), A2 => n160, B1 => b(28), B2 => n248, 
                           C1 => b(29), C2 => a(29), ZN => n249);
   U5 : AND2_X1 port map( A1 => n161, A2 => n162, ZN => n105);
   U6 : NOR2_X1 port map( A1 => a(27), A2 => b(27), ZN => n123);
   U7 : INV_X1 port map( A => b(27), ZN => n173);
   U8 : OAI22_X1 port map( A1 => a(22), A2 => n131, B1 => n234, B2 => b(22), ZN
                           => n124);
   U9 : AND2_X1 port map( A1 => n193, A2 => a(5), ZN => n192);
   U10 : NAND2_X1 port map( A1 => n194, A2 => n128, ZN => n125);
   U11 : NAND2_X1 port map( A1 => n125, A2 => n126, ZN => n141);
   U12 : OR2_X1 port map( A1 => n127, A2 => n134, ZN => n126);
   U13 : INV_X1 port map( A => n163, ZN => n127);
   U14 : AND2_X1 port map( A1 => n139, A2 => n163, ZN => n128);
   U15 : AND2_X1 port map( A1 => n166, A2 => n165, ZN => n129);
   U16 : CLKBUF_X1 port map( A => n182, Z => n130);
   U17 : CLKBUF_X1 port map( A => n235, Z => n131);
   U18 : NAND2_X1 port map( A1 => n208, A2 => n157, ZN => n132);
   U19 : NAND2_X1 port map( A1 => n133, A2 => n134, ZN => n147);
   U20 : NAND2_X1 port map( A1 => n139, A2 => n194, ZN => n133);
   U21 : OR2_X1 port map( A1 => b(7), A2 => a(7), ZN => n134);
   U22 : OAI221_X4 port map( B1 => n136, B2 => n228, C1 => n227, C2 => n226, A 
                           => n225, ZN => cout_4_port);
   U23 : OAI211_X1 port map( C1 => b(16), C2 => a(16), A => n260, B => n217, ZN
                           => n136);
   U24 : OAI221_X1 port map( B1 => n229, B2 => n228, C1 => n227, C2 => n226, A 
                           => n225, ZN => n259);
   U25 : OAI22_X1 port map( A1 => a(5), A2 => n151, B1 => n192, B2 => b(5), ZN 
                           => n137);
   U26 : NOR2_X1 port map( A1 => n137, A2 => n138, ZN => n195);
   U27 : NOR2_X1 port map( A1 => n142, A2 => n195, ZN => n140);
   U28 : NOR2_X1 port map( A1 => n140, A2 => n141, ZN => n262);
   U29 : OR2_X1 port map( A1 => b(6), A2 => n127, ZN => n142);
   U30 : OR2_X1 port map( A1 => n211, A2 => n210, ZN => n143);
   U31 : NAND2_X1 port map( A1 => n209, A2 => n143, ZN => n261);
   U32 : INV_X1 port map( A => b(11), ZN => n210);
   U33 : CLKBUF_X1 port map( A => n258, Z => cout_5_port);
   U34 : OAI21_X1 port map( B1 => n236, B2 => a(23), A => b(23), ZN => n145);
   U35 : CLKBUF_X1 port map( A => n185, Z => n146);
   U36 : OR2_X1 port map( A1 => n175, A2 => n147, ZN => n196);
   U37 : OR2_X1 port map( A1 => n233, A2 => n232, ZN => n148);
   U38 : NAND2_X1 port map( A1 => n148, A2 => n231, ZN => n235);
   U39 : CLKBUF_X1 port map( A => n188, Z => n149);
   U40 : CLKBUF_X1 port map( A => b(0), Z => n150);
   U41 : CLKBUF_X1 port map( A => n193, Z => n151);
   U42 : AND2_X1 port map( A1 => b(9), A2 => a(9), ZN => n152);
   U43 : NOR2_X1 port map( A1 => n203, A2 => n152, ZN => n207);
   U44 : NAND2_X1 port map( A1 => n196, A2 => n163, ZN => n153);
   U45 : OR2_X1 port map( A1 => n216, A2 => n215, ZN => n154);
   U46 : NAND2_X1 port map( A1 => n214, A2 => n154, ZN => n260);
   U47 : OR2_X1 port map( A1 => n211, A2 => n210, ZN => n155);
   U48 : NAND2_X1 port map( A1 => n132, A2 => n155, ZN => cout_2_port);
   U49 : CLKBUF_X1 port map( A => n263, Z => n156);
   U50 : NAND2_X1 port map( A1 => n105, A2 => n213, ZN => n166);
   U51 : OR2_X1 port map( A1 => a(11), A2 => b(11), ZN => n157);
   U52 : NAND2_X1 port map( A1 => n208, A2 => n157, ZN => n209);
   U53 : NAND2_X1 port map( A1 => n177, A2 => n158, ZN => n240);
   U54 : AND2_X1 port map( A1 => n145, A2 => n159, ZN => n158);
   U55 : INV_X1 port map( A => a(24), ZN => n159);
   U56 : CLKBUF_X1 port map( A => cout_6_port, Z => n160);
   U57 : OAI22_X1 port map( A1 => n172, A2 => n173, B1 => n247, B2 => n123, ZN 
                           => cout_6_port);
   U58 : NAND2_X1 port map( A1 => n177, A2 => n237, ZN => n258);
   U59 : OR2_X1 port map( A1 => n167, A2 => n168, ZN => n161);
   U60 : OR2_X1 port map( A1 => n169, A2 => n170, ZN => n162);
   U61 : INV_X1 port map( A => a(14), ZN => n167);
   U62 : INV_X1 port map( A => b(14), ZN => n168);
   U63 : INV_X1 port map( A => a(13), ZN => n169);
   U64 : INV_X1 port map( A => b(13), ZN => n170);
   U65 : OAI222_X1 port map( A1 => a(12), A2 => cout_2_port, B1 => b(12), B2 =>
                           n212, C1 => b(13), C2 => a(13), ZN => n213);
   U66 : OR2_X1 port map( A1 => n198, A2 => n197, ZN => n163);
   U67 : OR2_X1 port map( A1 => b(14), A2 => a(14), ZN => n165);
   U68 : NAND2_X1 port map( A1 => n166, A2 => n165, ZN => n216);
   U69 : CLKBUF_X1 port map( A => n156, Z => cout_0_port);
   U70 : NOR2_X1 port map( A1 => n195, A2 => b(6), ZN => n175);
   U71 : CLKBUF_X1 port map( A => n260, Z => cout_3_port);
   U72 : OR2_X1 port map( A1 => n239, A2 => n238, ZN => n177);
   U73 : CLKBUF_X1 port map( A => n153, Z => cout_1_port);
   U74 : INV_X1 port map( A => b(17), ZN => n219);
   U75 : INV_X1 port map( A => b(21), ZN => n232);
   U76 : INV_X1 port map( A => b(25), ZN => n241);
   U77 : INV_X1 port map( A => b(29), ZN => n250);
   U78 : NAND2_X1 port map( A1 => n219, A2 => n220, ZN => n217);
   U79 : INV_X1 port map( A => n227, ZN => n224);
   U80 : OAI21_X1 port map( B1 => n257, B2 => n256, A => n255, ZN => 
                           cout_7_port);
   U81 : INV_X1 port map( A => a(7), ZN => n198);
   U82 : INV_X1 port map( A => b(7), ZN => n197);
   U83 : AND2_X1 port map( A1 => n235, A2 => a(22), ZN => n234);
   U84 : INV_X1 port map( A => a(21), ZN => n233);
   U85 : INV_X1 port map( A => a(10), ZN => n205);
   U86 : NOR2_X1 port map( A1 => b(10), A2 => a(10), ZN => n206);
   U87 : INV_X1 port map( A => b(10), ZN => n204);
   U88 : INV_X1 port map( A => a(11), ZN => n211);
   U89 : OR2_X1 port map( A1 => a(26), A2 => b(26), ZN => n246);
   U90 : INV_X1 port map( A => a(25), ZN => n242);
   U91 : INV_X1 port map( A => a(15), ZN => n215);
   U92 : AOI22_X1 port map( A1 => n201, A2 => n202, B1 => n200, B2 => n199, ZN 
                           => n203);
   U93 : INV_X1 port map( A => a(9), ZN => n200);
   U94 : INV_X1 port map( A => b(9), ZN => n199);
   U96 : OAI21_X1 port map( B1 => a(18), B2 => n223, A => n222, ZN => n227);
   U97 : INV_X1 port map( A => n221, ZN => n222);
   U98 : AOI21_X1 port map( B1 => n223, B2 => a(18), A => b(18), ZN => n221);
   U99 : OAI21_X1 port map( B1 => n220, B2 => n219, A => n218, ZN => n223);
   U100 : INV_X1 port map( A => a(19), ZN => n226);
   U101 : OAI22_X1 port map( A1 => b(19), A2 => a(19), B1 => b(18), B2 => a(18)
                           , ZN => n228);
   U102 : OAI21_X1 port map( B1 => n224, B2 => a(19), A => b(19), ZN => n225);
   U103 : OAI22_X1 port map( A1 => a(2), A2 => n146, B1 => b(2), B2 => n184, ZN
                           => n186);
   U104 : AND2_X1 port map( A1 => n185, A2 => a(2), ZN => n184);
   U105 : OAI22_X1 port map( A1 => a(1), A2 => n130, B1 => b(1), B2 => n181, ZN
                           => n183);
   U106 : INV_X1 port map( A => a(23), ZN => n238);
   U107 : INV_X1 port map( A => n124, ZN => n236);
   U108 : AND2_X1 port map( A1 => n182, A2 => a(1), ZN => n181);
   U109 : NOR2_X1 port map( A1 => b(25), A2 => a(25), ZN => n243);
   U110 : AND2_X1 port map( A1 => n160, A2 => a(28), ZN => n248);
   U111 : OAI22_X1 port map( A1 => a(30), A2 => n253, B1 => b(30), B2 => n252, 
                           ZN => n257);
   U112 : AND2_X1 port map( A1 => n253, A2 => a(30), ZN => n252);
   U113 : OAI21_X1 port map( B1 => n251, B2 => n250, A => n249, ZN => n253);
   U114 : INV_X1 port map( A => a(29), ZN => n251);
   U115 : OAI21_X1 port map( B1 => n254, B2 => a(31), A => b(31), ZN => n255);
   U116 : INV_X1 port map( A => n257, ZN => n254);
   U117 : INV_X1 port map( A => a(17), ZN => n220);
   U118 : INV_X1 port map( A => a(31), ZN => n256);
   U119 : NAND2_X1 port map( A1 => n153, A2 => a(8), ZN => n202);
   U120 : AOI22_X1 port map( A1 => b(24), A2 => n240, B1 => n258, B2 => a(24), 
                           ZN => n244);
   U121 : OAI22_X1 port map( A1 => a(22), A2 => n131, B1 => n234, B2 => b(22), 
                           ZN => n239);
   U122 : OAI22_X1 port map( A1 => n207, A2 => n206, B1 => n205, B2 => n204, ZN
                           => n208);
   U123 : INV_X1 port map( A => n180, ZN => n182);
   U124 : INV_X1 port map( A => n189, ZN => n263);
   U125 : INV_X1 port map( A => n191, ZN => n193);
   U126 : OAI22_X1 port map( A1 => n150, A2 => a(0), B1 => n179, B2 => cin, ZN 
                           => n180);
   U127 : AND2_X1 port map( A1 => b(0), A2 => a(0), ZN => n179);
   U128 : OAI22_X1 port map( A1 => a(3), A2 => n149, B1 => b(3), B2 => n187, ZN
                           => n189);
   U129 : AND2_X1 port map( A1 => n188, A2 => a(3), ZN => n187);
   U130 : OAI22_X1 port map( A1 => a(4), A2 => n156, B1 => b(4), B2 => n190, ZN
                           => n191);
   U131 : AND2_X1 port map( A1 => n263, A2 => a(4), ZN => n190);
   U132 : OAI22_X1 port map( A1 => n244, A2 => n243, B1 => n242, B2 => n241, ZN
                           => n245);
   U133 : OAI222_X1 port map( A1 => a(20), A2 => cout_4_port, B1 => b(20), B2 
                           => n230, C1 => b(21), C2 => a(21), ZN => n231);
   U134 : AND2_X1 port map( A1 => n259, A2 => a(20), ZN => n230);
   U135 : AOI22_X1 port map( A1 => b(26), A2 => a(26), B1 => n245, B2 => n246, 
                           ZN => n247);
   U136 : INV_X1 port map( A => n186, ZN => n188);
   U137 : INV_X1 port map( A => n183, ZN => n185);
   U138 : AND2_X1 port map( A1 => n261, A2 => a(12), ZN => n212);
   U139 : OAI21_X1 port map( B1 => n262, B2 => a(8), A => b(8), ZN => n201);
   U140 : OAI211_X1 port map( C1 => b(16), C2 => a(16), A => n260, B => n217, 
                           ZN => n229);
   U141 : OAI22_X1 port map( A1 => a(5), A2 => n151, B1 => n192, B2 => b(5), ZN
                           => n194);
   U142 : OAI21_X1 port map( B1 => n129, B2 => a(15), A => b(15), ZN => n214);
   U143 : OAI21_X1 port map( B1 => a(23), B2 => n236, A => b(23), ZN => n237);

end SYN_p4_carry_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4CarryGenerator_DATA_SIZE32_SPARSITY4_2 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  cout :
         out std_logic_vector (7 downto 0));

end P4CarryGenerator_DATA_SIZE32_SPARSITY4_2;

architecture SYN_p4_carry_generator_arch of 
   P4CarryGenerator_DATA_SIZE32_SPARSITY4_2 is

   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal cout_7_port, n248, n249, n250, n251, n252, n123, n124, n125, 
      cout_3_port, n127, n128, n129, n130, n131, cout_5_port, cout_1_port, n134
      , n135, n136, n137, cout_0_port, n139, n140, n141, n142, n143, n144, n145
      , n146, n147, n148, cout_4_port, n150, cout_6_port, n152, n153, n154, 
      n155, cout_2_port, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, 
      n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, 
      n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, 
      n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, 
      n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, 
      n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, 
      n238, n239, n240, n241, n242, n243, n244, n245, n246, n247 : std_logic;

begin
   cout <= ( cout_7_port, cout_6_port, cout_5_port, cout_4_port, cout_3_port, 
      cout_2_port, cout_1_port, cout_0_port );
   
   U95 : NAND3_X1 port map( A1 => a(16), A2 => n207, A3 => b(16), ZN => n208);
   U1 : INV_X1 port map( A => a(27), ZN => n152);
   U2 : NOR2_X1 port map( A1 => b(13), A2 => a(13), ZN => n159);
   U3 : OAI222_X1 port map( A1 => a(28), A2 => n146, B1 => b(28), B2 => n238, 
                           C1 => b(29), C2 => a(29), ZN => n239);
   U4 : CLKBUF_X1 port map( A => n183, Z => n123);
   U5 : CLKBUF_X1 port map( A => n129, Z => n124);
   U6 : CLKBUF_X1 port map( A => n186, Z => n125);
   U7 : CLKBUF_X1 port map( A => n250, Z => cout_3_port);
   U8 : CLKBUF_X1 port map( A => n252, Z => n127);
   U9 : OAI21_X1 port map( B1 => n226, B2 => a(23), A => b(23), ZN => n128);
   U10 : NAND2_X1 port map( A1 => n199, A2 => n147, ZN => n129);
   U11 : AND2_X1 port map( A1 => n129, A2 => n130, ZN => n157);
   U12 : AND2_X1 port map( A1 => n131, A2 => n144, ZN => n130);
   U13 : INV_X1 port map( A => a(12), ZN => n131);
   U14 : BUF_X1 port map( A => n248, Z => cout_5_port);
   U15 : CLKBUF_X1 port map( A => n148, Z => cout_1_port);
   U16 : BUF_X2 port map( A => n249, Z => cout_4_port);
   U17 : NAND2_X1 port map( A1 => n154, A2 => n155, ZN => n134);
   U18 : NAND2_X1 port map( A1 => n202, A2 => n135, ZN => n163);
   U19 : INV_X1 port map( A => n134, ZN => n135);
   U20 : OR2_X1 port map( A1 => n164, A2 => n165, ZN => n154);
   U21 : OR2_X1 port map( A1 => n166, A2 => n167, ZN => n155);
   U22 : NOR2_X1 port map( A1 => a(27), A2 => b(27), ZN => n136);
   U23 : INV_X1 port map( A => b(12), ZN => n141);
   U24 : INV_X1 port map( A => b(27), ZN => n153);
   U25 : AND2_X1 port map( A1 => b(9), A2 => a(9), ZN => n137);
   U26 : NOR2_X1 port map( A1 => n194, A2 => n137, ZN => n198);
   U27 : CLKBUF_X1 port map( A => n127, Z => cout_0_port);
   U28 : OR2_X1 port map( A1 => n189, A2 => n188, ZN => n139);
   U29 : NAND2_X1 port map( A1 => n139, A2 => n187, ZN => n148);
   U30 : CLKBUF_X1 port map( A => b(0), Z => n140);
   U31 : AND2_X1 port map( A1 => n141, A2 => n142, ZN => n158);
   U32 : NAND2_X1 port map( A1 => n251, A2 => a(12), ZN => n142);
   U33 : OR2_X1 port map( A1 => n223, A2 => n222, ZN => n143);
   U34 : NAND2_X1 port map( A1 => n221, A2 => n143, ZN => n225);
   U35 : OR2_X1 port map( A1 => n201, A2 => n200, ZN => n144);
   U36 : NAND2_X1 port map( A1 => n144, A2 => n124, ZN => cout_2_port);
   U37 : OR2_X1 port map( A1 => n201, A2 => n200, ZN => n145);
   U38 : NAND2_X1 port map( A1 => n129, A2 => n145, ZN => n251);
   U39 : CLKBUF_X1 port map( A => cout_6_port, Z => n146);
   U40 : OR2_X1 port map( A1 => a(11), A2 => b(11), ZN => n147);
   U41 : OAI22_X1 port map( A1 => n152, A2 => n153, B1 => n237, B2 => n136, ZN 
                           => cout_6_port);
   U42 : OR2_X1 port map( A1 => n206, A2 => n205, ZN => n150);
   U43 : NAND2_X1 port map( A1 => n204, A2 => n150, ZN => n250);
   U44 : OAI221_X1 port map( B1 => n219, B2 => n218, C1 => n217, C2 => n216, A 
                           => n215, ZN => n249);
   U45 : INV_X1 port map( A => a(14), ZN => n164);
   U46 : INV_X1 port map( A => b(14), ZN => n165);
   U47 : INV_X1 port map( A => a(13), ZN => n166);
   U48 : INV_X1 port map( A => b(13), ZN => n167);
   U49 : OR3_X1 port map( A1 => n157, A2 => n158, A3 => n159, ZN => n202);
   U50 : NAND2_X1 port map( A1 => n168, A2 => n160, ZN => n230);
   U51 : AND2_X1 port map( A1 => n128, A2 => n161, ZN => n160);
   U52 : INV_X1 port map( A => a(24), ZN => n161);
   U53 : OR2_X1 port map( A1 => b(14), A2 => a(14), ZN => n162);
   U54 : NAND2_X1 port map( A1 => n162, A2 => n163, ZN => n206);
   U55 : OR2_X1 port map( A1 => n228, A2 => n229, ZN => n168);
   U56 : NAND2_X1 port map( A1 => n227, A2 => n168, ZN => n248);
   U57 : INV_X1 port map( A => b(17), ZN => n209);
   U58 : NAND2_X1 port map( A1 => n209, A2 => n210, ZN => n207);
   U59 : INV_X1 port map( A => n217, ZN => n214);
   U60 : INV_X1 port map( A => b(25), ZN => n231);
   U61 : INV_X1 port map( A => b(21), ZN => n222);
   U62 : INV_X1 port map( A => b(29), ZN => n240);
   U63 : OAI21_X1 port map( B1 => n247, B2 => n246, A => n245, ZN => 
                           cout_7_port);
   U64 : INV_X1 port map( A => a(15), ZN => n205);
   U65 : INV_X1 port map( A => n206, ZN => n203);
   U66 : INV_X1 port map( A => a(7), ZN => n189);
   U67 : INV_X1 port map( A => b(7), ZN => n188);
   U68 : OAI22_X1 port map( A1 => a(22), A2 => n225, B1 => b(22), B2 => n224, 
                           ZN => n229);
   U69 : AND2_X1 port map( A1 => n225, A2 => a(22), ZN => n224);
   U70 : INV_X1 port map( A => a(21), ZN => n223);
   U71 : OR2_X1 port map( A1 => a(26), A2 => b(26), ZN => n236);
   U72 : INV_X1 port map( A => a(25), ZN => n232);
   U73 : INV_X1 port map( A => n184, ZN => n186);
   U74 : OAI22_X1 port map( A1 => a(5), A2 => n123, B1 => b(5), B2 => n182, ZN 
                           => n184);
   U75 : AND2_X1 port map( A1 => n183, A2 => a(5), ZN => n182);
   U76 : INV_X1 port map( A => n181, ZN => n183);
   U77 : OAI22_X1 port map( A1 => a(4), A2 => n127, B1 => b(4), B2 => n180, ZN 
                           => n181);
   U78 : AND2_X1 port map( A1 => n252, A2 => a(4), ZN => n180);
   U79 : INV_X1 port map( A => n179, ZN => n252);
   U80 : OAI22_X1 port map( A1 => a(3), A2 => n178, B1 => b(3), B2 => n177, ZN 
                           => n179);
   U81 : AND2_X1 port map( A1 => n178, A2 => a(3), ZN => n177);
   U82 : INV_X1 port map( A => a(11), ZN => n201);
   U83 : INV_X1 port map( A => b(11), ZN => n200);
   U84 : INV_X1 port map( A => a(23), ZN => n228);
   U85 : INV_X1 port map( A => n229, ZN => n226);
   U86 : OAI22_X1 port map( A1 => n198, A2 => n197, B1 => n196, B2 => n195, ZN 
                           => n199);
   U87 : INV_X1 port map( A => a(10), ZN => n196);
   U88 : NOR2_X1 port map( A1 => b(10), A2 => a(10), ZN => n197);
   U89 : INV_X1 port map( A => b(10), ZN => n195);
   U90 : AOI22_X1 port map( A1 => n192, A2 => n193, B1 => n191, B2 => n190, ZN 
                           => n194);
   U91 : INV_X1 port map( A => a(9), ZN => n191);
   U92 : INV_X1 port map( A => b(9), ZN => n190);
   U93 : OAI21_X1 port map( B1 => a(18), B2 => n213, A => n212, ZN => n217);
   U94 : INV_X1 port map( A => n211, ZN => n212);
   U96 : AOI21_X1 port map( B1 => n213, B2 => a(18), A => b(18), ZN => n211);
   U97 : OAI21_X1 port map( B1 => n210, B2 => n209, A => n208, ZN => n213);
   U98 : INV_X1 port map( A => a(19), ZN => n216);
   U99 : OAI22_X1 port map( A1 => b(19), A2 => a(19), B1 => b(18), B2 => a(18),
                           ZN => n218);
   U100 : OAI21_X1 port map( B1 => n214, B2 => a(19), A => b(19), ZN => n215);
   U101 : NAND2_X1 port map( A1 => n148, A2 => a(8), ZN => n193);
   U102 : OAI222_X1 port map( A1 => cout_4_port, A2 => a(20), B1 => b(20), B2 
                           => n220, C1 => b(21), C2 => a(21), ZN => n221);
   U103 : AND2_X1 port map( A1 => n249, A2 => a(20), ZN => n220);
   U104 : NOR2_X1 port map( A1 => b(25), A2 => a(25), ZN => n233);
   U105 : AND2_X1 port map( A1 => n146, A2 => a(28), ZN => n238);
   U106 : OAI22_X1 port map( A1 => a(30), A2 => n243, B1 => b(30), B2 => n242, 
                           ZN => n247);
   U107 : AND2_X1 port map( A1 => n243, A2 => a(30), ZN => n242);
   U108 : OAI21_X1 port map( B1 => n241, B2 => n240, A => n239, ZN => n243);
   U109 : INV_X1 port map( A => a(29), ZN => n241);
   U110 : OAI21_X1 port map( B1 => n244, B2 => a(31), A => b(31), ZN => n245);
   U111 : INV_X1 port map( A => n247, ZN => n244);
   U112 : INV_X1 port map( A => a(17), ZN => n210);
   U113 : INV_X1 port map( A => a(31), ZN => n246);
   U114 : INV_X1 port map( A => n170, ZN => n172);
   U115 : INV_X1 port map( A => n173, ZN => n175);
   U116 : INV_X1 port map( A => n176, ZN => n178);
   U117 : AOI22_X1 port map( A1 => b(26), A2 => a(26), B1 => n235, B2 => n236, 
                           ZN => n237);
   U118 : OAI21_X1 port map( B1 => n148, B2 => a(8), A => b(8), ZN => n192);
   U119 : OAI22_X1 port map( A1 => n140, A2 => a(0), B1 => cin, B2 => n169, ZN 
                           => n170);
   U120 : AND2_X1 port map( A1 => a(0), A2 => b(0), ZN => n169);
   U121 : OAI22_X1 port map( A1 => n234, A2 => n233, B1 => n232, B2 => n231, ZN
                           => n235);
   U122 : AOI22_X1 port map( A1 => b(24), A2 => n230, B1 => n248, B2 => a(24), 
                           ZN => n234);
   U123 : OAI22_X1 port map( A1 => a(1), A2 => n172, B1 => b(1), B2 => n171, ZN
                           => n173);
   U124 : AND2_X1 port map( A1 => n172, A2 => a(1), ZN => n171);
   U125 : OAI22_X1 port map( A1 => a(2), A2 => n175, B1 => b(2), B2 => n174, ZN
                           => n176);
   U126 : AND2_X1 port map( A1 => n175, A2 => a(2), ZN => n174);
   U127 : OAI222_X1 port map( A1 => a(6), A2 => n125, B1 => b(6), B2 => n185, 
                           C1 => b(7), C2 => a(7), ZN => n187);
   U128 : AND2_X1 port map( A1 => n186, A2 => a(6), ZN => n185);
   U129 : OAI21_X1 port map( B1 => n203, B2 => a(15), A => b(15), ZN => n204);
   U130 : OAI21_X1 port map( B1 => n226, B2 => a(23), A => b(23), ZN => n227);
   U131 : OAI211_X1 port map( C1 => b(16), C2 => a(16), A => n250, B => n207, 
                           ZN => n219);

end SYN_p4_carry_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4CarryGenerator_DATA_SIZE32_SPARSITY4_1 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  cout :
         out std_logic_vector (7 downto 0));

end P4CarryGenerator_DATA_SIZE32_SPARSITY4_1;

architecture SYN_p4_carry_generator_arch of 
   P4CarryGenerator_DATA_SIZE32_SPARSITY4_1 is

   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X4
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal cout_7_port, n240, cout_4_port, n241, n242, n243, n244, n105, n107, 
      n108, n109, n117, n123, n124, cout_5_port, n126, n127, n128, n129, n130, 
      n131, n132, n133, n134, n135, cout_0_port, cout_6_port, n138, n139, n140,
      n141, n142, n143, cout_2_port, n145, cout_3_port, n147, n148, n149, n150,
      n151, n152, n153, n154, n155, cout_1_port, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, 
      n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, 
      n234, n235, n236, n237, n238, n239 : std_logic;

begin
   cout <= ( cout_7_port, cout_6_port, cout_5_port, cout_4_port, cout_3_port, 
      cout_2_port, cout_1_port, cout_0_port );
   
   U95 : NAND3_X1 port map( A1 => a(16), A2 => n199, A3 => b(16), ZN => n200);
   U1 : INV_X1 port map( A => a(24), ZN => n124);
   U2 : CLKBUF_X1 port map( A => n229, Z => n105);
   U3 : OR2_X1 port map( A1 => n193, A2 => n192, ZN => n107);
   U4 : NAND2_X1 port map( A1 => n107, A2 => n191, ZN => cout_2_port);
   U5 : NOR2_X1 port map( A1 => a(27), A2 => b(27), ZN => n108);
   U6 : AND2_X1 port map( A1 => n142, A2 => n141, ZN => n109);
   U7 : INV_X1 port map( A => b(27), ZN => n139);
   U8 : INV_X1 port map( A => a(27), ZN => n138);
   U9 : OAI22_X1 port map( A1 => n138, A2 => n139, B1 => n105, B2 => n108, ZN 
                           => n117);
   U10 : NAND2_X1 port map( A1 => n123, A2 => n219, ZN => n222);
   U11 : AND2_X1 port map( A1 => n161, A2 => n124, ZN => n123);
   U12 : CLKBUF_X1 port map( A => n176, Z => n132);
   U13 : CLKBUF_X1 port map( A => n240, Z => cout_5_port);
   U14 : NAND2_X1 port map( A1 => n219, A2 => n161, ZN => n240);
   U15 : AOI22_X1 port map( A1 => n162, A2 => n132, B1 => n163, B2 => n164, ZN 
                           => n126);
   U16 : AOI22_X1 port map( A1 => n162, A2 => n132, B1 => n163, B2 => n164, ZN 
                           => n127);
   U17 : AND2_X1 port map( A1 => n148, A2 => n145, ZN => n128);
   U18 : CLKBUF_X1 port map( A => n244, Z => n129);
   U19 : OR2_X1 port map( A1 => n193, A2 => n192, ZN => n130);
   U20 : NAND2_X1 port map( A1 => n191, A2 => n130, ZN => n242);
   U21 : OR2_X1 port map( A1 => n221, A2 => n220, ZN => n161);
   U22 : AND2_X1 port map( A1 => b(9), A2 => a(9), ZN => n131);
   U23 : NOR2_X1 port map( A1 => n185, A2 => n131, ZN => n189);
   U24 : NAND2_X1 port map( A1 => n195, A2 => n109, ZN => n148);
   U25 : NOR2_X1 port map( A1 => n169, A2 => n153, ZN => n133);
   U26 : OR2_X1 port map( A1 => n176, A2 => n162, ZN => n164);
   U27 : OAI22_X1 port map( A1 => n138, A2 => n139, B1 => n229, B2 => n108, ZN 
                           => cout_6_port);
   U28 : OR2_X1 port map( A1 => n215, A2 => n214, ZN => n134);
   U29 : NAND2_X1 port map( A1 => n213, A2 => n134, ZN => n217);
   U30 : OAI22_X1 port map( A1 => a(4), A2 => n129, B1 => b(4), B2 => n175, ZN 
                           => n176);
   U31 : OR2_X1 port map( A1 => a(11), A2 => b(11), ZN => n135);
   U32 : NAND2_X1 port map( A1 => n135, A2 => n190, ZN => n191);
   U33 : CLKBUF_X1 port map( A => n129, Z => cout_0_port);
   U34 : OR2_X1 port map( A1 => n180, A2 => n179, ZN => n140);
   U35 : NAND2_X1 port map( A1 => n140, A2 => n178, ZN => n243);
   U36 : OR2_X1 port map( A1 => n149, A2 => n150, ZN => n141);
   U37 : OR2_X1 port map( A1 => n151, A2 => n152, ZN => n142);
   U38 : INV_X1 port map( A => a(14), ZN => n149);
   U39 : INV_X1 port map( A => b(14), ZN => n150);
   U40 : INV_X1 port map( A => a(13), ZN => n151);
   U41 : INV_X1 port map( A => b(13), ZN => n152);
   U42 : OAI22_X1 port map( A1 => a(1), A2 => n168, B1 => b(1), B2 => n167, ZN 
                           => n143);
   U43 : OR2_X1 port map( A1 => b(14), A2 => a(14), ZN => n145);
   U44 : NAND2_X1 port map( A1 => n148, A2 => n145, ZN => n198);
   U45 : CLKBUF_X1 port map( A => n241, Z => cout_3_port);
   U46 : OAI22_X1 port map( A1 => a(2), A2 => n170, B1 => b(2), B2 => n133, ZN 
                           => n147);
   U47 : OAI22_X1 port map( A1 => a(3), A2 => n173, B1 => n172, B2 => b(3), ZN 
                           => n174);
   U48 : INV_X1 port map( A => n174, ZN => n244);
   U49 : OAI22_X1 port map( A1 => a(1), A2 => n168, B1 => b(1), B2 => n167, ZN 
                           => n169);
   U50 : INV_X1 port map( A => a(2), ZN => n153);
   U51 : INV_X1 port map( A => a(3), ZN => n154);
   U52 : INV_X1 port map( A => b(17), ZN => n201);
   U53 : INV_X1 port map( A => b(21), ZN => n214);
   U54 : INV_X1 port map( A => n209, ZN => n206);
   U55 : NAND2_X1 port map( A1 => n201, A2 => n202, ZN => n199);
   U56 : INV_X1 port map( A => n221, ZN => n218);
   U57 : INV_X1 port map( A => b(25), ZN => n223);
   U58 : INV_X1 port map( A => b(29), ZN => n232);
   U59 : OAI21_X1 port map( B1 => n239, B2 => n238, A => n237, ZN => 
                           cout_7_port);
   U60 : AND2_X1 port map( A1 => n217, A2 => a(22), ZN => n216);
   U61 : INV_X1 port map( A => a(21), ZN => n215);
   U62 : INV_X1 port map( A => a(7), ZN => n180);
   U63 : INV_X1 port map( A => b(7), ZN => n179);
   U64 : INV_X1 port map( A => n143, ZN => n170);
   U65 : OAI21_X1 port map( B1 => a(18), B2 => n205, A => n204, ZN => n209);
   U66 : INV_X1 port map( A => n203, ZN => n204);
   U67 : AOI21_X1 port map( B1 => n205, B2 => a(18), A => b(18), ZN => n203);
   U68 : OAI21_X1 port map( B1 => n202, B2 => n201, A => n200, ZN => n205);
   U69 : INV_X1 port map( A => a(11), ZN => n193);
   U70 : INV_X1 port map( A => b(11), ZN => n192);
   U71 : NOR2_X1 port map( A1 => n171, A2 => n154, ZN => n172);
   U72 : OR2_X1 port map( A1 => a(26), A2 => b(26), ZN => n228);
   U73 : INV_X1 port map( A => a(25), ZN => n224);
   U74 : INV_X1 port map( A => a(5), ZN => n162);
   U75 : INV_X1 port map( A => b(5), ZN => n163);
   U76 : OAI22_X1 port map( A1 => n189, A2 => n188, B1 => n187, B2 => n186, ZN 
                           => n190);
   U77 : INV_X1 port map( A => a(10), ZN => n187);
   U78 : INV_X1 port map( A => b(10), ZN => n186);
   U79 : NOR2_X1 port map( A1 => b(10), A2 => a(10), ZN => n188);
   U80 : AOI22_X1 port map( A1 => n183, A2 => n184, B1 => n182, B2 => n181, ZN 
                           => n185);
   U81 : INV_X1 port map( A => a(9), ZN => n182);
   U82 : INV_X1 port map( A => b(9), ZN => n181);
   U83 : INV_X1 port map( A => a(17), ZN => n202);
   U84 : INV_X1 port map( A => a(19), ZN => n208);
   U85 : OAI22_X1 port map( A1 => b(19), A2 => a(19), B1 => b(18), B2 => a(18),
                           ZN => n210);
   U86 : OAI21_X1 port map( B1 => n206, B2 => a(19), A => b(19), ZN => n207);
   U87 : AND2_X1 port map( A1 => n168, A2 => a(1), ZN => n167);
   U88 : OAI222_X1 port map( A1 => a(12), A2 => cout_2_port, B1 => b(12), B2 =>
                           n194, C1 => b(13), C2 => a(13), ZN => n195);
   U89 : NOR2_X1 port map( A1 => b(25), A2 => a(25), ZN => n225);
   U90 : OAI22_X1 port map( A1 => a(30), A2 => n235, B1 => b(30), B2 => n234, 
                           ZN => n239);
   U91 : AND2_X1 port map( A1 => n235, A2 => a(30), ZN => n234);
   U92 : OAI21_X1 port map( B1 => n233, B2 => n232, A => n231, ZN => n235);
   U93 : OAI222_X1 port map( A1 => a(28), A2 => n155, B1 => b(28), B2 => n230, 
                           C1 => b(29), C2 => a(29), ZN => n231);
   U94 : OAI21_X1 port map( B1 => n236, B2 => a(31), A => b(31), ZN => n237);
   U96 : INV_X1 port map( A => n239, ZN => n236);
   U97 : INV_X1 port map( A => a(31), ZN => n238);
   U98 : INV_X1 port map( A => a(29), ZN => n233);
   U99 : INV_X1 port map( A => n166, ZN => n168);
   U100 : CLKBUF_X1 port map( A => n117, Z => n155);
   U101 : CLKBUF_X1 port map( A => n243, Z => cout_1_port);
   U102 : OR2_X1 port map( A1 => a(6), A2 => n127, ZN => n157);
   U103 : OR2_X1 port map( A1 => n177, A2 => b(6), ZN => n158);
   U104 : OR2_X1 port map( A1 => b(7), A2 => a(7), ZN => n159);
   U105 : NAND3_X1 port map( A1 => n157, A2 => n158, A3 => n159, ZN => n178);
   U106 : OR2_X1 port map( A1 => n198, A2 => n197, ZN => n160);
   U107 : NAND2_X1 port map( A1 => n196, A2 => n160, ZN => n241);
   U108 : INV_X1 port map( A => a(15), ZN => n197);
   U109 : OAI22_X1 port map( A1 => a(22), A2 => n217, B1 => b(22), B2 => n216, 
                           ZN => n221);
   U110 : INV_X1 port map( A => a(23), ZN => n220);
   U111 : OAI22_X1 port map( A1 => b(0), A2 => a(0), B1 => cin, B2 => n165, ZN 
                           => n166);
   U112 : AND2_X1 port map( A1 => a(0), A2 => b(0), ZN => n165);
   U113 : AND2_X1 port map( A1 => n244, A2 => a(4), ZN => n175);
   U114 : OAI222_X1 port map( A1 => a(20), A2 => cout_4_port, B1 => b(20), B2 
                           => n212, C1 => b(21), C2 => a(21), ZN => n213);
   U115 : AND2_X1 port map( A1 => n155, A2 => a(28), ZN => n230);
   U116 : NAND2_X1 port map( A1 => n243, A2 => a(8), ZN => n184);
   U117 : OAI21_X1 port map( B1 => n128, B2 => a(15), A => b(15), ZN => n196);
   U118 : AND2_X1 port map( A1 => n126, A2 => a(6), ZN => n177);
   U119 : AOI22_X1 port map( A1 => b(26), A2 => a(26), B1 => n227, B2 => n228, 
                           ZN => n229);
   U120 : INV_X1 port map( A => n147, ZN => n173);
   U121 : AND2_X1 port map( A1 => n242, A2 => a(12), ZN => n194);
   U122 : OAI21_X1 port map( B1 => n243, B2 => a(8), A => b(8), ZN => n183);
   U123 : AND2_X1 port map( A1 => cout_4_port, A2 => a(20), ZN => n212);
   U124 : OAI221_X4 port map( B1 => n211, B2 => n210, C1 => n209, C2 => n208, A
                           => n207, ZN => cout_4_port);
   U125 : OAI22_X1 port map( A1 => n226, A2 => n225, B1 => n224, B2 => n223, ZN
                           => n227);
   U126 : AOI22_X1 port map( A1 => b(24), A2 => n222, B1 => a(24), B2 => n240, 
                           ZN => n226);
   U127 : OAI22_X1 port map( A1 => a(2), A2 => n170, B1 => n133, B2 => b(2), ZN
                           => n171);
   U128 : OAI21_X1 port map( B1 => n218, B2 => a(23), A => b(23), ZN => n219);
   U129 : OAI211_X1 port map( C1 => b(16), C2 => a(16), A => n241, B => n199, 
                           ZN => n211);

end SYN_p4_carry_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AddSub_DATA_SIZE32_3 is

   port( as : in std_logic;  a, b : in std_logic_vector (31 downto 0);  re : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end AddSub_DATA_SIZE32_3;

architecture SYN_add_sub_arch of AddSub_DATA_SIZE32_3 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component Adder_DATA_SIZE32_3
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;
   
   signal b_new_31_port, b_new_30_port, b_new_29_port, b_new_28_port, 
      b_new_27_port, b_new_26_port, b_new_25_port, b_new_24_port, b_new_23_port
      , b_new_22_port, b_new_21_port, b_new_20_port, b_new_19_port, 
      b_new_18_port, b_new_17_port, b_new_16_port, b_new_15_port, b_new_14_port
      , b_new_13_port, b_new_12_port, b_new_11_port, b_new_10_port, 
      b_new_9_port, b_new_8_port, b_new_7_port, b_new_6_port, b_new_5_port, 
      b_new_4_port, b_new_3_port, b_new_2_port, b_new_1_port, b_new_0_port, n1 
      : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b(9), B => n1, Z => b_new_9_port);
   U2 : XOR2_X1 port map( A => b(8), B => n1, Z => b_new_8_port);
   U3 : XOR2_X1 port map( A => b(7), B => n1, Z => b_new_7_port);
   U4 : XOR2_X1 port map( A => b(6), B => n1, Z => b_new_6_port);
   U5 : XOR2_X1 port map( A => b(5), B => n1, Z => b_new_5_port);
   U6 : XOR2_X1 port map( A => b(4), B => n1, Z => b_new_4_port);
   U7 : XOR2_X1 port map( A => b(3), B => n1, Z => b_new_3_port);
   U8 : XOR2_X1 port map( A => b(31), B => n1, Z => b_new_31_port);
   U9 : XOR2_X1 port map( A => b(30), B => n1, Z => b_new_30_port);
   U10 : XOR2_X1 port map( A => b(2), B => n1, Z => b_new_2_port);
   U11 : XOR2_X1 port map( A => b(29), B => n1, Z => b_new_29_port);
   U12 : XOR2_X1 port map( A => b(28), B => n1, Z => b_new_28_port);
   U13 : XOR2_X1 port map( A => b(27), B => n1, Z => b_new_27_port);
   U14 : XOR2_X1 port map( A => b(26), B => n1, Z => b_new_26_port);
   U15 : XOR2_X1 port map( A => b(25), B => n1, Z => b_new_25_port);
   U16 : XOR2_X1 port map( A => b(24), B => n1, Z => b_new_24_port);
   U17 : XOR2_X1 port map( A => b(23), B => n1, Z => b_new_23_port);
   U18 : XOR2_X1 port map( A => b(22), B => n1, Z => b_new_22_port);
   U19 : XOR2_X1 port map( A => b(21), B => n1, Z => b_new_21_port);
   U20 : XOR2_X1 port map( A => b(20), B => n1, Z => b_new_20_port);
   U21 : XOR2_X1 port map( A => b(1), B => n1, Z => b_new_1_port);
   U22 : XOR2_X1 port map( A => b(19), B => n1, Z => b_new_19_port);
   U23 : XOR2_X1 port map( A => b(18), B => n1, Z => b_new_18_port);
   U24 : XOR2_X1 port map( A => b(17), B => n1, Z => b_new_17_port);
   U25 : XOR2_X1 port map( A => b(16), B => n1, Z => b_new_16_port);
   U26 : XOR2_X1 port map( A => b(15), B => n1, Z => b_new_15_port);
   U27 : XOR2_X1 port map( A => b(14), B => n1, Z => b_new_14_port);
   U28 : XOR2_X1 port map( A => b(13), B => n1, Z => b_new_13_port);
   U29 : XOR2_X1 port map( A => b(12), B => n1, Z => b_new_12_port);
   U30 : XOR2_X1 port map( A => b(11), B => n1, Z => b_new_11_port);
   U31 : XOR2_X1 port map( A => b(10), B => n1, Z => b_new_10_port);
   ADDER0 : Adder_DATA_SIZE32_3 port map( cin => n1, a(31) => a(31), a(30) => 
                           a(30), a(29) => a(29), a(28) => a(28), a(27) => 
                           a(27), a(26) => a(26), a(25) => a(25), a(24) => 
                           a(24), a(23) => a(23), a(22) => a(22), a(21) => 
                           a(21), a(20) => a(20), a(19) => a(19), a(18) => 
                           a(18), a(17) => a(17), a(16) => a(16), a(15) => 
                           a(15), a(14) => a(14), a(13) => a(13), a(12) => 
                           a(12), a(11) => a(11), a(10) => a(10), a(9) => a(9),
                           a(8) => a(8), a(7) => a(7), a(6) => a(6), a(5) => 
                           a(5), a(4) => a(4), a(3) => a(3), a(2) => a(2), a(1)
                           => a(1), a(0) => a(0), b(31) => b_new_31_port, b(30)
                           => b_new_30_port, b(29) => b_new_29_port, b(28) => 
                           b_new_28_port, b(27) => b_new_27_port, b(26) => 
                           b_new_26_port, b(25) => b_new_25_port, b(24) => 
                           b_new_24_port, b(23) => b_new_23_port, b(22) => 
                           b_new_22_port, b(21) => b_new_21_port, b(20) => 
                           b_new_20_port, b(19) => b_new_19_port, b(18) => 
                           b_new_18_port, b(17) => b_new_17_port, b(16) => 
                           b_new_16_port, b(15) => b_new_15_port, b(14) => 
                           b_new_14_port, b(13) => b_new_13_port, b(12) => 
                           b_new_12_port, b(11) => b_new_11_port, b(10) => 
                           b_new_10_port, b(9) => b_new_9_port, b(8) => 
                           b_new_8_port, b(7) => b_new_7_port, b(6) => 
                           b_new_6_port, b(5) => b_new_5_port, b(4) => 
                           b_new_4_port, b(3) => b_new_3_port, b(2) => 
                           b_new_2_port, b(1) => b_new_1_port, b(0) => 
                           b_new_0_port, s(31) => re(31), s(30) => re(30), 
                           s(29) => re(29), s(28) => re(28), s(27) => re(27), 
                           s(26) => re(26), s(25) => re(25), s(24) => re(24), 
                           s(23) => re(23), s(22) => re(22), s(21) => re(21), 
                           s(20) => re(20), s(19) => re(19), s(18) => re(18), 
                           s(17) => re(17), s(16) => re(16), s(15) => re(15), 
                           s(14) => re(14), s(13) => re(13), s(12) => re(12), 
                           s(11) => re(11), s(10) => re(10), s(9) => re(9), 
                           s(8) => re(8), s(7) => re(7), s(6) => re(6), s(5) =>
                           re(5), s(4) => re(4), s(3) => re(3), s(2) => re(2), 
                           s(1) => re(1), s(0) => re(0), cout => cout);
   U32 : BUF_X4 port map( A => as, Z => n1);
   U33 : XOR2_X1 port map( A => b(0), B => as, Z => b_new_0_port);

end SYN_add_sub_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AddSub_DATA_SIZE32_2 is

   port( as : in std_logic;  a, b : in std_logic_vector (31 downto 0);  re : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end AddSub_DATA_SIZE32_2;

architecture SYN_add_sub_arch of AddSub_DATA_SIZE32_2 is

   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component Adder_DATA_SIZE32_2
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal b_new_31_port, b_new_30_port, b_new_29_port, b_new_28_port, 
      b_new_27_port, b_new_26_port, b_new_25_port, b_new_24_port, b_new_23_port
      , b_new_22_port, b_new_21_port, b_new_20_port, b_new_19_port, 
      b_new_18_port, b_new_17_port, b_new_16_port, b_new_15_port, b_new_14_port
      , b_new_13_port, b_new_12_port, b_new_11_port, b_new_10_port, 
      b_new_9_port, b_new_8_port, b_new_7_port, b_new_6_port, b_new_5_port, 
      b_new_4_port, b_new_3_port, b_new_2_port, b_new_1_port, b_new_0_port, n1,
      n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b(9), B => n5, Z => b_new_9_port);
   U2 : XOR2_X1 port map( A => b(8), B => n5, Z => b_new_8_port);
   U3 : XOR2_X1 port map( A => b(7), B => n5, Z => b_new_7_port);
   U4 : XOR2_X1 port map( A => b(6), B => n5, Z => b_new_6_port);
   U5 : XOR2_X1 port map( A => b(5), B => n5, Z => b_new_5_port);
   U6 : XOR2_X1 port map( A => b(4), B => n5, Z => b_new_4_port);
   U7 : XOR2_X1 port map( A => b(3), B => n5, Z => b_new_3_port);
   U8 : XOR2_X1 port map( A => b(31), B => n5, Z => b_new_31_port);
   U9 : XOR2_X1 port map( A => b(30), B => n5, Z => b_new_30_port);
   U10 : XOR2_X1 port map( A => b(2), B => n5, Z => b_new_2_port);
   U11 : XOR2_X1 port map( A => b(29), B => n5, Z => b_new_29_port);
   U12 : XOR2_X1 port map( A => b(28), B => n5, Z => b_new_28_port);
   U13 : XOR2_X1 port map( A => b(27), B => n5, Z => b_new_27_port);
   U14 : XOR2_X1 port map( A => b(26), B => n5, Z => b_new_26_port);
   U15 : XOR2_X1 port map( A => b(25), B => n5, Z => b_new_25_port);
   U16 : XOR2_X1 port map( A => b(24), B => n5, Z => b_new_24_port);
   U17 : XOR2_X1 port map( A => b(23), B => n5, Z => b_new_23_port);
   U18 : XOR2_X1 port map( A => b(22), B => n5, Z => b_new_22_port);
   U19 : XOR2_X1 port map( A => b(21), B => n5, Z => b_new_21_port);
   U20 : XOR2_X1 port map( A => b(20), B => n5, Z => b_new_20_port);
   U21 : XOR2_X1 port map( A => b(1), B => n5, Z => b_new_1_port);
   U22 : XOR2_X1 port map( A => b(19), B => n5, Z => b_new_19_port);
   U23 : XOR2_X1 port map( A => b(18), B => n5, Z => b_new_18_port);
   U24 : XOR2_X1 port map( A => b(17), B => n5, Z => b_new_17_port);
   U25 : XOR2_X1 port map( A => b(16), B => n5, Z => b_new_16_port);
   U26 : XOR2_X1 port map( A => b(15), B => n5, Z => b_new_15_port);
   U27 : XOR2_X1 port map( A => b(14), B => n5, Z => b_new_14_port);
   U28 : XOR2_X1 port map( A => b(13), B => n6, Z => b_new_13_port);
   U29 : XOR2_X1 port map( A => b(12), B => n6, Z => b_new_12_port);
   U30 : XOR2_X1 port map( A => b(11), B => n6, Z => b_new_11_port);
   U31 : XOR2_X1 port map( A => b(10), B => n6, Z => b_new_10_port);
   ADDER0 : Adder_DATA_SIZE32_2 port map( cin => n5, a(31) => a(31), a(30) => 
                           a(30), a(29) => a(29), a(28) => a(28), a(27) => 
                           a(27), a(26) => a(26), a(25) => a(25), a(24) => 
                           a(24), a(23) => a(23), a(22) => a(22), a(21) => 
                           a(21), a(20) => a(20), a(19) => a(19), a(18) => 
                           a(18), a(17) => a(17), a(16) => a(16), a(15) => 
                           a(15), a(14) => a(14), a(13) => a(13), a(12) => 
                           a(12), a(11) => a(11), a(10) => a(10), a(9) => a(9),
                           a(8) => a(8), a(7) => a(7), a(6) => a(6), a(5) => 
                           a(5), a(4) => a(4), a(3) => a(3), a(2) => a(2), a(1)
                           => a(1), a(0) => a(0), b(31) => b_new_31_port, b(30)
                           => b_new_30_port, b(29) => b_new_29_port, b(28) => 
                           b_new_28_port, b(27) => b_new_27_port, b(26) => 
                           b_new_26_port, b(25) => b_new_25_port, b(24) => 
                           b_new_24_port, b(23) => b_new_23_port, b(22) => 
                           b_new_22_port, b(21) => b_new_21_port, b(20) => 
                           b_new_20_port, b(19) => b_new_19_port, b(18) => 
                           b_new_18_port, b(17) => b_new_17_port, b(16) => 
                           b_new_16_port, b(15) => b_new_15_port, b(14) => 
                           b_new_14_port, b(13) => b_new_13_port, b(12) => 
                           b_new_12_port, b(11) => b_new_11_port, b(10) => 
                           b_new_10_port, b(9) => b_new_9_port, b(8) => 
                           b_new_8_port, b(7) => b_new_7_port, b(6) => 
                           b_new_6_port, b(5) => b_new_5_port, b(4) => 
                           b_new_4_port, b(3) => b_new_3_port, b(2) => 
                           b_new_2_port, b(1) => b_new_1_port, b(0) => 
                           b_new_0_port, s(31) => re(31), s(30) => re(30), 
                           s(29) => re(29), s(28) => re(28), s(27) => re(27), 
                           s(26) => re(26), s(25) => re(25), s(24) => re(24), 
                           s(23) => re(23), s(22) => re(22), s(21) => re(21), 
                           s(20) => re(20), s(19) => re(19), s(18) => re(18), 
                           s(17) => re(17), s(16) => re(16), s(15) => re(15), 
                           s(14) => re(14), s(13) => re(13), s(12) => re(12), 
                           s(11) => re(11), s(10) => re(10), s(9) => re(9), 
                           s(8) => re(8), s(7) => re(7), s(6) => re(6), s(5) =>
                           re(5), s(4) => re(4), s(3) => re(3), s(2) => re(2), 
                           s(1) => re(1), s(0) => re(0), cout => cout);
   U32 : BUF_X2 port map( A => as, Z => n6);
   U33 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => b_new_0_port);
   U34 : NAND2_X1 port map( A1 => b(0), A2 => n2, ZN => n3);
   U35 : NAND2_X1 port map( A1 => n1, A2 => n6, ZN => n4);
   U36 : INV_X1 port map( A => b(0), ZN => n1);
   U37 : INV_X1 port map( A => n6, ZN => n2);
   U38 : BUF_X4 port map( A => as, Z => n5);

end SYN_add_sub_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AddSub_DATA_SIZE32_1 is

   port( as : in std_logic;  a, b : in std_logic_vector (31 downto 0);  re : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end AddSub_DATA_SIZE32_1;

architecture SYN_add_sub_arch of AddSub_DATA_SIZE32_1 is

   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component Adder_DATA_SIZE32_1
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal b_new_31_port, b_new_30_port, b_new_29_port, b_new_28_port, 
      b_new_27_port, b_new_26_port, b_new_25_port, b_new_24_port, b_new_23_port
      , b_new_22_port, b_new_21_port, b_new_20_port, b_new_19_port, 
      b_new_18_port, b_new_17_port, b_new_16_port, b_new_15_port, b_new_14_port
      , b_new_13_port, b_new_12_port, b_new_11_port, b_new_10_port, 
      b_new_9_port, b_new_8_port, b_new_7_port, b_new_6_port, b_new_5_port, 
      b_new_4_port, b_new_3_port, b_new_2_port, b_new_1_port, b_new_0_port, n1,
      n2, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b(9), B => n5, Z => b_new_9_port);
   U2 : XOR2_X1 port map( A => b(8), B => n5, Z => b_new_8_port);
   U3 : XOR2_X1 port map( A => b(7), B => n5, Z => b_new_7_port);
   U4 : XOR2_X1 port map( A => b(6), B => n5, Z => b_new_6_port);
   U5 : XOR2_X1 port map( A => b(5), B => n5, Z => b_new_5_port);
   U6 : XOR2_X1 port map( A => b(4), B => n5, Z => b_new_4_port);
   U7 : XOR2_X1 port map( A => b(3), B => n5, Z => b_new_3_port);
   U8 : XOR2_X1 port map( A => b(31), B => n5, Z => b_new_31_port);
   U9 : XOR2_X1 port map( A => b(30), B => n5, Z => b_new_30_port);
   U10 : XOR2_X1 port map( A => b(2), B => n5, Z => b_new_2_port);
   U11 : XOR2_X1 port map( A => b(29), B => n5, Z => b_new_29_port);
   U12 : XOR2_X1 port map( A => b(28), B => n5, Z => b_new_28_port);
   U13 : XOR2_X1 port map( A => b(27), B => n5, Z => b_new_27_port);
   U14 : XOR2_X1 port map( A => b(26), B => n5, Z => b_new_26_port);
   U15 : XOR2_X1 port map( A => b(25), B => n5, Z => b_new_25_port);
   U16 : XOR2_X1 port map( A => b(24), B => n5, Z => b_new_24_port);
   U17 : XOR2_X1 port map( A => b(23), B => n5, Z => b_new_23_port);
   U18 : XOR2_X1 port map( A => b(22), B => n5, Z => b_new_22_port);
   U19 : XOR2_X1 port map( A => b(21), B => n5, Z => b_new_21_port);
   U20 : XOR2_X1 port map( A => b(20), B => n5, Z => b_new_20_port);
   U21 : XOR2_X1 port map( A => b(1), B => n5, Z => b_new_1_port);
   U22 : XOR2_X1 port map( A => b(19), B => n5, Z => b_new_19_port);
   U23 : XOR2_X1 port map( A => b(18), B => n5, Z => b_new_18_port);
   U24 : XOR2_X1 port map( A => b(17), B => n5, Z => b_new_17_port);
   U25 : XOR2_X1 port map( A => b(16), B => n5, Z => b_new_16_port);
   U26 : XOR2_X1 port map( A => b(15), B => n5, Z => b_new_15_port);
   U27 : XOR2_X1 port map( A => b(14), B => n5, Z => b_new_14_port);
   U28 : XOR2_X1 port map( A => b(13), B => n6, Z => b_new_13_port);
   U29 : XOR2_X1 port map( A => b(12), B => n6, Z => b_new_12_port);
   U30 : XOR2_X1 port map( A => b(11), B => n6, Z => b_new_11_port);
   U31 : XOR2_X1 port map( A => b(10), B => n6, Z => b_new_10_port);
   ADDER0 : Adder_DATA_SIZE32_1 port map( cin => n5, a(31) => a(31), a(30) => 
                           a(30), a(29) => a(29), a(28) => a(28), a(27) => 
                           a(27), a(26) => a(26), a(25) => a(25), a(24) => 
                           a(24), a(23) => a(23), a(22) => a(22), a(21) => 
                           a(21), a(20) => a(20), a(19) => a(19), a(18) => 
                           a(18), a(17) => a(17), a(16) => a(16), a(15) => 
                           a(15), a(14) => a(14), a(13) => a(13), a(12) => 
                           a(12), a(11) => a(11), a(10) => a(10), a(9) => a(9),
                           a(8) => a(8), a(7) => a(7), a(6) => a(6), a(5) => 
                           a(5), a(4) => a(4), a(3) => a(3), a(2) => a(2), a(1)
                           => a(1), a(0) => a(0), b(31) => b_new_31_port, b(30)
                           => b_new_30_port, b(29) => b_new_29_port, b(28) => 
                           b_new_28_port, b(27) => b_new_27_port, b(26) => 
                           b_new_26_port, b(25) => b_new_25_port, b(24) => 
                           b_new_24_port, b(23) => b_new_23_port, b(22) => 
                           b_new_22_port, b(21) => b_new_21_port, b(20) => 
                           b_new_20_port, b(19) => b_new_19_port, b(18) => 
                           b_new_18_port, b(17) => b_new_17_port, b(16) => 
                           b_new_16_port, b(15) => b_new_15_port, b(14) => 
                           b_new_14_port, b(13) => b_new_13_port, b(12) => 
                           b_new_12_port, b(11) => b_new_11_port, b(10) => 
                           b_new_10_port, b(9) => b_new_9_port, b(8) => 
                           b_new_8_port, b(7) => b_new_7_port, b(6) => 
                           b_new_6_port, b(5) => b_new_5_port, b(4) => 
                           b_new_4_port, b(3) => b_new_3_port, b(2) => 
                           b_new_2_port, b(1) => b_new_1_port, b(0) => 
                           b_new_0_port, s(31) => re(31), s(30) => re(30), 
                           s(29) => re(29), s(28) => re(28), s(27) => re(27), 
                           s(26) => re(26), s(25) => re(25), s(24) => re(24), 
                           s(23) => re(23), s(22) => re(22), s(21) => re(21), 
                           s(20) => re(20), s(19) => re(19), s(18) => re(18), 
                           s(17) => re(17), s(16) => re(16), s(15) => re(15), 
                           s(14) => re(14), s(13) => re(13), s(12) => re(12), 
                           s(11) => re(11), s(10) => re(10), s(9) => re(9), 
                           s(8) => re(8), s(7) => re(7), s(6) => re(6), s(5) =>
                           re(5), s(4) => re(4), s(3) => re(3), s(2) => re(2), 
                           s(1) => re(1), s(0) => re(0), cout => cout);
   U32 : BUF_X1 port map( A => as, Z => n6);
   U33 : NAND2_X1 port map( A1 => b(0), A2 => n2, ZN => n3);
   U34 : NAND2_X1 port map( A1 => n1, A2 => n6, ZN => n4);
   U35 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => b_new_0_port);
   U36 : INV_X1 port map( A => b(0), ZN => n1);
   U37 : INV_X1 port map( A => n6, ZN => n2);
   U38 : BUF_X4 port map( A => as, Z => n5);

end SYN_add_sub_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4Adder_DATA_SIZE32_SPARSITY4_7 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end P4Adder_DATA_SIZE32_SPARSITY4_7;

architecture SYN_p4_adder_arch of P4Adder_DATA_SIZE32_SPARSITY4_7 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AdderSumGenerator_DATA_SIZE32_SPARSITY4_7
      port( a, b : in std_logic_vector (31 downto 0);  cin : in 
            std_logic_vector (7 downto 0);  sum : out std_logic_vector (31 
            downto 0));
   end component;
   
   component P4CarryGenerator_DATA_SIZE32_SPARSITY4_7
      port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  
            cout : out std_logic_vector (7 downto 0));
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, carry_1_port, n1, n2 : std_logic;

begin
   
   CG0 : P4CarryGenerator_DATA_SIZE32_SPARSITY4_7 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), cin => cin, 
                           cout(7) => cout, cout(6) => carry_7_port, cout(5) =>
                           carry_6_port, cout(4) => carry_5_port, cout(3) => 
                           carry_4_port, cout(2) => carry_3_port, cout(1) => 
                           carry_2_port, cout(0) => carry_1_port);
   SG0 : AdderSumGenerator_DATA_SIZE32_SPARSITY4_7 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => n1, b(0) => n2, cin(7) => carry_7_port
                           , cin(6) => carry_6_port, cin(5) => carry_5_port, 
                           cin(4) => carry_4_port, cin(3) => carry_3_port, 
                           cin(2) => carry_2_port, cin(1) => carry_1_port, 
                           cin(0) => cin, sum(31) => s(31), sum(30) => s(30), 
                           sum(29) => s(29), sum(28) => s(28), sum(27) => s(27)
                           , sum(26) => s(26), sum(25) => s(25), sum(24) => 
                           s(24), sum(23) => s(23), sum(22) => s(22), sum(21) 
                           => s(21), sum(20) => s(20), sum(19) => s(19), 
                           sum(18) => s(18), sum(17) => s(17), sum(16) => s(16)
                           , sum(15) => s(15), sum(14) => s(14), sum(13) => 
                           s(13), sum(12) => s(12), sum(11) => s(11), sum(10) 
                           => s(10), sum(9) => s(9), sum(8) => s(8), sum(7) => 
                           s(7), sum(6) => s(6), sum(5) => s(5), sum(4) => s(4)
                           , sum(3) => s(3), sum(2) => s(2), sum(1) => s(1), 
                           sum(0) => s(0));
   U1 : CLKBUF_X1 port map( A => b(1), Z => n1);
   U2 : CLKBUF_X1 port map( A => b(0), Z => n2);

end SYN_p4_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4Adder_DATA_SIZE32_SPARSITY4_6 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end P4Adder_DATA_SIZE32_SPARSITY4_6;

architecture SYN_p4_adder_arch of P4Adder_DATA_SIZE32_SPARSITY4_6 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AdderSumGenerator_DATA_SIZE32_SPARSITY4_6
      port( a, b : in std_logic_vector (31 downto 0);  cin : in 
            std_logic_vector (7 downto 0);  sum : out std_logic_vector (31 
            downto 0));
   end component;
   
   component P4CarryGenerator_DATA_SIZE32_SPARSITY4_6
      port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  
            cout : out std_logic_vector (7 downto 0));
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, carry_1_port, n1, n2 : std_logic;

begin
   
   CG0 : P4CarryGenerator_DATA_SIZE32_SPARSITY4_6 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), cin => cin, 
                           cout(7) => cout, cout(6) => carry_7_port, cout(5) =>
                           carry_6_port, cout(4) => carry_5_port, cout(3) => 
                           carry_4_port, cout(2) => carry_3_port, cout(1) => 
                           carry_2_port, cout(0) => carry_1_port);
   SG0 : AdderSumGenerator_DATA_SIZE32_SPARSITY4_6 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => n1, b(0) => n2, cin(7) => carry_7_port
                           , cin(6) => carry_6_port, cin(5) => carry_5_port, 
                           cin(4) => carry_4_port, cin(3) => carry_3_port, 
                           cin(2) => carry_2_port, cin(1) => carry_1_port, 
                           cin(0) => cin, sum(31) => s(31), sum(30) => s(30), 
                           sum(29) => s(29), sum(28) => s(28), sum(27) => s(27)
                           , sum(26) => s(26), sum(25) => s(25), sum(24) => 
                           s(24), sum(23) => s(23), sum(22) => s(22), sum(21) 
                           => s(21), sum(20) => s(20), sum(19) => s(19), 
                           sum(18) => s(18), sum(17) => s(17), sum(16) => s(16)
                           , sum(15) => s(15), sum(14) => s(14), sum(13) => 
                           s(13), sum(12) => s(12), sum(11) => s(11), sum(10) 
                           => s(10), sum(9) => s(9), sum(8) => s(8), sum(7) => 
                           s(7), sum(6) => s(6), sum(5) => s(5), sum(4) => s(4)
                           , sum(3) => s(3), sum(2) => s(2), sum(1) => s(1), 
                           sum(0) => s(0));
   U1 : CLKBUF_X1 port map( A => b(1), Z => n1);
   U2 : CLKBUF_X1 port map( A => b(0), Z => n2);

end SYN_p4_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4Adder_DATA_SIZE32_SPARSITY4_5 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end P4Adder_DATA_SIZE32_SPARSITY4_5;

architecture SYN_p4_adder_arch of P4Adder_DATA_SIZE32_SPARSITY4_5 is

   component AdderSumGenerator_DATA_SIZE32_SPARSITY4_5
      port( a, b : in std_logic_vector (31 downto 0);  cin : in 
            std_logic_vector (7 downto 0);  sum : out std_logic_vector (31 
            downto 0));
   end component;
   
   component P4CarryGenerator_DATA_SIZE32_SPARSITY4_5
      port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  
            cout : out std_logic_vector (7 downto 0));
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, carry_1_port : std_logic;

begin
   
   CG0 : P4CarryGenerator_DATA_SIZE32_SPARSITY4_5 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), cin => cin, 
                           cout(7) => cout, cout(6) => carry_7_port, cout(5) =>
                           carry_6_port, cout(4) => carry_5_port, cout(3) => 
                           carry_4_port, cout(2) => carry_3_port, cout(1) => 
                           carry_2_port, cout(0) => carry_1_port);
   SG0 : AdderSumGenerator_DATA_SIZE32_SPARSITY4_5 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), cin(7) => 
                           carry_7_port, cin(6) => carry_6_port, cin(5) => 
                           carry_5_port, cin(4) => carry_4_port, cin(3) => 
                           carry_3_port, cin(2) => carry_2_port, cin(1) => 
                           carry_1_port, cin(0) => cin, sum(31) => s(31), 
                           sum(30) => s(30), sum(29) => s(29), sum(28) => s(28)
                           , sum(27) => s(27), sum(26) => s(26), sum(25) => 
                           s(25), sum(24) => s(24), sum(23) => s(23), sum(22) 
                           => s(22), sum(21) => s(21), sum(20) => s(20), 
                           sum(19) => s(19), sum(18) => s(18), sum(17) => s(17)
                           , sum(16) => s(16), sum(15) => s(15), sum(14) => 
                           s(14), sum(13) => s(13), sum(12) => s(12), sum(11) 
                           => s(11), sum(10) => s(10), sum(9) => s(9), sum(8) 
                           => s(8), sum(7) => s(7), sum(6) => s(6), sum(5) => 
                           s(5), sum(4) => s(4), sum(3) => s(3), sum(2) => s(2)
                           , sum(1) => s(1), sum(0) => s(0));

end SYN_p4_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4Adder_DATA_SIZE32_SPARSITY4_4 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end P4Adder_DATA_SIZE32_SPARSITY4_4;

architecture SYN_p4_adder_arch of P4Adder_DATA_SIZE32_SPARSITY4_4 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AdderSumGenerator_DATA_SIZE32_SPARSITY4_4
      port( a, b : in std_logic_vector (31 downto 0);  cin : in 
            std_logic_vector (7 downto 0);  sum : out std_logic_vector (31 
            downto 0));
   end component;
   
   component P4CarryGenerator_DATA_SIZE32_SPARSITY4_4
      port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  
            cout : out std_logic_vector (7 downto 0));
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, carry_1_port, n1 : std_logic;

begin
   
   CG0 : P4CarryGenerator_DATA_SIZE32_SPARSITY4_4 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), cin => cin, 
                           cout(7) => cout, cout(6) => carry_7_port, cout(5) =>
                           carry_6_port, cout(4) => carry_5_port, cout(3) => 
                           carry_4_port, cout(2) => carry_3_port, cout(1) => 
                           carry_2_port, cout(0) => carry_1_port);
   SG0 : AdderSumGenerator_DATA_SIZE32_SPARSITY4_4 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => n1, cin(7) => 
                           carry_7_port, cin(6) => carry_6_port, cin(5) => 
                           carry_5_port, cin(4) => carry_4_port, cin(3) => 
                           carry_3_port, cin(2) => carry_2_port, cin(1) => 
                           carry_1_port, cin(0) => cin, sum(31) => s(31), 
                           sum(30) => s(30), sum(29) => s(29), sum(28) => s(28)
                           , sum(27) => s(27), sum(26) => s(26), sum(25) => 
                           s(25), sum(24) => s(24), sum(23) => s(23), sum(22) 
                           => s(22), sum(21) => s(21), sum(20) => s(20), 
                           sum(19) => s(19), sum(18) => s(18), sum(17) => s(17)
                           , sum(16) => s(16), sum(15) => s(15), sum(14) => 
                           s(14), sum(13) => s(13), sum(12) => s(12), sum(11) 
                           => s(11), sum(10) => s(10), sum(9) => s(9), sum(8) 
                           => s(8), sum(7) => s(7), sum(6) => s(6), sum(5) => 
                           s(5), sum(4) => s(4), sum(3) => s(3), sum(2) => s(2)
                           , sum(1) => s(1), sum(0) => s(0));
   U1 : CLKBUF_X1 port map( A => b(0), Z => n1);

end SYN_p4_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4Adder_DATA_SIZE32_SPARSITY4_3 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end P4Adder_DATA_SIZE32_SPARSITY4_3;

architecture SYN_p4_adder_arch of P4Adder_DATA_SIZE32_SPARSITY4_3 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AdderSumGenerator_DATA_SIZE32_SPARSITY4_3
      port( a, b : in std_logic_vector (31 downto 0);  cin : in 
            std_logic_vector (7 downto 0);  sum : out std_logic_vector (31 
            downto 0));
   end component;
   
   component P4CarryGenerator_DATA_SIZE32_SPARSITY4_3
      port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  
            cout : out std_logic_vector (7 downto 0));
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, carry_1_port, n1, n2 : std_logic;

begin
   
   CG0 : P4CarryGenerator_DATA_SIZE32_SPARSITY4_3 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), cin => cin, 
                           cout(7) => cout, cout(6) => carry_7_port, cout(5) =>
                           carry_6_port, cout(4) => carry_5_port, cout(3) => 
                           carry_4_port, cout(2) => carry_3_port, cout(1) => 
                           carry_2_port, cout(0) => carry_1_port);
   SG0 : AdderSumGenerator_DATA_SIZE32_SPARSITY4_3 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => n1, b(0) => n2, cin(7) => carry_7_port
                           , cin(6) => carry_6_port, cin(5) => carry_5_port, 
                           cin(4) => carry_4_port, cin(3) => carry_3_port, 
                           cin(2) => carry_2_port, cin(1) => carry_1_port, 
                           cin(0) => cin, sum(31) => s(31), sum(30) => s(30), 
                           sum(29) => s(29), sum(28) => s(28), sum(27) => s(27)
                           , sum(26) => s(26), sum(25) => s(25), sum(24) => 
                           s(24), sum(23) => s(23), sum(22) => s(22), sum(21) 
                           => s(21), sum(20) => s(20), sum(19) => s(19), 
                           sum(18) => s(18), sum(17) => s(17), sum(16) => s(16)
                           , sum(15) => s(15), sum(14) => s(14), sum(13) => 
                           s(13), sum(12) => s(12), sum(11) => s(11), sum(10) 
                           => s(10), sum(9) => s(9), sum(8) => s(8), sum(7) => 
                           s(7), sum(6) => s(6), sum(5) => s(5), sum(4) => s(4)
                           , sum(3) => s(3), sum(2) => s(2), sum(1) => s(1), 
                           sum(0) => s(0));
   U1 : BUF_X1 port map( A => b(1), Z => n1);
   U2 : CLKBUF_X1 port map( A => b(0), Z => n2);

end SYN_p4_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4Adder_DATA_SIZE32_SPARSITY4_2 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end P4Adder_DATA_SIZE32_SPARSITY4_2;

architecture SYN_p4_adder_arch of P4Adder_DATA_SIZE32_SPARSITY4_2 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AdderSumGenerator_DATA_SIZE32_SPARSITY4_2
      port( a, b : in std_logic_vector (31 downto 0);  cin : in 
            std_logic_vector (7 downto 0);  sum : out std_logic_vector (31 
            downto 0));
   end component;
   
   component P4CarryGenerator_DATA_SIZE32_SPARSITY4_2
      port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  
            cout : out std_logic_vector (7 downto 0));
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, carry_1_port, n1 : std_logic;

begin
   
   CG0 : P4CarryGenerator_DATA_SIZE32_SPARSITY4_2 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), cin => cin, 
                           cout(7) => cout, cout(6) => carry_7_port, cout(5) =>
                           carry_6_port, cout(4) => carry_5_port, cout(3) => 
                           carry_4_port, cout(2) => carry_3_port, cout(1) => 
                           carry_2_port, cout(0) => carry_1_port);
   SG0 : AdderSumGenerator_DATA_SIZE32_SPARSITY4_2 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => n1, cin(7) => 
                           carry_7_port, cin(6) => carry_6_port, cin(5) => 
                           carry_5_port, cin(4) => carry_4_port, cin(3) => 
                           carry_3_port, cin(2) => carry_2_port, cin(1) => 
                           carry_1_port, cin(0) => cin, sum(31) => s(31), 
                           sum(30) => s(30), sum(29) => s(29), sum(28) => s(28)
                           , sum(27) => s(27), sum(26) => s(26), sum(25) => 
                           s(25), sum(24) => s(24), sum(23) => s(23), sum(22) 
                           => s(22), sum(21) => s(21), sum(20) => s(20), 
                           sum(19) => s(19), sum(18) => s(18), sum(17) => s(17)
                           , sum(16) => s(16), sum(15) => s(15), sum(14) => 
                           s(14), sum(13) => s(13), sum(12) => s(12), sum(11) 
                           => s(11), sum(10) => s(10), sum(9) => s(9), sum(8) 
                           => s(8), sum(7) => s(7), sum(6) => s(6), sum(5) => 
                           s(5), sum(4) => s(4), sum(3) => s(3), sum(2) => s(2)
                           , sum(1) => s(1), sum(0) => s(0));
   U1 : CLKBUF_X1 port map( A => b(0), Z => n1);

end SYN_p4_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4Adder_DATA_SIZE32_SPARSITY4_1 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end P4Adder_DATA_SIZE32_SPARSITY4_1;

architecture SYN_p4_adder_arch of P4Adder_DATA_SIZE32_SPARSITY4_1 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AdderSumGenerator_DATA_SIZE32_SPARSITY4_1
      port( a, b : in std_logic_vector (31 downto 0);  cin : in 
            std_logic_vector (7 downto 0);  sum : out std_logic_vector (31 
            downto 0));
   end component;
   
   component P4CarryGenerator_DATA_SIZE32_SPARSITY4_1
      port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  
            cout : out std_logic_vector (7 downto 0));
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, carry_1_port, n1, n2 : std_logic;

begin
   
   CG0 : P4CarryGenerator_DATA_SIZE32_SPARSITY4_1 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), cin => cin, 
                           cout(7) => cout, cout(6) => carry_7_port, cout(5) =>
                           carry_6_port, cout(4) => carry_5_port, cout(3) => 
                           carry_4_port, cout(2) => carry_3_port, cout(1) => 
                           carry_2_port, cout(0) => carry_1_port);
   SG0 : AdderSumGenerator_DATA_SIZE32_SPARSITY4_1 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => n1, b(0) => n2, cin(7) => carry_7_port
                           , cin(6) => carry_6_port, cin(5) => carry_5_port, 
                           cin(4) => carry_4_port, cin(3) => carry_3_port, 
                           cin(2) => carry_2_port, cin(1) => carry_1_port, 
                           cin(0) => cin, sum(31) => s(31), sum(30) => s(30), 
                           sum(29) => s(29), sum(28) => s(28), sum(27) => s(27)
                           , sum(26) => s(26), sum(25) => s(25), sum(24) => 
                           s(24), sum(23) => s(23), sum(22) => s(22), sum(21) 
                           => s(21), sum(20) => s(20), sum(19) => s(19), 
                           sum(18) => s(18), sum(17) => s(17), sum(16) => s(16)
                           , sum(15) => s(15), sum(14) => s(14), sum(13) => 
                           s(13), sum(12) => s(12), sum(11) => s(11), sum(10) 
                           => s(10), sum(9) => s(9), sum(8) => s(8), sum(7) => 
                           s(7), sum(6) => s(6), sum(5) => s(5), sum(4) => s(4)
                           , sum(3) => s(3), sum(2) => s(2), sum(1) => s(1), 
                           sum(0) => s(0));
   U1 : CLKBUF_X1 port map( A => b(1), Z => n1);
   U2 : CLKBUF_X1 port map( A => b(0), Z => n2);

end SYN_p4_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE5_5 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 0); 
         dout : out std_logic_vector (4 downto 0));

end Reg_DATA_SIZE5_5;

architecture SYN_reg_arch of Reg_DATA_SIZE5_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, net109193, net109194, net109195, net109196, 
      net109197, n11, n12, n13, n14, n15 : std_logic;

begin
   
   dout_reg_4_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           dout(4), QN => net109197);
   dout_reg_3_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           dout(3), QN => net109196);
   dout_reg_2_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           dout(2), QN => net109195);
   dout_reg_1_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           dout(1), QN => net109194);
   dout_reg_0_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           dout(0), QN => net109193);
   U2 : OAI21_X1 port map( B1 => net109193, B2 => en, A => n15, ZN => n5);
   U3 : NAND2_X1 port map( A1 => en, A2 => din(0), ZN => n15);
   U4 : OAI21_X1 port map( B1 => net109194, B2 => en, A => n14, ZN => n4);
   U5 : NAND2_X1 port map( A1 => din(1), A2 => en, ZN => n14);
   U6 : OAI21_X1 port map( B1 => net109195, B2 => en, A => n13, ZN => n3);
   U7 : NAND2_X1 port map( A1 => din(2), A2 => en, ZN => n13);
   U8 : OAI21_X1 port map( B1 => net109196, B2 => en, A => n12, ZN => n2);
   U9 : NAND2_X1 port map( A1 => din(3), A2 => en, ZN => n12);
   U10 : OAI21_X1 port map( B1 => net109197, B2 => en, A => n11, ZN => n1);
   U11 : NAND2_X1 port map( A1 => din(4), A2 => en, ZN => n11);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE5_4 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 0); 
         dout : out std_logic_vector (4 downto 0));

end Reg_DATA_SIZE5_4;

architecture SYN_reg_arch of Reg_DATA_SIZE5_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, net109193, net109194, net109195, net109196, 
      net109197, n11, n12, n13, n14, n15 : std_logic;

begin
   
   dout_reg_4_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           dout(4), QN => net109197);
   dout_reg_3_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           dout(3), QN => net109196);
   dout_reg_2_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           dout(2), QN => net109195);
   dout_reg_1_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           dout(1), QN => net109194);
   dout_reg_0_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           dout(0), QN => net109193);
   U2 : OAI21_X1 port map( B1 => net109193, B2 => en, A => n15, ZN => n5);
   U3 : NAND2_X1 port map( A1 => en, A2 => din(0), ZN => n15);
   U4 : OAI21_X1 port map( B1 => net109194, B2 => en, A => n14, ZN => n4);
   U5 : NAND2_X1 port map( A1 => din(1), A2 => en, ZN => n14);
   U6 : OAI21_X1 port map( B1 => net109195, B2 => en, A => n13, ZN => n3);
   U7 : NAND2_X1 port map( A1 => din(2), A2 => en, ZN => n13);
   U8 : OAI21_X1 port map( B1 => net109196, B2 => en, A => n12, ZN => n2);
   U9 : NAND2_X1 port map( A1 => din(3), A2 => en, ZN => n12);
   U10 : OAI21_X1 port map( B1 => net109197, B2 => en, A => n11, ZN => n1);
   U11 : NAND2_X1 port map( A1 => din(4), A2 => en, ZN => n11);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE5_3 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 0); 
         dout : out std_logic_vector (4 downto 0));

end Reg_DATA_SIZE5_3;

architecture SYN_reg_arch of Reg_DATA_SIZE5_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, net109193, net109194, net109195, net109196, 
      net109197, n11, n12, n13, n14, n15 : std_logic;

begin
   
   dout_reg_4_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           dout(4), QN => net109197);
   dout_reg_3_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           dout(3), QN => net109196);
   dout_reg_2_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           dout(2), QN => net109195);
   dout_reg_1_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           dout(1), QN => net109194);
   dout_reg_0_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           dout(0), QN => net109193);
   U2 : OAI21_X1 port map( B1 => net109193, B2 => en, A => n15, ZN => n5);
   U3 : NAND2_X1 port map( A1 => en, A2 => din(0), ZN => n15);
   U4 : OAI21_X1 port map( B1 => net109194, B2 => en, A => n14, ZN => n4);
   U5 : NAND2_X1 port map( A1 => din(1), A2 => en, ZN => n14);
   U6 : OAI21_X1 port map( B1 => net109195, B2 => en, A => n13, ZN => n3);
   U7 : NAND2_X1 port map( A1 => din(2), A2 => en, ZN => n13);
   U8 : OAI21_X1 port map( B1 => net109196, B2 => en, A => n12, ZN => n2);
   U9 : NAND2_X1 port map( A1 => din(3), A2 => en, ZN => n12);
   U10 : OAI21_X1 port map( B1 => net109197, B2 => en, A => n11, ZN => n1);
   U11 : NAND2_X1 port map( A1 => din(4), A2 => en, ZN => n11);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE5_2 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 0); 
         dout : out std_logic_vector (4 downto 0));

end Reg_DATA_SIZE5_2;

architecture SYN_reg_arch of Reg_DATA_SIZE5_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, net109193, net109194, net109195, net109196, 
      net109197, n11, n12, n13, n14, n15 : std_logic;

begin
   
   dout_reg_4_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           dout(4), QN => net109197);
   dout_reg_3_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           dout(3), QN => net109196);
   dout_reg_2_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           dout(2), QN => net109195);
   dout_reg_1_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           dout(1), QN => net109194);
   dout_reg_0_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           dout(0), QN => net109193);
   U2 : OAI21_X1 port map( B1 => net109193, B2 => en, A => n15, ZN => n5);
   U3 : NAND2_X1 port map( A1 => en, A2 => din(0), ZN => n15);
   U4 : OAI21_X1 port map( B1 => net109194, B2 => en, A => n14, ZN => n4);
   U5 : NAND2_X1 port map( A1 => din(1), A2 => en, ZN => n14);
   U6 : OAI21_X1 port map( B1 => net109195, B2 => en, A => n13, ZN => n3);
   U7 : NAND2_X1 port map( A1 => din(2), A2 => en, ZN => n13);
   U8 : OAI21_X1 port map( B1 => net109196, B2 => en, A => n12, ZN => n2);
   U9 : NAND2_X1 port map( A1 => din(3), A2 => en, ZN => n12);
   U10 : OAI21_X1 port map( B1 => net109197, B2 => en, A => n11, ZN => n1);
   U11 : NAND2_X1 port map( A1 => din(4), A2 => en, ZN => n11);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE5_1 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 0); 
         dout : out std_logic_vector (4 downto 0));

end Reg_DATA_SIZE5_1;

architecture SYN_reg_arch of Reg_DATA_SIZE5_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, net109193, net109194, net109195, net109196, 
      net109197, n11, n12, n13, n14, n15 : std_logic;

begin
   
   dout_reg_4_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           dout(4), QN => net109197);
   dout_reg_3_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           dout(3), QN => net109196);
   dout_reg_2_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           dout(2), QN => net109195);
   dout_reg_1_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           dout(1), QN => net109194);
   dout_reg_0_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           dout(0), QN => net109193);
   U2 : OAI21_X1 port map( B1 => net109193, B2 => en, A => n15, ZN => n5);
   U3 : NAND2_X1 port map( A1 => en, A2 => din(0), ZN => n15);
   U4 : OAI21_X1 port map( B1 => net109194, B2 => en, A => n14, ZN => n4);
   U5 : NAND2_X1 port map( A1 => din(1), A2 => en, ZN => n14);
   U6 : OAI21_X1 port map( B1 => net109195, B2 => en, A => n13, ZN => n3);
   U7 : NAND2_X1 port map( A1 => din(2), A2 => en, ZN => n13);
   U8 : OAI21_X1 port map( B1 => net109196, B2 => en, A => n12, ZN => n2);
   U9 : NAND2_X1 port map( A1 => din(3), A2 => en, ZN => n12);
   U10 : OAI21_X1 port map( B1 => net109197, B2 => en, A => n11, ZN => n1);
   U11 : NAND2_X1 port map( A1 => din(4), A2 => en, ZN => n11);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_2 is

   port( reg_c, reg_f, reg_ff : in std_logic_vector (31 downto 0);  addr_c, 
         addr_f, addr_ff : in std_logic_vector (4 downto 0);  valid_f, valid_ff
         , dirty_f, dirty_ff, en : in std_logic;  output : out std_logic_vector
         (31 downto 0);  match_dirty_f, match_dirty_ff : out std_logic);

end FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_2;

architecture SYN_fwd_mux_2_arch of FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
      N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, 
      N106, N107, N108, N109, N110, N111, N112, n92_port, n93_port, n94_port, 
      n95_port, n96_port, n97_port, n98_port, n99_port, n100_port, n101_port, 
      n102_port, n103_port, n104_port, n105_port, n106_port, n107_port, 
      n108_port, n109_port, n110_port, n111_port, n112_port, n113, n114, n115, 
      n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
      n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155 : std_logic;

begin
   
   match_dirty_ff_reg : DLH_X1 port map( G => en, D => N111, Q => 
                           match_dirty_ff);
   output_reg_31_inst : DLH_X1 port map( G => en, D => N110, Q => output(31));
   output_reg_30_inst : DLH_X1 port map( G => en, D => N109, Q => output(30));
   output_reg_29_inst : DLH_X1 port map( G => en, D => N108, Q => output(29));
   output_reg_28_inst : DLH_X1 port map( G => en, D => N107, Q => output(28));
   output_reg_27_inst : DLH_X1 port map( G => en, D => N106, Q => output(27));
   output_reg_26_inst : DLH_X1 port map( G => en, D => N105, Q => output(26));
   output_reg_25_inst : DLH_X1 port map( G => en, D => N104, Q => output(25));
   output_reg_24_inst : DLH_X1 port map( G => en, D => N103, Q => output(24));
   output_reg_23_inst : DLH_X1 port map( G => en, D => N102, Q => output(23));
   output_reg_22_inst : DLH_X1 port map( G => en, D => N101, Q => output(22));
   output_reg_21_inst : DLH_X1 port map( G => en, D => N100, Q => output(21));
   output_reg_20_inst : DLH_X1 port map( G => en, D => N99, Q => output(20));
   output_reg_19_inst : DLH_X1 port map( G => en, D => N98, Q => output(19));
   output_reg_18_inst : DLH_X1 port map( G => en, D => N97, Q => output(18));
   output_reg_17_inst : DLH_X1 port map( G => en, D => N96, Q => output(17));
   output_reg_16_inst : DLH_X1 port map( G => en, D => N95, Q => output(16));
   output_reg_15_inst : DLH_X1 port map( G => en, D => N94, Q => output(15));
   output_reg_14_inst : DLH_X1 port map( G => en, D => N93, Q => output(14));
   output_reg_13_inst : DLH_X1 port map( G => en, D => N92, Q => output(13));
   output_reg_12_inst : DLH_X1 port map( G => en, D => N91, Q => output(12));
   output_reg_11_inst : DLH_X1 port map( G => en, D => N90, Q => output(11));
   output_reg_10_inst : DLH_X1 port map( G => en, D => N89, Q => output(10));
   output_reg_9_inst : DLH_X1 port map( G => en, D => N88, Q => output(9));
   output_reg_8_inst : DLH_X1 port map( G => en, D => N87, Q => output(8));
   output_reg_7_inst : DLH_X1 port map( G => en, D => N86, Q => output(7));
   output_reg_6_inst : DLH_X1 port map( G => en, D => N85, Q => output(6));
   output_reg_5_inst : DLH_X1 port map( G => en, D => N84, Q => output(5));
   output_reg_4_inst : DLH_X1 port map( G => en, D => N83, Q => output(4));
   output_reg_3_inst : DLH_X1 port map( G => en, D => N82, Q => output(3));
   output_reg_2_inst : DLH_X1 port map( G => en, D => N81, Q => output(2));
   output_reg_1_inst : DLH_X1 port map( G => en, D => N80, Q => output(1));
   output_reg_0_inst : DLH_X1 port map( G => en, D => N79, Q => output(0));
   match_dirty_f_reg : DLH_X1 port map( G => en, D => N112, Q => match_dirty_f)
                           ;
   U83 : XOR2_X1 port map( A => addr_f(3), B => addr_c(3), Z => n107_port);
   U84 : XOR2_X1 port map( A => addr_f(2), B => addr_c(2), Z => n108_port);
   U85 : XOR2_X1 port map( A => addr_f(4), B => addr_c(4), Z => n109_port);
   U86 : XOR2_X1 port map( A => addr_ff(4), B => addr_c(4), Z => n101_port);
   U87 : XOR2_X1 port map( A => addr_ff(0), B => addr_c(0), Z => n102_port);
   U88 : XOR2_X1 port map( A => addr_ff(1), B => addr_c(1), Z => n103_port);
   U89 : XOR2_X1 port map( A => n116, B => addr_ff(3), Z => n105_port);
   U90 : XOR2_X1 port map( A => n114, B => addr_ff(2), Z => n106_port);
   U2 : BUF_X1 port map( A => n153, Z => n95_port);
   U3 : BUF_X1 port map( A => n153, Z => n96_port);
   U4 : BUF_X1 port map( A => n152, Z => n92_port);
   U5 : BUF_X1 port map( A => n152, Z => n93_port);
   U6 : BUF_X1 port map( A => n153, Z => n97_port);
   U7 : BUF_X1 port map( A => n154, Z => n99_port);
   U8 : BUF_X1 port map( A => n154, Z => n98_port);
   U9 : BUF_X1 port map( A => n152, Z => n94_port);
   U10 : BUF_X1 port map( A => n154, Z => n100_port);
   U11 : OAI21_X1 port map( B1 => n117, B2 => n120, A => n119, ZN => n154);
   U12 : AND3_X1 port map( A1 => n119, A2 => n118, A3 => n117, ZN => n153);
   U13 : AND2_X1 port map( A1 => n120, A2 => n119, ZN => n152);
   U14 : INV_X1 port map( A => n118, ZN => n120);
   U15 : NOR3_X1 port map( A1 => n109_port, A2 => n108_port, A3 => n107_port, 
                           ZN => n110_port);
   U16 : NAND4_X1 port map( A1 => n116, A2 => n115, A3 => n114, A4 => n113, ZN 
                           => n119);
   U17 : INV_X1 port map( A => addr_c(4), ZN => n115);
   U18 : NOR2_X1 port map( A1 => addr_c(1), A2 => addr_c(0), ZN => n113);
   U19 : NAND4_X1 port map( A1 => n112_port, A2 => valid_f, A3 => n111_port, A4
                           => n110_port, ZN => n118);
   U20 : XNOR2_X1 port map( A => addr_c(1), B => addr_f(1), ZN => n112_port);
   U21 : XNOR2_X1 port map( A => addr_c(0), B => addr_f(0), ZN => n111_port);
   U22 : INV_X1 port map( A => addr_c(2), ZN => n114);
   U23 : AND4_X1 port map( A1 => n106_port, A2 => valid_ff, A3 => n105_port, A4
                           => n104_port, ZN => n117);
   U24 : NOR3_X1 port map( A1 => n103_port, A2 => n102_port, A3 => n101_port, 
                           ZN => n104_port);
   U25 : INV_X1 port map( A => addr_c(3), ZN => n116);
   U26 : INV_X1 port map( A => n122, ZN => N101);
   U27 : AOI222_X1 port map( A1 => reg_c(22), A2 => n98_port, B1 => reg_ff(22),
                           B2 => n97_port, C1 => reg_f(22), C2 => n94_port, ZN 
                           => n122);
   U28 : INV_X1 port map( A => n123, ZN => N102);
   U29 : AOI222_X1 port map( A1 => reg_c(23), A2 => n98_port, B1 => reg_ff(23),
                           B2 => n97_port, C1 => reg_f(23), C2 => n94_port, ZN 
                           => n123);
   U30 : INV_X1 port map( A => n124, ZN => N103);
   U31 : AOI222_X1 port map( A1 => reg_c(24), A2 => n98_port, B1 => reg_ff(24),
                           B2 => n97_port, C1 => reg_f(24), C2 => n94_port, ZN 
                           => n124);
   U32 : INV_X1 port map( A => n125, ZN => N104);
   U33 : AOI222_X1 port map( A1 => reg_c(25), A2 => n98_port, B1 => reg_ff(25),
                           B2 => n97_port, C1 => reg_f(25), C2 => n94_port, ZN 
                           => n125);
   U34 : INV_X1 port map( A => n126, ZN => N105);
   U35 : AOI222_X1 port map( A1 => reg_c(26), A2 => n98_port, B1 => reg_ff(26),
                           B2 => n97_port, C1 => reg_f(26), C2 => n94_port, ZN 
                           => n126);
   U36 : INV_X1 port map( A => n127, ZN => N106);
   U37 : AOI222_X1 port map( A1 => reg_c(27), A2 => n98_port, B1 => reg_ff(27),
                           B2 => n97_port, C1 => reg_f(27), C2 => n94_port, ZN 
                           => n127);
   U38 : INV_X1 port map( A => n128, ZN => N107);
   U39 : AOI222_X1 port map( A1 => reg_c(28), A2 => n98_port, B1 => reg_ff(28),
                           B2 => n97_port, C1 => reg_f(28), C2 => n94_port, ZN 
                           => n128);
   U40 : INV_X1 port map( A => n129, ZN => N108);
   U41 : AOI222_X1 port map( A1 => reg_c(29), A2 => n98_port, B1 => reg_ff(29),
                           B2 => n97_port, C1 => reg_f(29), C2 => n94_port, ZN 
                           => n129);
   U42 : INV_X1 port map( A => n132, ZN => N79);
   U43 : AOI222_X1 port map( A1 => reg_c(0), A2 => n98_port, B1 => reg_ff(0), 
                           B2 => n96_port, C1 => reg_f(0), C2 => n93_port, ZN 
                           => n132);
   U44 : INV_X1 port map( A => n133, ZN => N80);
   U45 : AOI222_X1 port map( A1 => reg_c(1), A2 => n99_port, B1 => reg_ff(1), 
                           B2 => n96_port, C1 => reg_f(1), C2 => n93_port, ZN 
                           => n133);
   U46 : INV_X1 port map( A => n134, ZN => N81);
   U47 : AOI222_X1 port map( A1 => reg_c(2), A2 => n99_port, B1 => reg_ff(2), 
                           B2 => n96_port, C1 => reg_f(2), C2 => n93_port, ZN 
                           => n134);
   U48 : INV_X1 port map( A => n135, ZN => N82);
   U49 : AOI222_X1 port map( A1 => reg_c(3), A2 => n99_port, B1 => reg_ff(3), 
                           B2 => n96_port, C1 => reg_f(3), C2 => n93_port, ZN 
                           => n135);
   U50 : INV_X1 port map( A => n136, ZN => N83);
   U51 : AOI222_X1 port map( A1 => reg_c(4), A2 => n99_port, B1 => reg_ff(4), 
                           B2 => n96_port, C1 => reg_f(4), C2 => n93_port, ZN 
                           => n136);
   U52 : INV_X1 port map( A => n137, ZN => N84);
   U53 : AOI222_X1 port map( A1 => reg_c(5), A2 => n99_port, B1 => reg_ff(5), 
                           B2 => n96_port, C1 => reg_f(5), C2 => n93_port, ZN 
                           => n137);
   U54 : INV_X1 port map( A => n138, ZN => N85);
   U55 : AOI222_X1 port map( A1 => reg_c(6), A2 => n99_port, B1 => reg_ff(6), 
                           B2 => n96_port, C1 => reg_f(6), C2 => n93_port, ZN 
                           => n138);
   U56 : INV_X1 port map( A => n139, ZN => N86);
   U57 : AOI222_X1 port map( A1 => reg_c(7), A2 => n99_port, B1 => reg_ff(7), 
                           B2 => n96_port, C1 => reg_f(7), C2 => n93_port, ZN 
                           => n139);
   U58 : INV_X1 port map( A => n140, ZN => N87);
   U59 : AOI222_X1 port map( A1 => reg_c(8), A2 => n99_port, B1 => reg_ff(8), 
                           B2 => n96_port, C1 => reg_f(8), C2 => n93_port, ZN 
                           => n140);
   U60 : INV_X1 port map( A => n141, ZN => N88);
   U61 : AOI222_X1 port map( A1 => reg_c(9), A2 => n99_port, B1 => reg_ff(9), 
                           B2 => n95_port, C1 => reg_f(9), C2 => n92_port, ZN 
                           => n141);
   U62 : INV_X1 port map( A => n142, ZN => N89);
   U63 : AOI222_X1 port map( A1 => reg_c(10), A2 => n99_port, B1 => reg_ff(10),
                           B2 => n95_port, C1 => reg_f(10), C2 => n92_port, ZN 
                           => n142);
   U64 : INV_X1 port map( A => n143, ZN => N90);
   U65 : AOI222_X1 port map( A1 => reg_c(11), A2 => n99_port, B1 => reg_ff(11),
                           B2 => n95_port, C1 => reg_f(11), C2 => n92_port, ZN 
                           => n143);
   U66 : INV_X1 port map( A => n144, ZN => N91);
   U67 : AOI222_X1 port map( A1 => reg_c(12), A2 => n99_port, B1 => reg_ff(12),
                           B2 => n95_port, C1 => reg_f(12), C2 => n92_port, ZN 
                           => n144);
   U68 : INV_X1 port map( A => n145, ZN => N92);
   U69 : AOI222_X1 port map( A1 => reg_c(13), A2 => n100_port, B1 => reg_ff(13)
                           , B2 => n95_port, C1 => reg_f(13), C2 => n92_port, 
                           ZN => n145);
   U70 : INV_X1 port map( A => n146, ZN => N93);
   U71 : AOI222_X1 port map( A1 => reg_c(14), A2 => n100_port, B1 => reg_ff(14)
                           , B2 => n95_port, C1 => reg_f(14), C2 => n92_port, 
                           ZN => n146);
   U72 : INV_X1 port map( A => n147, ZN => N94);
   U73 : AOI222_X1 port map( A1 => reg_c(15), A2 => n100_port, B1 => reg_ff(15)
                           , B2 => n95_port, C1 => reg_f(15), C2 => n92_port, 
                           ZN => n147);
   U74 : INV_X1 port map( A => n148, ZN => N95);
   U75 : AOI222_X1 port map( A1 => reg_c(16), A2 => n100_port, B1 => reg_ff(16)
                           , B2 => n95_port, C1 => reg_f(16), C2 => n92_port, 
                           ZN => n148);
   U76 : INV_X1 port map( A => n149, ZN => N96);
   U77 : AOI222_X1 port map( A1 => reg_c(17), A2 => n100_port, B1 => reg_ff(17)
                           , B2 => n95_port, C1 => reg_f(17), C2 => n92_port, 
                           ZN => n149);
   U78 : INV_X1 port map( A => n150, ZN => N97);
   U79 : AOI222_X1 port map( A1 => reg_c(18), A2 => n100_port, B1 => reg_ff(18)
                           , B2 => n95_port, C1 => reg_f(18), C2 => n92_port, 
                           ZN => n150);
   U80 : INV_X1 port map( A => n151, ZN => N98);
   U81 : AOI222_X1 port map( A1 => reg_c(19), A2 => n100_port, B1 => reg_ff(19)
                           , B2 => n95_port, C1 => reg_f(19), C2 => n92_port, 
                           ZN => n151);
   U82 : INV_X1 port map( A => n155, ZN => N99);
   U91 : AOI222_X1 port map( A1 => reg_c(20), A2 => n100_port, B1 => reg_ff(20)
                           , B2 => n96_port, C1 => reg_f(20), C2 => n93_port, 
                           ZN => n155);
   U92 : INV_X1 port map( A => n121, ZN => N100);
   U93 : AOI222_X1 port map( A1 => reg_c(21), A2 => n98_port, B1 => reg_ff(21),
                           B2 => n95_port, C1 => reg_f(21), C2 => n92_port, ZN 
                           => n121);
   U94 : INV_X1 port map( A => n130, ZN => N109);
   U95 : AOI222_X1 port map( A1 => reg_c(30), A2 => n98_port, B1 => reg_ff(30),
                           B2 => n96_port, C1 => reg_f(30), C2 => n93_port, ZN 
                           => n130);
   U96 : INV_X1 port map( A => n131, ZN => N110);
   U97 : AOI222_X1 port map( A1 => reg_c(31), A2 => n98_port, B1 => reg_ff(31),
                           B2 => n96_port, C1 => reg_f(31), C2 => n93_port, ZN 
                           => n131);
   U98 : AND2_X1 port map( A1 => dirty_ff, A2 => n97_port, ZN => N111);
   U99 : AND2_X1 port map( A1 => dirty_f, A2 => n94_port, ZN => N112);

end SYN_fwd_mux_2_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_1 is

   port( reg_c, reg_f, reg_ff : in std_logic_vector (31 downto 0);  addr_c, 
         addr_f, addr_ff : in std_logic_vector (4 downto 0);  valid_f, valid_ff
         , dirty_f, dirty_ff, en : in std_logic;  output : out std_logic_vector
         (31 downto 0);  match_dirty_f, match_dirty_ff : out std_logic);

end FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_1;

architecture SYN_fwd_mux_2_arch of FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
      N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, 
      N106, N107, N108, N109, N110, N111, N112, n92_port, n93_port, n94_port, 
      n95_port, n96_port, n97_port, n98_port, n99_port, n100_port, n101_port, 
      n102_port, n103_port, n104_port, n105_port, n106_port, n107_port, 
      n108_port, n109_port, n110_port, n111_port, n112_port, n113, n114, n115, 
      n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
      n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155 : std_logic;

begin
   
   match_dirty_ff_reg : DLH_X1 port map( G => en, D => N111, Q => 
                           match_dirty_ff);
   output_reg_31_inst : DLH_X1 port map( G => en, D => N110, Q => output(31));
   output_reg_30_inst : DLH_X1 port map( G => en, D => N109, Q => output(30));
   output_reg_29_inst : DLH_X1 port map( G => en, D => N108, Q => output(29));
   output_reg_28_inst : DLH_X1 port map( G => en, D => N107, Q => output(28));
   output_reg_27_inst : DLH_X1 port map( G => en, D => N106, Q => output(27));
   output_reg_26_inst : DLH_X1 port map( G => en, D => N105, Q => output(26));
   output_reg_25_inst : DLH_X1 port map( G => en, D => N104, Q => output(25));
   output_reg_24_inst : DLH_X1 port map( G => en, D => N103, Q => output(24));
   output_reg_23_inst : DLH_X1 port map( G => en, D => N102, Q => output(23));
   output_reg_22_inst : DLH_X1 port map( G => en, D => N101, Q => output(22));
   output_reg_21_inst : DLH_X1 port map( G => en, D => N100, Q => output(21));
   output_reg_20_inst : DLH_X1 port map( G => en, D => N99, Q => output(20));
   output_reg_19_inst : DLH_X1 port map( G => en, D => N98, Q => output(19));
   output_reg_18_inst : DLH_X1 port map( G => en, D => N97, Q => output(18));
   output_reg_17_inst : DLH_X1 port map( G => en, D => N96, Q => output(17));
   output_reg_16_inst : DLH_X1 port map( G => en, D => N95, Q => output(16));
   output_reg_15_inst : DLH_X1 port map( G => en, D => N94, Q => output(15));
   output_reg_14_inst : DLH_X1 port map( G => en, D => N93, Q => output(14));
   output_reg_13_inst : DLH_X1 port map( G => en, D => N92, Q => output(13));
   output_reg_12_inst : DLH_X1 port map( G => en, D => N91, Q => output(12));
   output_reg_11_inst : DLH_X1 port map( G => en, D => N90, Q => output(11));
   output_reg_10_inst : DLH_X1 port map( G => en, D => N89, Q => output(10));
   output_reg_9_inst : DLH_X1 port map( G => en, D => N88, Q => output(9));
   output_reg_8_inst : DLH_X1 port map( G => en, D => N87, Q => output(8));
   output_reg_7_inst : DLH_X1 port map( G => en, D => N86, Q => output(7));
   output_reg_6_inst : DLH_X1 port map( G => en, D => N85, Q => output(6));
   output_reg_5_inst : DLH_X1 port map( G => en, D => N84, Q => output(5));
   output_reg_4_inst : DLH_X1 port map( G => en, D => N83, Q => output(4));
   output_reg_3_inst : DLH_X1 port map( G => en, D => N82, Q => output(3));
   output_reg_2_inst : DLH_X1 port map( G => en, D => N81, Q => output(2));
   output_reg_1_inst : DLH_X1 port map( G => en, D => N80, Q => output(1));
   output_reg_0_inst : DLH_X1 port map( G => en, D => N79, Q => output(0));
   match_dirty_f_reg : DLH_X1 port map( G => en, D => N112, Q => match_dirty_f)
                           ;
   U83 : XOR2_X1 port map( A => addr_f(3), B => addr_c(3), Z => n107_port);
   U84 : XOR2_X1 port map( A => addr_f(2), B => addr_c(2), Z => n108_port);
   U85 : XOR2_X1 port map( A => addr_f(4), B => addr_c(4), Z => n109_port);
   U86 : XOR2_X1 port map( A => addr_ff(4), B => addr_c(4), Z => n101_port);
   U87 : XOR2_X1 port map( A => addr_ff(0), B => addr_c(0), Z => n102_port);
   U88 : XOR2_X1 port map( A => addr_ff(1), B => addr_c(1), Z => n103_port);
   U89 : XOR2_X1 port map( A => n116, B => addr_ff(3), Z => n105_port);
   U90 : XOR2_X1 port map( A => n114, B => addr_ff(2), Z => n106_port);
   U2 : BUF_X1 port map( A => n153, Z => n95_port);
   U3 : BUF_X1 port map( A => n153, Z => n96_port);
   U4 : BUF_X1 port map( A => n152, Z => n92_port);
   U5 : BUF_X1 port map( A => n152, Z => n93_port);
   U6 : BUF_X1 port map( A => n153, Z => n97_port);
   U7 : BUF_X1 port map( A => n154, Z => n99_port);
   U8 : BUF_X1 port map( A => n154, Z => n98_port);
   U9 : BUF_X1 port map( A => n152, Z => n94_port);
   U10 : BUF_X1 port map( A => n154, Z => n100_port);
   U11 : OAI21_X1 port map( B1 => n117, B2 => n120, A => n119, ZN => n154);
   U12 : AND3_X1 port map( A1 => n119, A2 => n118, A3 => n117, ZN => n153);
   U13 : AND2_X1 port map( A1 => n120, A2 => n119, ZN => n152);
   U14 : INV_X1 port map( A => n118, ZN => n120);
   U15 : NAND4_X1 port map( A1 => n116, A2 => n115, A3 => n114, A4 => n113, ZN 
                           => n119);
   U16 : INV_X1 port map( A => addr_c(4), ZN => n115);
   U17 : NOR2_X1 port map( A1 => addr_c(1), A2 => addr_c(0), ZN => n113);
   U18 : NAND4_X1 port map( A1 => n112_port, A2 => valid_f, A3 => n111_port, A4
                           => n110_port, ZN => n118);
   U19 : XNOR2_X1 port map( A => addr_c(1), B => addr_f(1), ZN => n112_port);
   U20 : XNOR2_X1 port map( A => addr_c(0), B => addr_f(0), ZN => n111_port);
   U21 : NOR3_X1 port map( A1 => n109_port, A2 => n108_port, A3 => n107_port, 
                           ZN => n110_port);
   U22 : AND4_X1 port map( A1 => n106_port, A2 => valid_ff, A3 => n105_port, A4
                           => n104_port, ZN => n117);
   U23 : NOR3_X1 port map( A1 => n103_port, A2 => n102_port, A3 => n101_port, 
                           ZN => n104_port);
   U24 : INV_X1 port map( A => addr_c(2), ZN => n114);
   U25 : INV_X1 port map( A => addr_c(3), ZN => n116);
   U26 : INV_X1 port map( A => n122, ZN => N101);
   U27 : AOI222_X1 port map( A1 => reg_c(22), A2 => n98_port, B1 => reg_ff(22),
                           B2 => n97_port, C1 => reg_f(22), C2 => n94_port, ZN 
                           => n122);
   U28 : INV_X1 port map( A => n123, ZN => N102);
   U29 : AOI222_X1 port map( A1 => reg_c(23), A2 => n98_port, B1 => reg_ff(23),
                           B2 => n97_port, C1 => reg_f(23), C2 => n94_port, ZN 
                           => n123);
   U30 : INV_X1 port map( A => n124, ZN => N103);
   U31 : AOI222_X1 port map( A1 => reg_c(24), A2 => n98_port, B1 => reg_ff(24),
                           B2 => n97_port, C1 => reg_f(24), C2 => n94_port, ZN 
                           => n124);
   U32 : INV_X1 port map( A => n125, ZN => N104);
   U33 : AOI222_X1 port map( A1 => reg_c(25), A2 => n98_port, B1 => reg_ff(25),
                           B2 => n97_port, C1 => reg_f(25), C2 => n94_port, ZN 
                           => n125);
   U34 : INV_X1 port map( A => n126, ZN => N105);
   U35 : AOI222_X1 port map( A1 => reg_c(26), A2 => n98_port, B1 => reg_ff(26),
                           B2 => n97_port, C1 => reg_f(26), C2 => n94_port, ZN 
                           => n126);
   U36 : INV_X1 port map( A => n127, ZN => N106);
   U37 : AOI222_X1 port map( A1 => reg_c(27), A2 => n98_port, B1 => reg_ff(27),
                           B2 => n97_port, C1 => reg_f(27), C2 => n94_port, ZN 
                           => n127);
   U38 : INV_X1 port map( A => n128, ZN => N107);
   U39 : AOI222_X1 port map( A1 => reg_c(28), A2 => n98_port, B1 => reg_ff(28),
                           B2 => n97_port, C1 => reg_f(28), C2 => n94_port, ZN 
                           => n128);
   U40 : INV_X1 port map( A => n129, ZN => N108);
   U41 : AOI222_X1 port map( A1 => reg_c(29), A2 => n98_port, B1 => reg_ff(29),
                           B2 => n97_port, C1 => reg_f(29), C2 => n94_port, ZN 
                           => n129);
   U42 : INV_X1 port map( A => n132, ZN => N79);
   U43 : AOI222_X1 port map( A1 => reg_c(0), A2 => n98_port, B1 => reg_ff(0), 
                           B2 => n96_port, C1 => reg_f(0), C2 => n93_port, ZN 
                           => n132);
   U44 : INV_X1 port map( A => n133, ZN => N80);
   U45 : AOI222_X1 port map( A1 => reg_c(1), A2 => n99_port, B1 => reg_ff(1), 
                           B2 => n96_port, C1 => reg_f(1), C2 => n93_port, ZN 
                           => n133);
   U46 : INV_X1 port map( A => n134, ZN => N81);
   U47 : AOI222_X1 port map( A1 => reg_c(2), A2 => n99_port, B1 => reg_ff(2), 
                           B2 => n96_port, C1 => reg_f(2), C2 => n93_port, ZN 
                           => n134);
   U48 : INV_X1 port map( A => n135, ZN => N82);
   U49 : AOI222_X1 port map( A1 => reg_c(3), A2 => n99_port, B1 => reg_ff(3), 
                           B2 => n96_port, C1 => reg_f(3), C2 => n93_port, ZN 
                           => n135);
   U50 : INV_X1 port map( A => n136, ZN => N83);
   U51 : AOI222_X1 port map( A1 => reg_c(4), A2 => n99_port, B1 => reg_ff(4), 
                           B2 => n96_port, C1 => reg_f(4), C2 => n93_port, ZN 
                           => n136);
   U52 : INV_X1 port map( A => n137, ZN => N84);
   U53 : AOI222_X1 port map( A1 => reg_c(5), A2 => n99_port, B1 => reg_ff(5), 
                           B2 => n96_port, C1 => reg_f(5), C2 => n93_port, ZN 
                           => n137);
   U54 : INV_X1 port map( A => n138, ZN => N85);
   U55 : AOI222_X1 port map( A1 => reg_c(6), A2 => n99_port, B1 => reg_ff(6), 
                           B2 => n96_port, C1 => reg_f(6), C2 => n93_port, ZN 
                           => n138);
   U56 : INV_X1 port map( A => n139, ZN => N86);
   U57 : AOI222_X1 port map( A1 => reg_c(7), A2 => n99_port, B1 => reg_ff(7), 
                           B2 => n96_port, C1 => reg_f(7), C2 => n93_port, ZN 
                           => n139);
   U58 : INV_X1 port map( A => n140, ZN => N87);
   U59 : AOI222_X1 port map( A1 => reg_c(8), A2 => n99_port, B1 => reg_ff(8), 
                           B2 => n96_port, C1 => reg_f(8), C2 => n93_port, ZN 
                           => n140);
   U60 : INV_X1 port map( A => n141, ZN => N88);
   U61 : AOI222_X1 port map( A1 => reg_c(9), A2 => n99_port, B1 => reg_ff(9), 
                           B2 => n95_port, C1 => reg_f(9), C2 => n92_port, ZN 
                           => n141);
   U62 : INV_X1 port map( A => n142, ZN => N89);
   U63 : AOI222_X1 port map( A1 => reg_c(10), A2 => n99_port, B1 => reg_ff(10),
                           B2 => n95_port, C1 => reg_f(10), C2 => n92_port, ZN 
                           => n142);
   U64 : INV_X1 port map( A => n143, ZN => N90);
   U65 : AOI222_X1 port map( A1 => reg_c(11), A2 => n99_port, B1 => reg_ff(11),
                           B2 => n95_port, C1 => reg_f(11), C2 => n92_port, ZN 
                           => n143);
   U66 : INV_X1 port map( A => n144, ZN => N91);
   U67 : AOI222_X1 port map( A1 => reg_c(12), A2 => n99_port, B1 => reg_ff(12),
                           B2 => n95_port, C1 => reg_f(12), C2 => n92_port, ZN 
                           => n144);
   U68 : INV_X1 port map( A => n145, ZN => N92);
   U69 : AOI222_X1 port map( A1 => reg_c(13), A2 => n100_port, B1 => reg_ff(13)
                           , B2 => n95_port, C1 => reg_f(13), C2 => n92_port, 
                           ZN => n145);
   U70 : INV_X1 port map( A => n146, ZN => N93);
   U71 : AOI222_X1 port map( A1 => reg_c(14), A2 => n100_port, B1 => reg_ff(14)
                           , B2 => n95_port, C1 => reg_f(14), C2 => n92_port, 
                           ZN => n146);
   U72 : INV_X1 port map( A => n147, ZN => N94);
   U73 : AOI222_X1 port map( A1 => reg_c(15), A2 => n100_port, B1 => reg_ff(15)
                           , B2 => n95_port, C1 => reg_f(15), C2 => n92_port, 
                           ZN => n147);
   U74 : INV_X1 port map( A => n148, ZN => N95);
   U75 : AOI222_X1 port map( A1 => reg_c(16), A2 => n100_port, B1 => reg_ff(16)
                           , B2 => n95_port, C1 => reg_f(16), C2 => n92_port, 
                           ZN => n148);
   U76 : INV_X1 port map( A => n149, ZN => N96);
   U77 : AOI222_X1 port map( A1 => reg_c(17), A2 => n100_port, B1 => reg_ff(17)
                           , B2 => n95_port, C1 => reg_f(17), C2 => n92_port, 
                           ZN => n149);
   U78 : INV_X1 port map( A => n150, ZN => N97);
   U79 : AOI222_X1 port map( A1 => reg_c(18), A2 => n100_port, B1 => reg_ff(18)
                           , B2 => n95_port, C1 => reg_f(18), C2 => n92_port, 
                           ZN => n150);
   U80 : INV_X1 port map( A => n151, ZN => N98);
   U81 : AOI222_X1 port map( A1 => reg_c(19), A2 => n100_port, B1 => reg_ff(19)
                           , B2 => n95_port, C1 => reg_f(19), C2 => n92_port, 
                           ZN => n151);
   U82 : INV_X1 port map( A => n155, ZN => N99);
   U91 : AOI222_X1 port map( A1 => reg_c(20), A2 => n100_port, B1 => reg_ff(20)
                           , B2 => n96_port, C1 => reg_f(20), C2 => n93_port, 
                           ZN => n155);
   U92 : INV_X1 port map( A => n121, ZN => N100);
   U93 : AOI222_X1 port map( A1 => reg_c(21), A2 => n98_port, B1 => reg_ff(21),
                           B2 => n95_port, C1 => reg_f(21), C2 => n92_port, ZN 
                           => n121);
   U94 : INV_X1 port map( A => n130, ZN => N109);
   U95 : AOI222_X1 port map( A1 => reg_c(30), A2 => n98_port, B1 => reg_ff(30),
                           B2 => n96_port, C1 => reg_f(30), C2 => n93_port, ZN 
                           => n130);
   U96 : INV_X1 port map( A => n131, ZN => N110);
   U97 : AOI222_X1 port map( A1 => reg_c(31), A2 => n98_port, B1 => reg_ff(31),
                           B2 => n96_port, C1 => reg_f(31), C2 => n93_port, ZN 
                           => n131);
   U98 : AND2_X1 port map( A1 => dirty_ff, A2 => n97_port, ZN => N111);
   U99 : AND2_X1 port map( A1 => dirty_f, A2 => n94_port, ZN => N112);

end SYN_fwd_mux_2_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE32_11 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 0);
         dout : out std_logic_vector (31 downto 0));

end Reg_DATA_SIZE32_11;

architecture SYN_reg_arch of Reg_DATA_SIZE32_11 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, net108873, net108874, net108875, net108876, net108877, 
      net108878, net108879, net108880, net108881, net108882, net108883, 
      net108884, net108885, net108886, net108887, net108888, net108889, 
      net108890, net108891, net108892, net108893, net108894, net108895, 
      net108896, net108897, net108898, net108899, net108900, net108901, 
      net108902, net108903, net108904, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   dout_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => n67, Q => 
                           dout(31), QN => net108904);
   dout_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => n67, Q => 
                           dout(30), QN => net108903);
   dout_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => n67, Q => 
                           dout(29), QN => net108902);
   dout_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => n67, Q => 
                           dout(28), QN => net108901);
   dout_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => n67, Q => 
                           dout(27), QN => net108900);
   dout_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => n66, Q => 
                           dout(26), QN => net108899);
   dout_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => n66, Q => 
                           dout(25), QN => net108898);
   dout_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => n67, Q => 
                           dout(24), QN => net108897);
   dout_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => n66, Q => 
                           dout(23), QN => net108896);
   dout_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => n66, Q => 
                           dout(22), QN => net108895);
   dout_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => n66, Q => 
                           dout(21), QN => net108894);
   dout_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => n66, Q => 
                           dout(20), QN => net108893);
   dout_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => n65, Q => 
                           dout(19), QN => net108892);
   dout_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => n66, Q => 
                           dout(18), QN => net108891);
   dout_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => n65, Q => 
                           dout(17), QN => net108890);
   dout_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => n65, Q => 
                           dout(16), QN => net108889);
   dout_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => n66, Q => 
                           dout(15), QN => net108888);
   dout_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => n65, Q => 
                           dout(14), QN => net108887);
   dout_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => n65, Q => 
                           dout(13), QN => net108886);
   dout_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => n65, Q => 
                           dout(12), QN => net108885);
   dout_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => n65, Q => 
                           dout(11), QN => net108884);
   dout_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => n65, Q => 
                           dout(10), QN => net108883);
   dout_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => n67, Q => 
                           dout(9), QN => net108882);
   dout_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => n66, Q => 
                           dout(8), QN => net108881);
   dout_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => n66, Q => 
                           dout(7), QN => net108880);
   dout_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => n65, Q => 
                           dout(6), QN => net108879);
   dout_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => n66, Q => 
                           dout(5), QN => net108878);
   dout_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => n66, Q => 
                           dout(4), QN => net108877);
   dout_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => n65, Q => 
                           dout(3), QN => net108876);
   dout_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => n65, Q => 
                           dout(2), QN => net108875);
   dout_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => n65, Q => 
                           dout(1), QN => net108874);
   dout_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => n67, Q => 
                           dout(0), QN => net108873);
   U2 : BUF_X1 port map( A => rst, Z => n65);
   U3 : BUF_X1 port map( A => rst, Z => n66);
   U4 : BUF_X1 port map( A => rst, Z => n67);
   U5 : OAI21_X1 port map( B1 => net108873, B2 => en, A => n93, ZN => n32);
   U6 : NAND2_X1 port map( A1 => din(0), A2 => en, ZN => n93);
   U7 : OAI21_X1 port map( B1 => net108874, B2 => en, A => n92, ZN => n31);
   U8 : NAND2_X1 port map( A1 => din(1), A2 => en, ZN => n92);
   U9 : OAI21_X1 port map( B1 => net108875, B2 => en, A => n91, ZN => n30);
   U10 : NAND2_X1 port map( A1 => din(2), A2 => en, ZN => n91);
   U11 : OAI21_X1 port map( B1 => net108876, B2 => en, A => n89, ZN => n29);
   U12 : NAND2_X1 port map( A1 => din(3), A2 => en, ZN => n89);
   U13 : OAI21_X1 port map( B1 => net108877, B2 => en, A => n88, ZN => n28);
   U14 : NAND2_X1 port map( A1 => din(4), A2 => en, ZN => n88);
   U15 : OAI21_X1 port map( B1 => net108878, B2 => en, A => n87, ZN => n27);
   U16 : NAND2_X1 port map( A1 => din(5), A2 => en, ZN => n87);
   U17 : OAI21_X1 port map( B1 => net108879, B2 => en, A => n86, ZN => n26);
   U18 : NAND2_X1 port map( A1 => din(6), A2 => en, ZN => n86);
   U19 : OAI21_X1 port map( B1 => net108880, B2 => en, A => n85, ZN => n25);
   U20 : NAND2_X1 port map( A1 => din(7), A2 => en, ZN => n85);
   U21 : OAI21_X1 port map( B1 => net108881, B2 => en, A => n84, ZN => n24);
   U22 : NAND2_X1 port map( A1 => din(8), A2 => en, ZN => n84);
   U23 : OAI21_X1 port map( B1 => net108882, B2 => en, A => n83, ZN => n23);
   U24 : NAND2_X1 port map( A1 => din(9), A2 => en, ZN => n83);
   U25 : OAI21_X1 port map( B1 => net108883, B2 => en, A => n82, ZN => n22);
   U26 : NAND2_X1 port map( A1 => din(10), A2 => en, ZN => n82);
   U27 : OAI21_X1 port map( B1 => net108884, B2 => en, A => n81, ZN => n21);
   U28 : NAND2_X1 port map( A1 => din(11), A2 => en, ZN => n81);
   U29 : OAI21_X1 port map( B1 => net108885, B2 => en, A => n80, ZN => n20);
   U30 : NAND2_X1 port map( A1 => din(12), A2 => en, ZN => n80);
   U31 : OAI21_X1 port map( B1 => net108886, B2 => en, A => n78, ZN => n19);
   U32 : NAND2_X1 port map( A1 => din(13), A2 => en, ZN => n78);
   U33 : OAI21_X1 port map( B1 => net108887, B2 => en, A => n77, ZN => n18);
   U34 : NAND2_X1 port map( A1 => din(14), A2 => en, ZN => n77);
   U35 : OAI21_X1 port map( B1 => net108888, B2 => en, A => n76, ZN => n17);
   U36 : NAND2_X1 port map( A1 => din(15), A2 => en, ZN => n76);
   U37 : OAI21_X1 port map( B1 => net108889, B2 => en, A => n75, ZN => n16);
   U38 : NAND2_X1 port map( A1 => din(16), A2 => en, ZN => n75);
   U39 : OAI21_X1 port map( B1 => net108890, B2 => en, A => n74, ZN => n15);
   U40 : NAND2_X1 port map( A1 => din(17), A2 => en, ZN => n74);
   U41 : OAI21_X1 port map( B1 => net108891, B2 => en, A => n73, ZN => n14);
   U42 : NAND2_X1 port map( A1 => din(18), A2 => en, ZN => n73);
   U43 : OAI21_X1 port map( B1 => net108892, B2 => en, A => n72, ZN => n13);
   U44 : NAND2_X1 port map( A1 => din(19), A2 => en, ZN => n72);
   U45 : OAI21_X1 port map( B1 => net108893, B2 => en, A => n71, ZN => n12);
   U46 : NAND2_X1 port map( A1 => din(20), A2 => en, ZN => n71);
   U47 : OAI21_X1 port map( B1 => net108894, B2 => en, A => n70, ZN => n11);
   U48 : NAND2_X1 port map( A1 => din(21), A2 => en, ZN => n70);
   U49 : OAI21_X1 port map( B1 => net108895, B2 => en, A => n69, ZN => n10);
   U50 : NAND2_X1 port map( A1 => din(22), A2 => en, ZN => n69);
   U51 : OAI21_X1 port map( B1 => net108896, B2 => en, A => n99, ZN => n9);
   U52 : NAND2_X1 port map( A1 => en, A2 => din(23), ZN => n99);
   U53 : OAI21_X1 port map( B1 => net108897, B2 => en, A => n98, ZN => n8);
   U54 : NAND2_X1 port map( A1 => din(24), A2 => en, ZN => n98);
   U55 : OAI21_X1 port map( B1 => net108898, B2 => en, A => n97, ZN => n7);
   U56 : NAND2_X1 port map( A1 => din(25), A2 => en, ZN => n97);
   U57 : OAI21_X1 port map( B1 => net108899, B2 => en, A => n96, ZN => n6);
   U58 : NAND2_X1 port map( A1 => din(26), A2 => en, ZN => n96);
   U59 : OAI21_X1 port map( B1 => net108900, B2 => en, A => n95, ZN => n5);
   U60 : NAND2_X1 port map( A1 => din(27), A2 => en, ZN => n95);
   U61 : OAI21_X1 port map( B1 => net108901, B2 => en, A => n94, ZN => n4);
   U62 : NAND2_X1 port map( A1 => din(28), A2 => en, ZN => n94);
   U63 : OAI21_X1 port map( B1 => net108902, B2 => en, A => n90, ZN => n3);
   U64 : NAND2_X1 port map( A1 => din(29), A2 => en, ZN => n90);
   U65 : OAI21_X1 port map( B1 => net108903, B2 => en, A => n79, ZN => n2);
   U66 : NAND2_X1 port map( A1 => din(30), A2 => en, ZN => n79);
   U67 : OAI21_X1 port map( B1 => net108904, B2 => en, A => n68, ZN => n1);
   U68 : NAND2_X1 port map( A1 => din(31), A2 => en, ZN => n68);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE32_10 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 0);
         dout : out std_logic_vector (31 downto 0));

end Reg_DATA_SIZE32_10;

architecture SYN_reg_arch of Reg_DATA_SIZE32_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, net108873, net108874, net108875, net108876, net108877, 
      net108878, net108879, net108880, net108881, net108882, net108883, 
      net108884, net108885, net108886, net108887, net108888, net108889, 
      net108890, net108891, net108892, net108893, net108894, net108895, 
      net108896, net108897, net108898, net108899, net108900, net108901, 
      net108902, net108903, net108904, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   dout_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => n67, Q => 
                           dout(31), QN => net108904);
   dout_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => n67, Q => 
                           dout(30), QN => net108903);
   dout_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => n67, Q => 
                           dout(29), QN => net108902);
   dout_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => n67, Q => 
                           dout(28), QN => net108901);
   dout_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => n67, Q => 
                           dout(27), QN => net108900);
   dout_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => n66, Q => 
                           dout(26), QN => net108899);
   dout_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => n66, Q => 
                           dout(25), QN => net108898);
   dout_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => n67, Q => 
                           dout(24), QN => net108897);
   dout_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => n66, Q => 
                           dout(23), QN => net108896);
   dout_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => n66, Q => 
                           dout(22), QN => net108895);
   dout_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => n66, Q => 
                           dout(21), QN => net108894);
   dout_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => n66, Q => 
                           dout(20), QN => net108893);
   dout_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => n65, Q => 
                           dout(19), QN => net108892);
   dout_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => n66, Q => 
                           dout(18), QN => net108891);
   dout_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => n65, Q => 
                           dout(17), QN => net108890);
   dout_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => n65, Q => 
                           dout(16), QN => net108889);
   dout_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => n66, Q => 
                           dout(15), QN => net108888);
   dout_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => n65, Q => 
                           dout(14), QN => net108887);
   dout_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => n65, Q => 
                           dout(13), QN => net108886);
   dout_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => n65, Q => 
                           dout(12), QN => net108885);
   dout_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => n65, Q => 
                           dout(11), QN => net108884);
   dout_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => n65, Q => 
                           dout(10), QN => net108883);
   dout_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => n67, Q => 
                           dout(9), QN => net108882);
   dout_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => n66, Q => 
                           dout(8), QN => net108881);
   dout_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => n66, Q => 
                           dout(7), QN => net108880);
   dout_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => n65, Q => 
                           dout(6), QN => net108879);
   dout_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => n66, Q => 
                           dout(5), QN => net108878);
   dout_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => n66, Q => 
                           dout(4), QN => net108877);
   dout_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => n65, Q => 
                           dout(3), QN => net108876);
   dout_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => n65, Q => 
                           dout(2), QN => net108875);
   dout_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => n65, Q => 
                           dout(1), QN => net108874);
   dout_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => n67, Q => 
                           dout(0), QN => net108873);
   U2 : BUF_X1 port map( A => rst, Z => n65);
   U3 : BUF_X1 port map( A => rst, Z => n66);
   U4 : BUF_X1 port map( A => rst, Z => n67);
   U5 : OAI21_X1 port map( B1 => net108873, B2 => en, A => n93, ZN => n32);
   U6 : NAND2_X1 port map( A1 => din(0), A2 => en, ZN => n93);
   U7 : OAI21_X1 port map( B1 => net108874, B2 => en, A => n92, ZN => n31);
   U8 : NAND2_X1 port map( A1 => din(1), A2 => en, ZN => n92);
   U9 : OAI21_X1 port map( B1 => net108875, B2 => en, A => n91, ZN => n30);
   U10 : NAND2_X1 port map( A1 => din(2), A2 => en, ZN => n91);
   U11 : OAI21_X1 port map( B1 => net108876, B2 => en, A => n89, ZN => n29);
   U12 : NAND2_X1 port map( A1 => din(3), A2 => en, ZN => n89);
   U13 : OAI21_X1 port map( B1 => net108877, B2 => en, A => n88, ZN => n28);
   U14 : NAND2_X1 port map( A1 => din(4), A2 => en, ZN => n88);
   U15 : OAI21_X1 port map( B1 => net108878, B2 => en, A => n87, ZN => n27);
   U16 : NAND2_X1 port map( A1 => din(5), A2 => en, ZN => n87);
   U17 : OAI21_X1 port map( B1 => net108879, B2 => en, A => n86, ZN => n26);
   U18 : NAND2_X1 port map( A1 => din(6), A2 => en, ZN => n86);
   U19 : OAI21_X1 port map( B1 => net108880, B2 => en, A => n85, ZN => n25);
   U20 : NAND2_X1 port map( A1 => din(7), A2 => en, ZN => n85);
   U21 : OAI21_X1 port map( B1 => net108881, B2 => en, A => n84, ZN => n24);
   U22 : NAND2_X1 port map( A1 => din(8), A2 => en, ZN => n84);
   U23 : OAI21_X1 port map( B1 => net108882, B2 => en, A => n83, ZN => n23);
   U24 : NAND2_X1 port map( A1 => din(9), A2 => en, ZN => n83);
   U25 : OAI21_X1 port map( B1 => net108883, B2 => en, A => n82, ZN => n22);
   U26 : NAND2_X1 port map( A1 => din(10), A2 => en, ZN => n82);
   U27 : OAI21_X1 port map( B1 => net108884, B2 => en, A => n81, ZN => n21);
   U28 : NAND2_X1 port map( A1 => din(11), A2 => en, ZN => n81);
   U29 : OAI21_X1 port map( B1 => net108885, B2 => en, A => n80, ZN => n20);
   U30 : NAND2_X1 port map( A1 => din(12), A2 => en, ZN => n80);
   U31 : OAI21_X1 port map( B1 => net108886, B2 => en, A => n78, ZN => n19);
   U32 : NAND2_X1 port map( A1 => din(13), A2 => en, ZN => n78);
   U33 : OAI21_X1 port map( B1 => net108887, B2 => en, A => n77, ZN => n18);
   U34 : NAND2_X1 port map( A1 => din(14), A2 => en, ZN => n77);
   U35 : OAI21_X1 port map( B1 => net108888, B2 => en, A => n76, ZN => n17);
   U36 : NAND2_X1 port map( A1 => din(15), A2 => en, ZN => n76);
   U37 : OAI21_X1 port map( B1 => net108889, B2 => en, A => n75, ZN => n16);
   U38 : NAND2_X1 port map( A1 => din(16), A2 => en, ZN => n75);
   U39 : OAI21_X1 port map( B1 => net108890, B2 => en, A => n74, ZN => n15);
   U40 : NAND2_X1 port map( A1 => din(17), A2 => en, ZN => n74);
   U41 : OAI21_X1 port map( B1 => net108891, B2 => en, A => n73, ZN => n14);
   U42 : NAND2_X1 port map( A1 => din(18), A2 => en, ZN => n73);
   U43 : OAI21_X1 port map( B1 => net108892, B2 => en, A => n72, ZN => n13);
   U44 : NAND2_X1 port map( A1 => din(19), A2 => en, ZN => n72);
   U45 : OAI21_X1 port map( B1 => net108893, B2 => en, A => n71, ZN => n12);
   U46 : NAND2_X1 port map( A1 => din(20), A2 => en, ZN => n71);
   U47 : OAI21_X1 port map( B1 => net108894, B2 => en, A => n70, ZN => n11);
   U48 : NAND2_X1 port map( A1 => din(21), A2 => en, ZN => n70);
   U49 : OAI21_X1 port map( B1 => net108895, B2 => en, A => n69, ZN => n10);
   U50 : NAND2_X1 port map( A1 => din(22), A2 => en, ZN => n69);
   U51 : OAI21_X1 port map( B1 => net108896, B2 => en, A => n99, ZN => n9);
   U52 : NAND2_X1 port map( A1 => en, A2 => din(23), ZN => n99);
   U53 : OAI21_X1 port map( B1 => net108897, B2 => en, A => n98, ZN => n8);
   U54 : NAND2_X1 port map( A1 => din(24), A2 => en, ZN => n98);
   U55 : OAI21_X1 port map( B1 => net108898, B2 => en, A => n97, ZN => n7);
   U56 : NAND2_X1 port map( A1 => din(25), A2 => en, ZN => n97);
   U57 : OAI21_X1 port map( B1 => net108899, B2 => en, A => n96, ZN => n6);
   U58 : NAND2_X1 port map( A1 => din(26), A2 => en, ZN => n96);
   U59 : OAI21_X1 port map( B1 => net108900, B2 => en, A => n95, ZN => n5);
   U60 : NAND2_X1 port map( A1 => din(27), A2 => en, ZN => n95);
   U61 : OAI21_X1 port map( B1 => net108901, B2 => en, A => n94, ZN => n4);
   U62 : NAND2_X1 port map( A1 => din(28), A2 => en, ZN => n94);
   U63 : OAI21_X1 port map( B1 => net108902, B2 => en, A => n90, ZN => n3);
   U64 : NAND2_X1 port map( A1 => din(29), A2 => en, ZN => n90);
   U65 : OAI21_X1 port map( B1 => net108903, B2 => en, A => n79, ZN => n2);
   U66 : NAND2_X1 port map( A1 => din(30), A2 => en, ZN => n79);
   U67 : OAI21_X1 port map( B1 => net108904, B2 => en, A => n68, ZN => n1);
   U68 : NAND2_X1 port map( A1 => din(31), A2 => en, ZN => n68);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE32_9 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 0);
         dout : out std_logic_vector (31 downto 0));

end Reg_DATA_SIZE32_9;

architecture SYN_reg_arch of Reg_DATA_SIZE32_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component SDFFR_X1
      port( D, SI, SE, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, net108873, net108874, net108875, net108876, net108877, 
      net108878, net108879, net108880, net108881, net108882, net108883, 
      net108884, net108885, net108886, net108887, net108888, net108889, 
      net108890, net108891, net108892, net108893, net108894, net108895, 
      net108896, net108897, net108898, net108899, net108900, net108901, 
      net108902, net108903, net108904, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101 
      : std_logic;

begin
   
   dout_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => n69, Q => 
                           dout(31), QN => net108904);
   dout_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => n69, Q => 
                           dout(30), QN => net108903);
   dout_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => n69, Q => 
                           dout(29), QN => net108902);
   dout_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => n69, Q => 
                           dout(28), QN => net108901);
   dout_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => n69, Q => 
                           dout(27), QN => net108900);
   dout_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => n68, Q => 
                           dout(26), QN => net108899);
   dout_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => n68, Q => 
                           dout(25), QN => net108898);
   dout_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => n69, Q => 
                           dout(24), QN => net108897);
   dout_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => n68, Q => 
                           dout(23), QN => net108896);
   dout_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => n68, Q => 
                           dout(22), QN => net108895);
   dout_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => n68, Q => 
                           dout(21), QN => net108894);
   dout_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => n68, Q => 
                           dout(20), QN => net108893);
   dout_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => n67, Q => 
                           dout(19), QN => net108892);
   dout_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => n68, Q => 
                           dout(18), QN => net108891);
   dout_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => n67, Q => 
                           dout(17), QN => net108890);
   dout_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => n67, Q => 
                           dout(16), QN => net108889);
   dout_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => n68, Q => 
                           dout(15), QN => net108888);
   dout_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => n67, Q => 
                           dout(14), QN => net108887);
   dout_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => n67, Q => 
                           dout(13), QN => net108886);
   dout_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => n67, Q => 
                           dout(12), QN => net108885);
   dout_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => n67, Q => 
                           dout(11), QN => net108884);
   dout_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => n67, Q => 
                           dout(10), QN => net108883);
   dout_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => n69, Q => 
                           dout(9), QN => net108882);
   dout_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => n68, Q => 
                           dout(8), QN => net108881);
   dout_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => n68, Q => 
                           dout(7), QN => net108880);
   dout_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => n67, Q => 
                           dout(6), QN => net108879);
   dout_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => n68, Q => 
                           dout(5), QN => net108878);
   dout_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => n68, Q => 
                           dout(4), QN => net108877);
   dout_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => n67, Q => 
                           dout(3), QN => net108876);
   dout_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => n67, Q => 
                           dout(2), QN => net108875);
   dout_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => n67, Q => 
                           dout(1), QN => net108874);
   dout_reg_0_inst : SDFFR_X1 port map( D => n66, SI => n32, SE => n65, CK => 
                           clk, RN => n69, Q => dout(0), QN => net108873);
   n65 <= '1';
   n66 <= '0';
   U4 : BUF_X1 port map( A => rst, Z => n67);
   U5 : BUF_X1 port map( A => rst, Z => n68);
   U6 : BUF_X1 port map( A => rst, Z => n69);
   U7 : OAI21_X1 port map( B1 => net108889, B2 => en, A => n77, ZN => n16);
   U8 : NAND2_X1 port map( A1 => din(16), A2 => en, ZN => n77);
   U9 : OAI21_X1 port map( B1 => net108890, B2 => en, A => n76, ZN => n15);
   U10 : NAND2_X1 port map( A1 => din(17), A2 => en, ZN => n76);
   U11 : OAI21_X1 port map( B1 => net108891, B2 => en, A => n75, ZN => n14);
   U12 : NAND2_X1 port map( A1 => din(18), A2 => en, ZN => n75);
   U13 : OAI21_X1 port map( B1 => net108892, B2 => en, A => n74, ZN => n13);
   U14 : NAND2_X1 port map( A1 => din(19), A2 => en, ZN => n74);
   U15 : OAI21_X1 port map( B1 => net108894, B2 => en, A => n72, ZN => n11);
   U16 : NAND2_X1 port map( A1 => din(21), A2 => en, ZN => n72);
   U17 : OAI21_X1 port map( B1 => net108895, B2 => en, A => n71, ZN => n10);
   U18 : NAND2_X1 port map( A1 => din(22), A2 => en, ZN => n71);
   U19 : OAI21_X1 port map( B1 => net108896, B2 => en, A => n101, ZN => n9);
   U20 : NAND2_X1 port map( A1 => en, A2 => din(23), ZN => n101);
   U21 : OAI21_X1 port map( B1 => net108901, B2 => en, A => n96, ZN => n4);
   U22 : NAND2_X1 port map( A1 => din(28), A2 => en, ZN => n96);
   U23 : OAI21_X1 port map( B1 => net108904, B2 => en, A => n70, ZN => n1);
   U24 : NAND2_X1 port map( A1 => din(31), A2 => en, ZN => n70);
   U25 : OAI21_X1 port map( B1 => net108893, B2 => en, A => n73, ZN => n12);
   U26 : NAND2_X1 port map( A1 => din(20), A2 => en, ZN => n73);
   U27 : OAI21_X1 port map( B1 => net108897, B2 => en, A => n100, ZN => n8);
   U28 : NAND2_X1 port map( A1 => din(24), A2 => en, ZN => n100);
   U29 : OAI21_X1 port map( B1 => net108898, B2 => en, A => n99, ZN => n7);
   U30 : NAND2_X1 port map( A1 => din(25), A2 => en, ZN => n99);
   U31 : OAI21_X1 port map( B1 => net108899, B2 => en, A => n98, ZN => n6);
   U32 : NAND2_X1 port map( A1 => din(26), A2 => en, ZN => n98);
   U33 : OAI21_X1 port map( B1 => net108900, B2 => en, A => n97, ZN => n5);
   U34 : NAND2_X1 port map( A1 => din(27), A2 => en, ZN => n97);
   U35 : OAI21_X1 port map( B1 => net108902, B2 => en, A => n92, ZN => n3);
   U36 : NAND2_X1 port map( A1 => din(29), A2 => en, ZN => n92);
   U37 : OAI21_X1 port map( B1 => net108903, B2 => en, A => n81, ZN => n2);
   U38 : NAND2_X1 port map( A1 => din(30), A2 => en, ZN => n81);
   U39 : OAI21_X1 port map( B1 => net108879, B2 => en, A => n88, ZN => n26);
   U40 : NAND2_X1 port map( A1 => din(6), A2 => en, ZN => n88);
   U41 : OAI21_X1 port map( B1 => net108880, B2 => en, A => n87, ZN => n25);
   U42 : NAND2_X1 port map( A1 => din(7), A2 => en, ZN => n87);
   U43 : OAI21_X1 port map( B1 => net108883, B2 => en, A => n84, ZN => n22);
   U44 : NAND2_X1 port map( A1 => din(10), A2 => en, ZN => n84);
   U45 : OAI21_X1 port map( B1 => net108884, B2 => en, A => n83, ZN => n21);
   U46 : NAND2_X1 port map( A1 => din(11), A2 => en, ZN => n83);
   U47 : OAI21_X1 port map( B1 => net108885, B2 => en, A => n82, ZN => n20);
   U48 : NAND2_X1 port map( A1 => din(12), A2 => en, ZN => n82);
   U49 : OAI21_X1 port map( B1 => net108886, B2 => en, A => n80, ZN => n19);
   U50 : NAND2_X1 port map( A1 => din(13), A2 => en, ZN => n80);
   U51 : OAI21_X1 port map( B1 => net108887, B2 => en, A => n79, ZN => n18);
   U52 : NAND2_X1 port map( A1 => din(14), A2 => en, ZN => n79);
   U53 : OAI21_X1 port map( B1 => net108888, B2 => en, A => n78, ZN => n17);
   U54 : NAND2_X1 port map( A1 => din(15), A2 => en, ZN => n78);
   U55 : OAI21_X1 port map( B1 => net108877, B2 => en, A => n90, ZN => n28);
   U56 : NAND2_X1 port map( A1 => din(4), A2 => en, ZN => n90);
   U57 : OAI21_X1 port map( B1 => net108878, B2 => en, A => n89, ZN => n27);
   U58 : NAND2_X1 port map( A1 => din(5), A2 => en, ZN => n89);
   U59 : OAI21_X1 port map( B1 => net108881, B2 => en, A => n86, ZN => n24);
   U60 : NAND2_X1 port map( A1 => din(8), A2 => en, ZN => n86);
   U61 : OAI21_X1 port map( B1 => net108882, B2 => en, A => n85, ZN => n23);
   U62 : NAND2_X1 port map( A1 => din(9), A2 => en, ZN => n85);
   U63 : OAI21_X1 port map( B1 => net108874, B2 => en, A => n94, ZN => n31);
   U64 : NAND2_X1 port map( A1 => din(1), A2 => en, ZN => n94);
   U65 : OAI21_X1 port map( B1 => net108876, B2 => en, A => n91, ZN => n29);
   U66 : NAND2_X1 port map( A1 => din(3), A2 => en, ZN => n91);
   U67 : OAI21_X1 port map( B1 => net108875, B2 => en, A => n93, ZN => n30);
   U68 : NAND2_X1 port map( A1 => din(2), A2 => en, ZN => n93);
   U69 : OAI21_X1 port map( B1 => net108873, B2 => en, A => n95, ZN => n32);
   U70 : NAND2_X1 port map( A1 => din(0), A2 => en, ZN => n95);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE32_8 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 0);
         dout : out std_logic_vector (31 downto 0));

end Reg_DATA_SIZE32_8;

architecture SYN_reg_arch of Reg_DATA_SIZE32_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, net108873, net108874, net108875, net108876, net108877, 
      net108878, net108879, net108880, net108881, net108882, net108883, 
      net108884, net108885, net108886, net108887, net108888, net108889, 
      net108890, net108891, net108892, net108893, net108894, net108895, 
      net108896, net108897, net108898, net108899, net108900, net108901, 
      net108902, net108903, net108904, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   dout_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => n67, Q => 
                           dout(31), QN => net108904);
   dout_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => n67, Q => 
                           dout(30), QN => net108903);
   dout_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => n67, Q => 
                           dout(29), QN => net108902);
   dout_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => n67, Q => 
                           dout(28), QN => net108901);
   dout_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => n67, Q => 
                           dout(27), QN => net108900);
   dout_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => n66, Q => 
                           dout(26), QN => net108899);
   dout_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => n66, Q => 
                           dout(25), QN => net108898);
   dout_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => n67, Q => 
                           dout(24), QN => net108897);
   dout_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => n66, Q => 
                           dout(23), QN => net108896);
   dout_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => n66, Q => 
                           dout(22), QN => net108895);
   dout_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => n66, Q => 
                           dout(21), QN => net108894);
   dout_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => n66, Q => 
                           dout(20), QN => net108893);
   dout_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => n65, Q => 
                           dout(19), QN => net108892);
   dout_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => n66, Q => 
                           dout(18), QN => net108891);
   dout_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => n65, Q => 
                           dout(17), QN => net108890);
   dout_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => n65, Q => 
                           dout(16), QN => net108889);
   dout_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => n66, Q => 
                           dout(15), QN => net108888);
   dout_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => n65, Q => 
                           dout(14), QN => net108887);
   dout_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => n65, Q => 
                           dout(13), QN => net108886);
   dout_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => n65, Q => 
                           dout(12), QN => net108885);
   dout_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => n65, Q => 
                           dout(11), QN => net108884);
   dout_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => n65, Q => 
                           dout(10), QN => net108883);
   dout_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => n67, Q => 
                           dout(9), QN => net108882);
   dout_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => n66, Q => 
                           dout(8), QN => net108881);
   dout_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => n66, Q => 
                           dout(7), QN => net108880);
   dout_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => n65, Q => 
                           dout(6), QN => net108879);
   dout_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => n66, Q => 
                           dout(5), QN => net108878);
   dout_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => n66, Q => 
                           dout(4), QN => net108877);
   dout_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => n65, Q => 
                           dout(3), QN => net108876);
   dout_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => n65, Q => 
                           dout(2), QN => net108875);
   dout_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => n65, Q => 
                           dout(1), QN => net108874);
   dout_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => n67, Q => 
                           dout(0), QN => net108873);
   U2 : BUF_X1 port map( A => rst, Z => n65);
   U3 : BUF_X1 port map( A => rst, Z => n66);
   U4 : BUF_X1 port map( A => rst, Z => n67);
   U5 : OAI21_X1 port map( B1 => net108902, B2 => en, A => n90, ZN => n3);
   U6 : NAND2_X1 port map( A1 => din(29), A2 => en, ZN => n90);
   U7 : OAI21_X1 port map( B1 => net108903, B2 => en, A => n79, ZN => n2);
   U8 : NAND2_X1 port map( A1 => din(30), A2 => en, ZN => n79);
   U9 : OAI21_X1 port map( B1 => net108901, B2 => en, A => n94, ZN => n4);
   U10 : NAND2_X1 port map( A1 => din(28), A2 => en, ZN => n94);
   U11 : OAI21_X1 port map( B1 => net108897, B2 => en, A => n98, ZN => n8);
   U12 : NAND2_X1 port map( A1 => din(24), A2 => en, ZN => n98);
   U13 : OAI21_X1 port map( B1 => net108898, B2 => en, A => n97, ZN => n7);
   U14 : NAND2_X1 port map( A1 => din(25), A2 => en, ZN => n97);
   U15 : OAI21_X1 port map( B1 => net108899, B2 => en, A => n96, ZN => n6);
   U16 : NAND2_X1 port map( A1 => din(26), A2 => en, ZN => n96);
   U17 : OAI21_X1 port map( B1 => net108900, B2 => en, A => n95, ZN => n5);
   U18 : NAND2_X1 port map( A1 => din(27), A2 => en, ZN => n95);
   U19 : OAI21_X1 port map( B1 => net108873, B2 => en, A => n93, ZN => n32);
   U20 : NAND2_X1 port map( A1 => din(0), A2 => en, ZN => n93);
   U21 : OAI21_X1 port map( B1 => net108874, B2 => en, A => n92, ZN => n31);
   U22 : NAND2_X1 port map( A1 => din(1), A2 => en, ZN => n92);
   U23 : OAI21_X1 port map( B1 => net108875, B2 => en, A => n91, ZN => n30);
   U24 : NAND2_X1 port map( A1 => din(2), A2 => en, ZN => n91);
   U25 : OAI21_X1 port map( B1 => net108876, B2 => en, A => n89, ZN => n29);
   U26 : NAND2_X1 port map( A1 => din(3), A2 => en, ZN => n89);
   U27 : OAI21_X1 port map( B1 => net108877, B2 => en, A => n88, ZN => n28);
   U28 : NAND2_X1 port map( A1 => din(4), A2 => en, ZN => n88);
   U29 : OAI21_X1 port map( B1 => net108879, B2 => en, A => n86, ZN => n26);
   U30 : NAND2_X1 port map( A1 => din(6), A2 => en, ZN => n86);
   U31 : OAI21_X1 port map( B1 => net108880, B2 => en, A => n85, ZN => n25);
   U32 : NAND2_X1 port map( A1 => din(7), A2 => en, ZN => n85);
   U33 : OAI21_X1 port map( B1 => net108881, B2 => en, A => n84, ZN => n24);
   U34 : NAND2_X1 port map( A1 => din(8), A2 => en, ZN => n84);
   U35 : OAI21_X1 port map( B1 => net108882, B2 => en, A => n83, ZN => n23);
   U36 : NAND2_X1 port map( A1 => din(9), A2 => en, ZN => n83);
   U37 : OAI21_X1 port map( B1 => net108883, B2 => en, A => n82, ZN => n22);
   U38 : NAND2_X1 port map( A1 => din(10), A2 => en, ZN => n82);
   U39 : OAI21_X1 port map( B1 => net108884, B2 => en, A => n81, ZN => n21);
   U40 : NAND2_X1 port map( A1 => din(11), A2 => en, ZN => n81);
   U41 : OAI21_X1 port map( B1 => net108885, B2 => en, A => n80, ZN => n20);
   U42 : NAND2_X1 port map( A1 => din(12), A2 => en, ZN => n80);
   U43 : OAI21_X1 port map( B1 => net108886, B2 => en, A => n78, ZN => n19);
   U44 : NAND2_X1 port map( A1 => din(13), A2 => en, ZN => n78);
   U45 : OAI21_X1 port map( B1 => net108887, B2 => en, A => n77, ZN => n18);
   U46 : NAND2_X1 port map( A1 => din(14), A2 => en, ZN => n77);
   U47 : OAI21_X1 port map( B1 => net108888, B2 => en, A => n76, ZN => n17);
   U48 : NAND2_X1 port map( A1 => din(15), A2 => en, ZN => n76);
   U49 : OAI21_X1 port map( B1 => net108889, B2 => en, A => n75, ZN => n16);
   U50 : NAND2_X1 port map( A1 => din(16), A2 => en, ZN => n75);
   U51 : OAI21_X1 port map( B1 => net108890, B2 => en, A => n74, ZN => n15);
   U52 : NAND2_X1 port map( A1 => din(17), A2 => en, ZN => n74);
   U53 : OAI21_X1 port map( B1 => net108891, B2 => en, A => n73, ZN => n14);
   U54 : NAND2_X1 port map( A1 => din(18), A2 => en, ZN => n73);
   U55 : OAI21_X1 port map( B1 => net108892, B2 => en, A => n72, ZN => n13);
   U56 : NAND2_X1 port map( A1 => din(19), A2 => en, ZN => n72);
   U57 : OAI21_X1 port map( B1 => net108893, B2 => en, A => n71, ZN => n12);
   U58 : NAND2_X1 port map( A1 => din(20), A2 => en, ZN => n71);
   U59 : OAI21_X1 port map( B1 => net108894, B2 => en, A => n70, ZN => n11);
   U60 : NAND2_X1 port map( A1 => din(21), A2 => en, ZN => n70);
   U61 : OAI21_X1 port map( B1 => net108895, B2 => en, A => n69, ZN => n10);
   U62 : NAND2_X1 port map( A1 => din(22), A2 => en, ZN => n69);
   U63 : OAI21_X1 port map( B1 => net108904, B2 => en, A => n68, ZN => n1);
   U64 : NAND2_X1 port map( A1 => din(31), A2 => en, ZN => n68);
   U65 : OAI21_X1 port map( B1 => net108896, B2 => en, A => n99, ZN => n9);
   U66 : NAND2_X1 port map( A1 => en, A2 => din(23), ZN => n99);
   U67 : OAI21_X1 port map( B1 => net108878, B2 => en, A => n87, ZN => n27);
   U68 : NAND2_X1 port map( A1 => din(5), A2 => en, ZN => n87);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE32_7 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 0);
         dout : out std_logic_vector (31 downto 0));

end Reg_DATA_SIZE32_7;

architecture SYN_reg_arch of Reg_DATA_SIZE32_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, net108873, net108874, net108875, net108876, net108877, 
      net108878, net108879, net108880, net108881, net108882, net108883, 
      net108884, net108885, net108886, net108887, net108888, net108889, 
      net108890, net108891, net108892, net108893, net108894, net108895, 
      net108896, net108897, net108898, net108899, net108900, net108901, 
      net108902, net108903, net108904, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104 : std_logic;

begin
   
   dout_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => n72, Q => 
                           dout(31), QN => net108904);
   dout_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => n72, Q => 
                           dout(30), QN => net108903);
   dout_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => n72, Q => 
                           dout(29), QN => net108902);
   dout_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => n72, Q => 
                           dout(28), QN => net108901);
   dout_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => n72, Q => 
                           dout(27), QN => net108900);
   dout_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => n71, Q => 
                           dout(26), QN => net108899);
   dout_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => n71, Q => 
                           dout(25), QN => net108898);
   dout_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => n72, Q => 
                           dout(24), QN => net108897);
   dout_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => n71, Q => 
                           dout(23), QN => net108896);
   dout_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => n71, Q => 
                           dout(22), QN => net108895);
   dout_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => n71, Q => 
                           dout(21), QN => net108894);
   dout_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => n71, Q => 
                           dout(20), QN => net108893);
   dout_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => n70, Q => 
                           dout(19), QN => net108892);
   dout_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => n71, Q => 
                           dout(18), QN => net108891);
   dout_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => n70, Q => 
                           dout(17), QN => net108890);
   dout_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => n70, Q => 
                           dout(16), QN => net108889);
   dout_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => n71, Q => 
                           dout(15), QN => net108888);
   dout_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => n70, Q => 
                           dout(14), QN => net108887);
   dout_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => n70, Q => 
                           dout(13), QN => net108886);
   dout_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => n70, Q => 
                           dout(12), QN => net108885);
   dout_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => n70, Q => 
                           dout(11), QN => net108884);
   dout_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => n70, Q => 
                           dout(10), QN => net108883);
   dout_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => n72, Q => 
                           dout(9), QN => net108882);
   dout_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => n71, Q => 
                           dout(8), QN => net108881);
   dout_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => n71, Q => 
                           dout(7), QN => net108880);
   dout_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => n70, Q => 
                           dout(6), QN => net108879);
   dout_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => n71, Q => 
                           dout(5), QN => net108878);
   dout_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => n71, Q => 
                           dout(4), QN => net108877);
   dout_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => n70, Q => 
                           dout(3), QN => net108876);
   dout_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => n70, Q => 
                           dout(2), QN => net108875);
   dout_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => n70, Q => 
                           dout(1), QN => net108874);
   dout_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => n72, Q => 
                           dout(0), QN => net108873);
   U2 : OR2_X1 port map( A1 => net108873, A2 => en, ZN => n69);
   U3 : OR2_X1 port map( A1 => net108901, A2 => en, ZN => n68);
   U4 : OR2_X1 port map( A1 => net108902, A2 => en, ZN => n67);
   U5 : OR2_X1 port map( A1 => net108903, A2 => en, ZN => n66);
   U6 : OR2_X1 port map( A1 => net108904, A2 => en, ZN => n65);
   U7 : NAND2_X1 port map( A1 => n65, A2 => n73, ZN => n1);
   U8 : NAND2_X1 port map( A1 => n66, A2 => n84, ZN => n2);
   U9 : NAND2_X1 port map( A1 => n67, A2 => n95, ZN => n3);
   U10 : NAND2_X1 port map( A1 => n99, A2 => n68, ZN => n4);
   U11 : NAND2_X1 port map( A1 => n98, A2 => n69, ZN => n32);
   U12 : BUF_X1 port map( A => rst, Z => n70);
   U13 : BUF_X1 port map( A => rst, Z => n71);
   U14 : BUF_X1 port map( A => rst, Z => n72);
   U15 : NAND2_X1 port map( A1 => din(30), A2 => en, ZN => n84);
   U16 : NAND2_X1 port map( A1 => din(31), A2 => en, ZN => n73);
   U17 : OAI21_X1 port map( B1 => net108897, B2 => en, A => n103, ZN => n8);
   U18 : NAND2_X1 port map( A1 => din(24), A2 => en, ZN => n103);
   U19 : OAI21_X1 port map( B1 => net108891, B2 => en, A => n78, ZN => n14);
   U20 : NAND2_X1 port map( A1 => din(18), A2 => en, ZN => n78);
   U21 : OAI21_X1 port map( B1 => net108892, B2 => en, A => n77, ZN => n13);
   U22 : NAND2_X1 port map( A1 => din(19), A2 => en, ZN => n77);
   U23 : OAI21_X1 port map( B1 => net108896, B2 => en, A => n104, ZN => n9);
   U24 : NAND2_X1 port map( A1 => en, A2 => din(23), ZN => n104);
   U25 : OAI21_X1 port map( B1 => net108893, B2 => en, A => n76, ZN => n12);
   U26 : NAND2_X1 port map( A1 => din(20), A2 => en, ZN => n76);
   U27 : OAI21_X1 port map( B1 => net108894, B2 => en, A => n75, ZN => n11);
   U28 : NAND2_X1 port map( A1 => din(21), A2 => en, ZN => n75);
   U29 : OAI21_X1 port map( B1 => net108895, B2 => en, A => n74, ZN => n10);
   U30 : NAND2_X1 port map( A1 => din(22), A2 => en, ZN => n74);
   U31 : NAND2_X1 port map( A1 => din(28), A2 => en, ZN => n99);
   U32 : OAI21_X1 port map( B1 => net108900, B2 => en, A => n100, ZN => n5);
   U33 : NAND2_X1 port map( A1 => din(27), A2 => en, ZN => n100);
   U34 : OAI21_X1 port map( B1 => net108898, B2 => en, A => n102, ZN => n7);
   U35 : NAND2_X1 port map( A1 => din(25), A2 => en, ZN => n102);
   U36 : OAI21_X1 port map( B1 => net108899, B2 => en, A => n101, ZN => n6);
   U37 : NAND2_X1 port map( A1 => din(26), A2 => en, ZN => n101);
   U38 : OAI21_X1 port map( B1 => net108889, B2 => en, A => n80, ZN => n16);
   U39 : NAND2_X1 port map( A1 => din(16), A2 => en, ZN => n80);
   U40 : OAI21_X1 port map( B1 => net108890, B2 => en, A => n79, ZN => n15);
   U41 : NAND2_X1 port map( A1 => din(17), A2 => en, ZN => n79);
   U42 : OAI21_X1 port map( B1 => net108874, B2 => en, A => n97, ZN => n31);
   U43 : NAND2_X1 port map( A1 => din(1), A2 => en, ZN => n97);
   U44 : OAI21_X1 port map( B1 => net108875, B2 => en, A => n96, ZN => n30);
   U45 : NAND2_X1 port map( A1 => din(2), A2 => en, ZN => n96);
   U46 : OAI21_X1 port map( B1 => net108876, B2 => en, A => n94, ZN => n29);
   U47 : NAND2_X1 port map( A1 => din(3), A2 => en, ZN => n94);
   U48 : OAI21_X1 port map( B1 => net108877, B2 => en, A => n93, ZN => n28);
   U49 : NAND2_X1 port map( A1 => din(4), A2 => en, ZN => n93);
   U50 : OAI21_X1 port map( B1 => net108878, B2 => en, A => n92, ZN => n27);
   U51 : NAND2_X1 port map( A1 => din(5), A2 => en, ZN => n92);
   U52 : OAI21_X1 port map( B1 => net108879, B2 => en, A => n91, ZN => n26);
   U53 : NAND2_X1 port map( A1 => din(6), A2 => en, ZN => n91);
   U54 : OAI21_X1 port map( B1 => net108880, B2 => en, A => n90, ZN => n25);
   U55 : NAND2_X1 port map( A1 => din(7), A2 => en, ZN => n90);
   U56 : OAI21_X1 port map( B1 => net108881, B2 => en, A => n89, ZN => n24);
   U57 : NAND2_X1 port map( A1 => din(8), A2 => en, ZN => n89);
   U58 : OAI21_X1 port map( B1 => net108882, B2 => en, A => n88, ZN => n23);
   U59 : NAND2_X1 port map( A1 => din(9), A2 => en, ZN => n88);
   U60 : OAI21_X1 port map( B1 => net108883, B2 => en, A => n87, ZN => n22);
   U61 : NAND2_X1 port map( A1 => din(10), A2 => en, ZN => n87);
   U62 : OAI21_X1 port map( B1 => net108884, B2 => en, A => n86, ZN => n21);
   U63 : NAND2_X1 port map( A1 => din(11), A2 => en, ZN => n86);
   U64 : OAI21_X1 port map( B1 => net108885, B2 => en, A => n85, ZN => n20);
   U65 : NAND2_X1 port map( A1 => din(12), A2 => en, ZN => n85);
   U66 : OAI21_X1 port map( B1 => net108886, B2 => en, A => n83, ZN => n19);
   U67 : NAND2_X1 port map( A1 => din(13), A2 => en, ZN => n83);
   U68 : OAI21_X1 port map( B1 => net108887, B2 => en, A => n82, ZN => n18);
   U69 : NAND2_X1 port map( A1 => din(14), A2 => en, ZN => n82);
   U70 : OAI21_X1 port map( B1 => net108888, B2 => en, A => n81, ZN => n17);
   U71 : NAND2_X1 port map( A1 => din(15), A2 => en, ZN => n81);
   U72 : NAND2_X1 port map( A1 => din(29), A2 => en, ZN => n95);
   U73 : NAND2_X1 port map( A1 => din(0), A2 => en, ZN => n98);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE32_6 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 0);
         dout : out std_logic_vector (31 downto 0));

end Reg_DATA_SIZE32_6;

architecture SYN_reg_arch of Reg_DATA_SIZE32_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, net108873, net108874, net108875, net108876, net108877, 
      net108878, net108879, net108880, net108881, net108882, net108883, 
      net108884, net108885, net108886, net108887, net108888, net108889, 
      net108890, net108891, net108892, net108893, net108894, net108895, 
      net108896, net108897, net108898, net108899, net108900, net108901, 
      net108902, net108903, net108904, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   dout_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => n67, Q => 
                           dout(31), QN => net108904);
   dout_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => n67, Q => 
                           dout(30), QN => net108903);
   dout_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => n67, Q => 
                           dout(29), QN => net108902);
   dout_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => n67, Q => 
                           dout(28), QN => net108901);
   dout_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => n67, Q => 
                           dout(27), QN => net108900);
   dout_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => n66, Q => 
                           dout(26), QN => net108899);
   dout_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => n66, Q => 
                           dout(25), QN => net108898);
   dout_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => n67, Q => 
                           dout(24), QN => net108897);
   dout_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => n66, Q => 
                           dout(23), QN => net108896);
   dout_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => n66, Q => 
                           dout(22), QN => net108895);
   dout_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => n66, Q => 
                           dout(21), QN => net108894);
   dout_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => n66, Q => 
                           dout(20), QN => net108893);
   dout_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => n65, Q => 
                           dout(19), QN => net108892);
   dout_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => n66, Q => 
                           dout(18), QN => net108891);
   dout_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => n65, Q => 
                           dout(17), QN => net108890);
   dout_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => n65, Q => 
                           dout(16), QN => net108889);
   dout_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => n66, Q => 
                           dout(15), QN => net108888);
   dout_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => n65, Q => 
                           dout(14), QN => net108887);
   dout_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => n65, Q => 
                           dout(13), QN => net108886);
   dout_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => n65, Q => 
                           dout(12), QN => net108885);
   dout_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => n65, Q => 
                           dout(11), QN => net108884);
   dout_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => n65, Q => 
                           dout(10), QN => net108883);
   dout_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => n67, Q => 
                           dout(9), QN => net108882);
   dout_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => n66, Q => 
                           dout(8), QN => net108881);
   dout_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => n66, Q => 
                           dout(7), QN => net108880);
   dout_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => n65, Q => 
                           dout(6), QN => net108879);
   dout_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => n66, Q => 
                           dout(5), QN => net108878);
   dout_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => n66, Q => 
                           dout(4), QN => net108877);
   dout_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => n65, Q => 
                           dout(3), QN => net108876);
   dout_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => n65, Q => 
                           dout(2), QN => net108875);
   dout_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => n65, Q => 
                           dout(1), QN => net108874);
   dout_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => n67, Q => 
                           dout(0), QN => net108873);
   U2 : BUF_X1 port map( A => rst, Z => n65);
   U3 : BUF_X1 port map( A => rst, Z => n66);
   U4 : BUF_X1 port map( A => rst, Z => n67);
   U5 : OAI21_X1 port map( B1 => net108873, B2 => en, A => n93, ZN => n32);
   U6 : NAND2_X1 port map( A1 => din(0), A2 => en, ZN => n93);
   U7 : OAI21_X1 port map( B1 => net108874, B2 => en, A => n92, ZN => n31);
   U8 : NAND2_X1 port map( A1 => din(1), A2 => en, ZN => n92);
   U9 : OAI21_X1 port map( B1 => net108875, B2 => en, A => n91, ZN => n30);
   U10 : NAND2_X1 port map( A1 => din(2), A2 => en, ZN => n91);
   U11 : OAI21_X1 port map( B1 => net108876, B2 => en, A => n89, ZN => n29);
   U12 : NAND2_X1 port map( A1 => din(3), A2 => en, ZN => n89);
   U13 : OAI21_X1 port map( B1 => net108877, B2 => en, A => n88, ZN => n28);
   U14 : NAND2_X1 port map( A1 => din(4), A2 => en, ZN => n88);
   U15 : OAI21_X1 port map( B1 => net108878, B2 => en, A => n87, ZN => n27);
   U16 : NAND2_X1 port map( A1 => din(5), A2 => en, ZN => n87);
   U17 : OAI21_X1 port map( B1 => net108879, B2 => en, A => n86, ZN => n26);
   U18 : NAND2_X1 port map( A1 => din(6), A2 => en, ZN => n86);
   U19 : OAI21_X1 port map( B1 => net108880, B2 => en, A => n85, ZN => n25);
   U20 : NAND2_X1 port map( A1 => din(7), A2 => en, ZN => n85);
   U21 : OAI21_X1 port map( B1 => net108881, B2 => en, A => n84, ZN => n24);
   U22 : NAND2_X1 port map( A1 => din(8), A2 => en, ZN => n84);
   U23 : OAI21_X1 port map( B1 => net108882, B2 => en, A => n83, ZN => n23);
   U24 : NAND2_X1 port map( A1 => din(9), A2 => en, ZN => n83);
   U25 : OAI21_X1 port map( B1 => net108883, B2 => en, A => n82, ZN => n22);
   U26 : NAND2_X1 port map( A1 => din(10), A2 => en, ZN => n82);
   U27 : OAI21_X1 port map( B1 => net108884, B2 => en, A => n81, ZN => n21);
   U28 : NAND2_X1 port map( A1 => din(11), A2 => en, ZN => n81);
   U29 : OAI21_X1 port map( B1 => net108885, B2 => en, A => n80, ZN => n20);
   U30 : NAND2_X1 port map( A1 => din(12), A2 => en, ZN => n80);
   U31 : OAI21_X1 port map( B1 => net108886, B2 => en, A => n78, ZN => n19);
   U32 : NAND2_X1 port map( A1 => din(13), A2 => en, ZN => n78);
   U33 : OAI21_X1 port map( B1 => net108887, B2 => en, A => n77, ZN => n18);
   U34 : NAND2_X1 port map( A1 => din(14), A2 => en, ZN => n77);
   U35 : OAI21_X1 port map( B1 => net108888, B2 => en, A => n76, ZN => n17);
   U36 : NAND2_X1 port map( A1 => din(15), A2 => en, ZN => n76);
   U37 : OAI21_X1 port map( B1 => net108889, B2 => en, A => n75, ZN => n16);
   U38 : NAND2_X1 port map( A1 => din(16), A2 => en, ZN => n75);
   U39 : OAI21_X1 port map( B1 => net108890, B2 => en, A => n74, ZN => n15);
   U40 : NAND2_X1 port map( A1 => din(17), A2 => en, ZN => n74);
   U41 : OAI21_X1 port map( B1 => net108891, B2 => en, A => n73, ZN => n14);
   U42 : NAND2_X1 port map( A1 => din(18), A2 => en, ZN => n73);
   U43 : OAI21_X1 port map( B1 => net108892, B2 => en, A => n72, ZN => n13);
   U44 : NAND2_X1 port map( A1 => din(19), A2 => en, ZN => n72);
   U45 : OAI21_X1 port map( B1 => net108893, B2 => en, A => n71, ZN => n12);
   U46 : NAND2_X1 port map( A1 => din(20), A2 => en, ZN => n71);
   U47 : OAI21_X1 port map( B1 => net108894, B2 => en, A => n70, ZN => n11);
   U48 : NAND2_X1 port map( A1 => din(21), A2 => en, ZN => n70);
   U49 : OAI21_X1 port map( B1 => net108895, B2 => en, A => n69, ZN => n10);
   U50 : NAND2_X1 port map( A1 => din(22), A2 => en, ZN => n69);
   U51 : OAI21_X1 port map( B1 => net108896, B2 => en, A => n99, ZN => n9);
   U52 : NAND2_X1 port map( A1 => en, A2 => din(23), ZN => n99);
   U53 : OAI21_X1 port map( B1 => net108897, B2 => en, A => n98, ZN => n8);
   U54 : NAND2_X1 port map( A1 => din(24), A2 => en, ZN => n98);
   U55 : OAI21_X1 port map( B1 => net108898, B2 => en, A => n97, ZN => n7);
   U56 : NAND2_X1 port map( A1 => din(25), A2 => en, ZN => n97);
   U57 : OAI21_X1 port map( B1 => net108899, B2 => en, A => n96, ZN => n6);
   U58 : NAND2_X1 port map( A1 => din(26), A2 => en, ZN => n96);
   U59 : OAI21_X1 port map( B1 => net108900, B2 => en, A => n95, ZN => n5);
   U60 : NAND2_X1 port map( A1 => din(27), A2 => en, ZN => n95);
   U61 : OAI21_X1 port map( B1 => net108901, B2 => en, A => n94, ZN => n4);
   U62 : NAND2_X1 port map( A1 => din(28), A2 => en, ZN => n94);
   U63 : OAI21_X1 port map( B1 => net108902, B2 => en, A => n90, ZN => n3);
   U64 : NAND2_X1 port map( A1 => din(29), A2 => en, ZN => n90);
   U65 : OAI21_X1 port map( B1 => net108903, B2 => en, A => n79, ZN => n2);
   U66 : NAND2_X1 port map( A1 => din(30), A2 => en, ZN => n79);
   U67 : OAI21_X1 port map( B1 => net108904, B2 => en, A => n68, ZN => n1);
   U68 : NAND2_X1 port map( A1 => din(31), A2 => en, ZN => n68);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE32_5 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 0);
         dout : out std_logic_vector (31 downto 0));

end Reg_DATA_SIZE32_5;

architecture SYN_reg_arch of Reg_DATA_SIZE32_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, net108873, net108874, net108875, net108876, net108877, 
      net108878, net108879, net108880, net108881, net108882, net108883, 
      net108884, net108885, net108886, net108887, net108888, net108889, 
      net108890, net108891, net108892, net108893, net108894, net108895, 
      net108896, net108897, net108898, net108899, net108900, net108901, 
      net108902, net108903, net108904, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   dout_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => n67, Q => 
                           dout(31), QN => net108904);
   dout_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => n67, Q => 
                           dout(30), QN => net108903);
   dout_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => n67, Q => 
                           dout(29), QN => net108902);
   dout_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => n67, Q => 
                           dout(28), QN => net108901);
   dout_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => n67, Q => 
                           dout(27), QN => net108900);
   dout_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => n66, Q => 
                           dout(26), QN => net108899);
   dout_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => n66, Q => 
                           dout(25), QN => net108898);
   dout_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => n67, Q => 
                           dout(24), QN => net108897);
   dout_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => n66, Q => 
                           dout(23), QN => net108896);
   dout_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => n66, Q => 
                           dout(22), QN => net108895);
   dout_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => n66, Q => 
                           dout(21), QN => net108894);
   dout_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => n66, Q => 
                           dout(20), QN => net108893);
   dout_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => n65, Q => 
                           dout(19), QN => net108892);
   dout_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => n66, Q => 
                           dout(18), QN => net108891);
   dout_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => n65, Q => 
                           dout(17), QN => net108890);
   dout_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => n65, Q => 
                           dout(16), QN => net108889);
   dout_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => n66, Q => 
                           dout(15), QN => net108888);
   dout_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => n65, Q => 
                           dout(14), QN => net108887);
   dout_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => n65, Q => 
                           dout(13), QN => net108886);
   dout_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => n65, Q => 
                           dout(12), QN => net108885);
   dout_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => n65, Q => 
                           dout(11), QN => net108884);
   dout_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => n65, Q => 
                           dout(10), QN => net108883);
   dout_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => n67, Q => 
                           dout(9), QN => net108882);
   dout_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => n66, Q => 
                           dout(8), QN => net108881);
   dout_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => n66, Q => 
                           dout(7), QN => net108880);
   dout_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => n65, Q => 
                           dout(6), QN => net108879);
   dout_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => n66, Q => 
                           dout(5), QN => net108878);
   dout_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => n66, Q => 
                           dout(4), QN => net108877);
   dout_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => n65, Q => 
                           dout(3), QN => net108876);
   dout_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => n65, Q => 
                           dout(2), QN => net108875);
   dout_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => n65, Q => 
                           dout(1), QN => net108874);
   dout_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => n67, Q => 
                           dout(0), QN => net108873);
   U2 : BUF_X1 port map( A => rst, Z => n65);
   U3 : BUF_X1 port map( A => rst, Z => n66);
   U4 : BUF_X1 port map( A => rst, Z => n67);
   U5 : OAI21_X1 port map( B1 => net108892, B2 => en, A => n72, ZN => n13);
   U6 : NAND2_X1 port map( A1 => din(19), A2 => en, ZN => n72);
   U7 : OAI21_X1 port map( B1 => net108890, B2 => en, A => n74, ZN => n15);
   U8 : NAND2_X1 port map( A1 => din(17), A2 => en, ZN => n74);
   U9 : OAI21_X1 port map( B1 => net108891, B2 => en, A => n73, ZN => n14);
   U10 : NAND2_X1 port map( A1 => din(18), A2 => en, ZN => n73);
   U11 : OAI21_X1 port map( B1 => net108902, B2 => en, A => n90, ZN => n3);
   U12 : NAND2_X1 port map( A1 => din(29), A2 => en, ZN => n90);
   U13 : OAI21_X1 port map( B1 => net108903, B2 => en, A => n79, ZN => n2);
   U14 : NAND2_X1 port map( A1 => din(30), A2 => en, ZN => n79);
   U15 : OAI21_X1 port map( B1 => net108873, B2 => en, A => n93, ZN => n32);
   U16 : NAND2_X1 port map( A1 => din(0), A2 => en, ZN => n93);
   U17 : OAI21_X1 port map( B1 => net108874, B2 => en, A => n92, ZN => n31);
   U18 : NAND2_X1 port map( A1 => din(1), A2 => en, ZN => n92);
   U19 : OAI21_X1 port map( B1 => net108875, B2 => en, A => n91, ZN => n30);
   U20 : NAND2_X1 port map( A1 => din(2), A2 => en, ZN => n91);
   U21 : OAI21_X1 port map( B1 => net108876, B2 => en, A => n89, ZN => n29);
   U22 : NAND2_X1 port map( A1 => din(3), A2 => en, ZN => n89);
   U23 : OAI21_X1 port map( B1 => net108877, B2 => en, A => n88, ZN => n28);
   U24 : NAND2_X1 port map( A1 => din(4), A2 => en, ZN => n88);
   U25 : OAI21_X1 port map( B1 => net108878, B2 => en, A => n87, ZN => n27);
   U26 : NAND2_X1 port map( A1 => din(5), A2 => en, ZN => n87);
   U27 : OAI21_X1 port map( B1 => net108879, B2 => en, A => n86, ZN => n26);
   U28 : NAND2_X1 port map( A1 => din(6), A2 => en, ZN => n86);
   U29 : OAI21_X1 port map( B1 => net108880, B2 => en, A => n85, ZN => n25);
   U30 : NAND2_X1 port map( A1 => din(7), A2 => en, ZN => n85);
   U31 : OAI21_X1 port map( B1 => net108881, B2 => en, A => n84, ZN => n24);
   U32 : NAND2_X1 port map( A1 => din(8), A2 => en, ZN => n84);
   U33 : OAI21_X1 port map( B1 => net108882, B2 => en, A => n83, ZN => n23);
   U34 : NAND2_X1 port map( A1 => din(9), A2 => en, ZN => n83);
   U35 : OAI21_X1 port map( B1 => net108883, B2 => en, A => n82, ZN => n22);
   U36 : NAND2_X1 port map( A1 => din(10), A2 => en, ZN => n82);
   U37 : OAI21_X1 port map( B1 => net108884, B2 => en, A => n81, ZN => n21);
   U38 : NAND2_X1 port map( A1 => din(11), A2 => en, ZN => n81);
   U39 : OAI21_X1 port map( B1 => net108885, B2 => en, A => n80, ZN => n20);
   U40 : NAND2_X1 port map( A1 => din(12), A2 => en, ZN => n80);
   U41 : OAI21_X1 port map( B1 => net108886, B2 => en, A => n78, ZN => n19);
   U42 : NAND2_X1 port map( A1 => din(13), A2 => en, ZN => n78);
   U43 : OAI21_X1 port map( B1 => net108887, B2 => en, A => n77, ZN => n18);
   U44 : NAND2_X1 port map( A1 => din(14), A2 => en, ZN => n77);
   U45 : OAI21_X1 port map( B1 => net108888, B2 => en, A => n76, ZN => n17);
   U46 : NAND2_X1 port map( A1 => din(15), A2 => en, ZN => n76);
   U47 : OAI21_X1 port map( B1 => net108889, B2 => en, A => n75, ZN => n16);
   U48 : NAND2_X1 port map( A1 => din(16), A2 => en, ZN => n75);
   U49 : OAI21_X1 port map( B1 => net108893, B2 => en, A => n71, ZN => n12);
   U50 : NAND2_X1 port map( A1 => din(20), A2 => en, ZN => n71);
   U51 : OAI21_X1 port map( B1 => net108894, B2 => en, A => n70, ZN => n11);
   U52 : NAND2_X1 port map( A1 => din(21), A2 => en, ZN => n70);
   U53 : OAI21_X1 port map( B1 => net108895, B2 => en, A => n69, ZN => n10);
   U54 : NAND2_X1 port map( A1 => din(22), A2 => en, ZN => n69);
   U55 : OAI21_X1 port map( B1 => net108896, B2 => en, A => n99, ZN => n9);
   U56 : NAND2_X1 port map( A1 => en, A2 => din(23), ZN => n99);
   U57 : OAI21_X1 port map( B1 => net108897, B2 => en, A => n98, ZN => n8);
   U58 : NAND2_X1 port map( A1 => din(24), A2 => en, ZN => n98);
   U59 : OAI21_X1 port map( B1 => net108898, B2 => en, A => n97, ZN => n7);
   U60 : NAND2_X1 port map( A1 => din(25), A2 => en, ZN => n97);
   U61 : OAI21_X1 port map( B1 => net108899, B2 => en, A => n96, ZN => n6);
   U62 : NAND2_X1 port map( A1 => din(26), A2 => en, ZN => n96);
   U63 : OAI21_X1 port map( B1 => net108900, B2 => en, A => n95, ZN => n5);
   U64 : NAND2_X1 port map( A1 => din(27), A2 => en, ZN => n95);
   U65 : OAI21_X1 port map( B1 => net108901, B2 => en, A => n94, ZN => n4);
   U66 : NAND2_X1 port map( A1 => din(28), A2 => en, ZN => n94);
   U67 : OAI21_X1 port map( B1 => net108904, B2 => en, A => n68, ZN => n1);
   U68 : NAND2_X1 port map( A1 => din(31), A2 => en, ZN => n68);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE32_4 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 0);
         dout : out std_logic_vector (31 downto 0));

end Reg_DATA_SIZE32_4;

architecture SYN_reg_arch of Reg_DATA_SIZE32_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, net108873, net108874, net108875, net108876, net108877, 
      net108878, net108879, net108880, net108881, net108882, net108883, 
      net108884, net108885, net108886, net108887, net108888, net108889, 
      net108890, net108891, net108892, net108893, net108894, net108895, 
      net108896, net108897, net108898, net108899, net108900, net108901, 
      net108902, net108903, net108904, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   dout_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => n67, Q => 
                           dout(31), QN => net108904);
   dout_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => n67, Q => 
                           dout(30), QN => net108903);
   dout_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => n67, Q => 
                           dout(29), QN => net108902);
   dout_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => n67, Q => 
                           dout(28), QN => net108901);
   dout_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => n67, Q => 
                           dout(27), QN => net108900);
   dout_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => n66, Q => 
                           dout(26), QN => net108899);
   dout_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => n66, Q => 
                           dout(25), QN => net108898);
   dout_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => n67, Q => 
                           dout(24), QN => net108897);
   dout_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => n66, Q => 
                           dout(23), QN => net108896);
   dout_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => n66, Q => 
                           dout(22), QN => net108895);
   dout_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => n66, Q => 
                           dout(21), QN => net108894);
   dout_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => n66, Q => 
                           dout(20), QN => net108893);
   dout_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => n65, Q => 
                           dout(19), QN => net108892);
   dout_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => n66, Q => 
                           dout(18), QN => net108891);
   dout_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => n65, Q => 
                           dout(17), QN => net108890);
   dout_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => n65, Q => 
                           dout(16), QN => net108889);
   dout_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => n66, Q => 
                           dout(15), QN => net108888);
   dout_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => n65, Q => 
                           dout(14), QN => net108887);
   dout_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => n65, Q => 
                           dout(13), QN => net108886);
   dout_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => n65, Q => 
                           dout(12), QN => net108885);
   dout_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => n65, Q => 
                           dout(11), QN => net108884);
   dout_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => n65, Q => 
                           dout(10), QN => net108883);
   dout_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => n67, Q => 
                           dout(9), QN => net108882);
   dout_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => n66, Q => 
                           dout(8), QN => net108881);
   dout_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => n66, Q => 
                           dout(7), QN => net108880);
   dout_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => n65, Q => 
                           dout(6), QN => net108879);
   dout_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => n66, Q => 
                           dout(5), QN => net108878);
   dout_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => n66, Q => 
                           dout(4), QN => net108877);
   dout_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => n65, Q => 
                           dout(3), QN => net108876);
   dout_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => n65, Q => 
                           dout(2), QN => net108875);
   dout_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => n65, Q => 
                           dout(1), QN => net108874);
   dout_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => n67, Q => 
                           dout(0), QN => net108873);
   U2 : BUF_X1 port map( A => rst, Z => n65);
   U3 : BUF_X1 port map( A => rst, Z => n66);
   U4 : BUF_X1 port map( A => rst, Z => n67);
   U5 : OAI21_X1 port map( B1 => net108873, B2 => en, A => n93, ZN => n32);
   U6 : NAND2_X1 port map( A1 => din(0), A2 => en, ZN => n93);
   U7 : OAI21_X1 port map( B1 => net108874, B2 => en, A => n92, ZN => n31);
   U8 : NAND2_X1 port map( A1 => din(1), A2 => en, ZN => n92);
   U9 : OAI21_X1 port map( B1 => net108875, B2 => en, A => n91, ZN => n30);
   U10 : NAND2_X1 port map( A1 => din(2), A2 => en, ZN => n91);
   U11 : OAI21_X1 port map( B1 => net108876, B2 => en, A => n89, ZN => n29);
   U12 : NAND2_X1 port map( A1 => din(3), A2 => en, ZN => n89);
   U13 : OAI21_X1 port map( B1 => net108877, B2 => en, A => n88, ZN => n28);
   U14 : NAND2_X1 port map( A1 => din(4), A2 => en, ZN => n88);
   U15 : OAI21_X1 port map( B1 => net108878, B2 => en, A => n87, ZN => n27);
   U16 : NAND2_X1 port map( A1 => din(5), A2 => en, ZN => n87);
   U17 : OAI21_X1 port map( B1 => net108879, B2 => en, A => n86, ZN => n26);
   U18 : NAND2_X1 port map( A1 => din(6), A2 => en, ZN => n86);
   U19 : OAI21_X1 port map( B1 => net108880, B2 => en, A => n85, ZN => n25);
   U20 : NAND2_X1 port map( A1 => din(7), A2 => en, ZN => n85);
   U21 : OAI21_X1 port map( B1 => net108881, B2 => en, A => n84, ZN => n24);
   U22 : NAND2_X1 port map( A1 => din(8), A2 => en, ZN => n84);
   U23 : OAI21_X1 port map( B1 => net108882, B2 => en, A => n83, ZN => n23);
   U24 : NAND2_X1 port map( A1 => din(9), A2 => en, ZN => n83);
   U25 : OAI21_X1 port map( B1 => net108883, B2 => en, A => n82, ZN => n22);
   U26 : NAND2_X1 port map( A1 => din(10), A2 => en, ZN => n82);
   U27 : OAI21_X1 port map( B1 => net108884, B2 => en, A => n81, ZN => n21);
   U28 : NAND2_X1 port map( A1 => din(11), A2 => en, ZN => n81);
   U29 : OAI21_X1 port map( B1 => net108885, B2 => en, A => n80, ZN => n20);
   U30 : NAND2_X1 port map( A1 => din(12), A2 => en, ZN => n80);
   U31 : OAI21_X1 port map( B1 => net108886, B2 => en, A => n78, ZN => n19);
   U32 : NAND2_X1 port map( A1 => din(13), A2 => en, ZN => n78);
   U33 : OAI21_X1 port map( B1 => net108887, B2 => en, A => n77, ZN => n18);
   U34 : NAND2_X1 port map( A1 => din(14), A2 => en, ZN => n77);
   U35 : OAI21_X1 port map( B1 => net108888, B2 => en, A => n76, ZN => n17);
   U36 : NAND2_X1 port map( A1 => din(15), A2 => en, ZN => n76);
   U37 : OAI21_X1 port map( B1 => net108889, B2 => en, A => n75, ZN => n16);
   U38 : NAND2_X1 port map( A1 => din(16), A2 => en, ZN => n75);
   U39 : OAI21_X1 port map( B1 => net108890, B2 => en, A => n74, ZN => n15);
   U40 : NAND2_X1 port map( A1 => din(17), A2 => en, ZN => n74);
   U41 : OAI21_X1 port map( B1 => net108891, B2 => en, A => n73, ZN => n14);
   U42 : NAND2_X1 port map( A1 => din(18), A2 => en, ZN => n73);
   U43 : OAI21_X1 port map( B1 => net108892, B2 => en, A => n72, ZN => n13);
   U44 : NAND2_X1 port map( A1 => din(19), A2 => en, ZN => n72);
   U45 : OAI21_X1 port map( B1 => net108893, B2 => en, A => n71, ZN => n12);
   U46 : NAND2_X1 port map( A1 => din(20), A2 => en, ZN => n71);
   U47 : OAI21_X1 port map( B1 => net108894, B2 => en, A => n70, ZN => n11);
   U48 : NAND2_X1 port map( A1 => din(21), A2 => en, ZN => n70);
   U49 : OAI21_X1 port map( B1 => net108895, B2 => en, A => n69, ZN => n10);
   U50 : NAND2_X1 port map( A1 => din(22), A2 => en, ZN => n69);
   U51 : OAI21_X1 port map( B1 => net108896, B2 => en, A => n99, ZN => n9);
   U52 : NAND2_X1 port map( A1 => en, A2 => din(23), ZN => n99);
   U53 : OAI21_X1 port map( B1 => net108897, B2 => en, A => n98, ZN => n8);
   U54 : NAND2_X1 port map( A1 => din(24), A2 => en, ZN => n98);
   U55 : OAI21_X1 port map( B1 => net108898, B2 => en, A => n97, ZN => n7);
   U56 : NAND2_X1 port map( A1 => din(25), A2 => en, ZN => n97);
   U57 : OAI21_X1 port map( B1 => net108899, B2 => en, A => n96, ZN => n6);
   U58 : NAND2_X1 port map( A1 => din(26), A2 => en, ZN => n96);
   U59 : OAI21_X1 port map( B1 => net108900, B2 => en, A => n95, ZN => n5);
   U60 : NAND2_X1 port map( A1 => din(27), A2 => en, ZN => n95);
   U61 : OAI21_X1 port map( B1 => net108901, B2 => en, A => n94, ZN => n4);
   U62 : NAND2_X1 port map( A1 => din(28), A2 => en, ZN => n94);
   U63 : OAI21_X1 port map( B1 => net108902, B2 => en, A => n90, ZN => n3);
   U64 : NAND2_X1 port map( A1 => din(29), A2 => en, ZN => n90);
   U65 : OAI21_X1 port map( B1 => net108903, B2 => en, A => n79, ZN => n2);
   U66 : NAND2_X1 port map( A1 => din(30), A2 => en, ZN => n79);
   U67 : OAI21_X1 port map( B1 => net108904, B2 => en, A => n68, ZN => n1);
   U68 : NAND2_X1 port map( A1 => din(31), A2 => en, ZN => n68);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE32_2 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 0);
         dout : out std_logic_vector (31 downto 0));

end Reg_DATA_SIZE32_2;

architecture SYN_reg_arch of Reg_DATA_SIZE32_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, net108873, net108874, net108875, net108876, net108877, 
      net108878, net108879, net108880, net108881, net108882, net108883, 
      net108884, net108885, net108886, net108887, net108888, net108889, 
      net108890, net108891, net108892, net108893, net108894, net108895, 
      net108896, net108897, net108898, net108899, net108900, net108901, 
      net108902, net108903, net108904, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   dout_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => n67, Q => 
                           dout(31), QN => net108904);
   dout_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => n67, Q => 
                           dout(30), QN => net108903);
   dout_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => n67, Q => 
                           dout(29), QN => net108902);
   dout_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => n67, Q => 
                           dout(28), QN => net108901);
   dout_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => n67, Q => 
                           dout(27), QN => net108900);
   dout_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => n66, Q => 
                           dout(26), QN => net108899);
   dout_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => n66, Q => 
                           dout(25), QN => net108898);
   dout_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => n67, Q => 
                           dout(24), QN => net108897);
   dout_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => n66, Q => 
                           dout(23), QN => net108896);
   dout_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => n66, Q => 
                           dout(22), QN => net108895);
   dout_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => n66, Q => 
                           dout(21), QN => net108894);
   dout_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => n66, Q => 
                           dout(20), QN => net108893);
   dout_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => n65, Q => 
                           dout(19), QN => net108892);
   dout_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => n66, Q => 
                           dout(18), QN => net108891);
   dout_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => n65, Q => 
                           dout(17), QN => net108890);
   dout_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => n65, Q => 
                           dout(16), QN => net108889);
   dout_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => n66, Q => 
                           dout(15), QN => net108888);
   dout_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => n65, Q => 
                           dout(14), QN => net108887);
   dout_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => n65, Q => 
                           dout(13), QN => net108886);
   dout_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => n65, Q => 
                           dout(12), QN => net108885);
   dout_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => n65, Q => 
                           dout(11), QN => net108884);
   dout_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => n65, Q => 
                           dout(10), QN => net108883);
   dout_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => n67, Q => 
                           dout(9), QN => net108882);
   dout_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => n66, Q => 
                           dout(8), QN => net108881);
   dout_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => n66, Q => 
                           dout(7), QN => net108880);
   dout_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => n65, Q => 
                           dout(6), QN => net108879);
   dout_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => n66, Q => 
                           dout(5), QN => net108878);
   dout_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => n66, Q => 
                           dout(4), QN => net108877);
   dout_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => n65, Q => 
                           dout(3), QN => net108876);
   dout_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => n65, Q => 
                           dout(2), QN => net108875);
   dout_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => n65, Q => 
                           dout(1), QN => net108874);
   dout_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => n67, Q => 
                           dout(0), QN => net108873);
   U2 : BUF_X1 port map( A => rst, Z => n65);
   U3 : BUF_X1 port map( A => rst, Z => n66);
   U4 : BUF_X1 port map( A => rst, Z => n67);
   U5 : OAI21_X1 port map( B1 => net108873, B2 => en, A => n93, ZN => n32);
   U6 : NAND2_X1 port map( A1 => din(0), A2 => en, ZN => n93);
   U7 : OAI21_X1 port map( B1 => net108874, B2 => en, A => n92, ZN => n31);
   U8 : NAND2_X1 port map( A1 => din(1), A2 => en, ZN => n92);
   U9 : OAI21_X1 port map( B1 => net108875, B2 => en, A => n91, ZN => n30);
   U10 : NAND2_X1 port map( A1 => din(2), A2 => en, ZN => n91);
   U11 : OAI21_X1 port map( B1 => net108876, B2 => en, A => n89, ZN => n29);
   U12 : NAND2_X1 port map( A1 => din(3), A2 => en, ZN => n89);
   U13 : OAI21_X1 port map( B1 => net108877, B2 => en, A => n88, ZN => n28);
   U14 : NAND2_X1 port map( A1 => din(4), A2 => en, ZN => n88);
   U15 : OAI21_X1 port map( B1 => net108878, B2 => en, A => n87, ZN => n27);
   U16 : NAND2_X1 port map( A1 => din(5), A2 => en, ZN => n87);
   U17 : OAI21_X1 port map( B1 => net108879, B2 => en, A => n86, ZN => n26);
   U18 : NAND2_X1 port map( A1 => din(6), A2 => en, ZN => n86);
   U19 : OAI21_X1 port map( B1 => net108880, B2 => en, A => n85, ZN => n25);
   U20 : NAND2_X1 port map( A1 => din(7), A2 => en, ZN => n85);
   U21 : OAI21_X1 port map( B1 => net108881, B2 => en, A => n84, ZN => n24);
   U22 : NAND2_X1 port map( A1 => din(8), A2 => en, ZN => n84);
   U23 : OAI21_X1 port map( B1 => net108882, B2 => en, A => n83, ZN => n23);
   U24 : NAND2_X1 port map( A1 => din(9), A2 => en, ZN => n83);
   U25 : OAI21_X1 port map( B1 => net108883, B2 => en, A => n82, ZN => n22);
   U26 : NAND2_X1 port map( A1 => din(10), A2 => en, ZN => n82);
   U27 : OAI21_X1 port map( B1 => net108884, B2 => en, A => n81, ZN => n21);
   U28 : NAND2_X1 port map( A1 => din(11), A2 => en, ZN => n81);
   U29 : OAI21_X1 port map( B1 => net108885, B2 => en, A => n80, ZN => n20);
   U30 : NAND2_X1 port map( A1 => din(12), A2 => en, ZN => n80);
   U31 : OAI21_X1 port map( B1 => net108886, B2 => en, A => n78, ZN => n19);
   U32 : NAND2_X1 port map( A1 => din(13), A2 => en, ZN => n78);
   U33 : OAI21_X1 port map( B1 => net108887, B2 => en, A => n77, ZN => n18);
   U34 : NAND2_X1 port map( A1 => din(14), A2 => en, ZN => n77);
   U35 : OAI21_X1 port map( B1 => net108888, B2 => en, A => n76, ZN => n17);
   U36 : NAND2_X1 port map( A1 => din(15), A2 => en, ZN => n76);
   U37 : OAI21_X1 port map( B1 => net108889, B2 => en, A => n75, ZN => n16);
   U38 : NAND2_X1 port map( A1 => din(16), A2 => en, ZN => n75);
   U39 : OAI21_X1 port map( B1 => net108890, B2 => en, A => n74, ZN => n15);
   U40 : NAND2_X1 port map( A1 => din(17), A2 => en, ZN => n74);
   U41 : OAI21_X1 port map( B1 => net108891, B2 => en, A => n73, ZN => n14);
   U42 : NAND2_X1 port map( A1 => din(18), A2 => en, ZN => n73);
   U43 : OAI21_X1 port map( B1 => net108892, B2 => en, A => n72, ZN => n13);
   U44 : NAND2_X1 port map( A1 => din(19), A2 => en, ZN => n72);
   U45 : OAI21_X1 port map( B1 => net108893, B2 => en, A => n71, ZN => n12);
   U46 : NAND2_X1 port map( A1 => din(20), A2 => en, ZN => n71);
   U47 : OAI21_X1 port map( B1 => net108894, B2 => en, A => n70, ZN => n11);
   U48 : NAND2_X1 port map( A1 => din(21), A2 => en, ZN => n70);
   U49 : OAI21_X1 port map( B1 => net108895, B2 => en, A => n69, ZN => n10);
   U50 : NAND2_X1 port map( A1 => din(22), A2 => en, ZN => n69);
   U51 : OAI21_X1 port map( B1 => net108896, B2 => en, A => n99, ZN => n9);
   U52 : NAND2_X1 port map( A1 => en, A2 => din(23), ZN => n99);
   U53 : OAI21_X1 port map( B1 => net108897, B2 => en, A => n98, ZN => n8);
   U54 : NAND2_X1 port map( A1 => din(24), A2 => en, ZN => n98);
   U55 : OAI21_X1 port map( B1 => net108898, B2 => en, A => n97, ZN => n7);
   U56 : NAND2_X1 port map( A1 => din(25), A2 => en, ZN => n97);
   U57 : OAI21_X1 port map( B1 => net108899, B2 => en, A => n96, ZN => n6);
   U58 : NAND2_X1 port map( A1 => din(26), A2 => en, ZN => n96);
   U59 : OAI21_X1 port map( B1 => net108900, B2 => en, A => n95, ZN => n5);
   U60 : NAND2_X1 port map( A1 => din(27), A2 => en, ZN => n95);
   U61 : OAI21_X1 port map( B1 => net108901, B2 => en, A => n94, ZN => n4);
   U62 : NAND2_X1 port map( A1 => din(28), A2 => en, ZN => n94);
   U63 : OAI21_X1 port map( B1 => net108902, B2 => en, A => n90, ZN => n3);
   U64 : NAND2_X1 port map( A1 => din(29), A2 => en, ZN => n90);
   U65 : OAI21_X1 port map( B1 => net108903, B2 => en, A => n79, ZN => n2);
   U66 : NAND2_X1 port map( A1 => din(30), A2 => en, ZN => n79);
   U67 : OAI21_X1 port map( B1 => net108904, B2 => en, A => n68, ZN => n1);
   U68 : NAND2_X1 port map( A1 => din(31), A2 => en, ZN => n68);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE32_1 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 0);
         dout : out std_logic_vector (31 downto 0));

end Reg_DATA_SIZE32_1;

architecture SYN_reg_arch of Reg_DATA_SIZE32_1 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, net108873, net108874, net108875, net108876, net108877, 
      net108878, net108879, net108880, net108881, net108882, net108883, 
      net108884, net108885, net108886, net108887, net108888, net108889, 
      net108890, net108891, net108892, net108893, net108894, net108895, 
      net108896, net108897, net108898, net108899, net108900, net108901, 
      net108902, net108903, net108904, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109 : std_logic;

begin
   
   dout_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => n77, Q => 
                           dout(27), QN => net108900);
   dout_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => n76, Q => 
                           dout(26), QN => net108899);
   dout_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => n76, Q => 
                           dout(25), QN => net108898);
   dout_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => n77, Q => 
                           dout(24), QN => net108897);
   dout_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => n76, Q => 
                           dout(23), QN => net108896);
   dout_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => n76, Q => 
                           dout(22), QN => net108895);
   dout_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => n76, Q => 
                           dout(21), QN => net108894);
   dout_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => n76, Q => 
                           dout(20), QN => net108893);
   dout_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => n75, Q => 
                           dout(19), QN => net108892);
   dout_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => n76, Q => 
                           dout(18), QN => net108891);
   dout_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => n75, Q => 
                           dout(17), QN => net108890);
   dout_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => n75, Q => 
                           dout(16), QN => net108889);
   dout_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => n76, Q => 
                           dout(15), QN => net108888);
   dout_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => n75, Q => 
                           dout(13), QN => net108886);
   dout_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => n75, Q => 
                           dout(12), QN => net108885);
   dout_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => n75, Q => 
                           dout(11), QN => net108884);
   dout_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => n75, Q => 
                           dout(10), QN => net108883);
   dout_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => n76, Q => 
                           dout(8), QN => net108881);
   dout_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => n76, Q => 
                           dout(5), QN => net108878);
   dout_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => n76, Q => 
                           dout(4), QN => net108877);
   dout_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => n75, Q => 
                           dout(3), QN => net108876);
   dout_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => n75, Q => 
                           dout(2), QN => net108875);
   dout_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => n75, Q => 
                           dout(1), QN => net108874);
   dout_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => n77, Q => 
                           dout(28), QN => net108901);
   dout_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => n75, Q => 
                           dout(6), QN => net108879);
   dout_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => n76, Q => 
                           dout(7), QN => net108880);
   dout_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => n77, Q => 
                           dout(29), QN => net108902);
   dout_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => n77, Q => 
                           dout(30), QN => net108903);
   dout_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => n75, Q => 
                           dout(14), QN => net108887);
   dout_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => n77, Q => 
                           dout(0), QN => net108873);
   dout_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => n77, Q => 
                           dout(31), QN => net108904);
   dout_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => n77, Q => 
                           dout(9), QN => net108882);
   U2 : OR2_X1 port map( A1 => net108902, A2 => n72, ZN => n65);
   U3 : NAND2_X1 port map( A1 => n100, A2 => n65, ZN => n3);
   U4 : OR2_X1 port map( A1 => net108903, A2 => n73, ZN => n66);
   U5 : NAND2_X1 port map( A1 => n89, A2 => n66, ZN => n2);
   U6 : OR2_X1 port map( A1 => net108904, A2 => n72, ZN => n67);
   U7 : NAND2_X1 port map( A1 => n78, A2 => n67, ZN => n1);
   U8 : BUF_X1 port map( A => rst, Z => n75);
   U9 : BUF_X1 port map( A => rst, Z => n76);
   U10 : BUF_X1 port map( A => rst, Z => n77);
   U11 : BUF_X1 port map( A => en, Z => n69);
   U12 : BUF_X1 port map( A => en, Z => n73);
   U13 : BUF_X1 port map( A => en, Z => n70);
   U14 : BUF_X1 port map( A => en, Z => n72);
   U15 : OAI21_X1 port map( B1 => net108889, B2 => n73, A => n85, ZN => n16);
   U16 : NAND2_X1 port map( A1 => din(16), A2 => n69, ZN => n85);
   U17 : OAI21_X1 port map( B1 => net108890, B2 => n73, A => n84, ZN => n15);
   U18 : NAND2_X1 port map( A1 => din(17), A2 => n69, ZN => n84);
   U19 : OAI21_X1 port map( B1 => net108892, B2 => n73, A => n82, ZN => n13);
   U20 : NAND2_X1 port map( A1 => din(19), A2 => n69, ZN => n82);
   U21 : OAI21_X1 port map( B1 => net108897, B2 => n71, A => n108, ZN => n8);
   U22 : NAND2_X1 port map( A1 => din(24), A2 => n69, ZN => n108);
   U23 : OAI21_X1 port map( B1 => net108898, B2 => n71, A => n107, ZN => n7);
   U24 : NAND2_X1 port map( A1 => din(25), A2 => n69, ZN => n107);
   U25 : OAI21_X1 port map( B1 => net108900, B2 => n71, A => n105, ZN => n5);
   U26 : NAND2_X1 port map( A1 => din(27), A2 => n69, ZN => n105);
   U27 : OAI21_X1 port map( B1 => net108881, B2 => n72, A => n94, ZN => n24);
   U28 : NAND2_X1 port map( A1 => din(8), A2 => n71, ZN => n94);
   U29 : OAI21_X1 port map( B1 => net108882, B2 => n73, A => n93, ZN => n23);
   U30 : NAND2_X1 port map( A1 => din(9), A2 => n71, ZN => n93);
   U31 : OAI21_X1 port map( B1 => net108891, B2 => n73, A => n83, ZN => n14);
   U32 : NAND2_X1 port map( A1 => din(18), A2 => n69, ZN => n83);
   U33 : OAI21_X1 port map( B1 => net108883, B2 => n73, A => n92, ZN => n22);
   U34 : NAND2_X1 port map( A1 => din(10), A2 => n70, ZN => n92);
   U35 : OAI21_X1 port map( B1 => net108884, B2 => n73, A => n91, ZN => n21);
   U36 : NAND2_X1 port map( A1 => din(11), A2 => n70, ZN => n91);
   U37 : OAI21_X1 port map( B1 => net108885, B2 => n73, A => n90, ZN => n20);
   U38 : NAND2_X1 port map( A1 => din(12), A2 => n70, ZN => n90);
   U39 : OAI21_X1 port map( B1 => net108886, B2 => n73, A => n88, ZN => n19);
   U40 : NAND2_X1 port map( A1 => din(13), A2 => n70, ZN => n88);
   U41 : OAI21_X1 port map( B1 => net108887, B2 => n73, A => n87, ZN => n18);
   U42 : NAND2_X1 port map( A1 => din(14), A2 => n70, ZN => n87);
   U43 : OAI21_X1 port map( B1 => net108888, B2 => n73, A => n86, ZN => n17);
   U44 : NAND2_X1 port map( A1 => din(15), A2 => n70, ZN => n86);
   U45 : OAI21_X1 port map( B1 => net108893, B2 => n74, A => n81, ZN => n12);
   U46 : NAND2_X1 port map( A1 => din(20), A2 => n69, ZN => n81);
   U47 : OAI21_X1 port map( B1 => net108894, B2 => n74, A => n80, ZN => n11);
   U48 : NAND2_X1 port map( A1 => din(21), A2 => n69, ZN => n80);
   U49 : OAI21_X1 port map( B1 => net108895, B2 => n74, A => n79, ZN => n10);
   U50 : NAND2_X1 port map( A1 => din(22), A2 => n69, ZN => n79);
   U51 : OAI21_X1 port map( B1 => net108880, B2 => n72, A => n95, ZN => n25);
   U52 : NAND2_X1 port map( A1 => din(7), A2 => n71, ZN => n95);
   U53 : OAI21_X1 port map( B1 => net108899, B2 => n72, A => n106, ZN => n6);
   U54 : NAND2_X1 port map( A1 => din(26), A2 => n69, ZN => n106);
   U55 : OAI21_X1 port map( B1 => net108896, B2 => n72, A => n109, ZN => n9);
   U56 : NAND2_X1 port map( A1 => n74, A2 => din(23), ZN => n109);
   U57 : OAI21_X1 port map( B1 => net108874, B2 => n71, A => n102, ZN => n31);
   U58 : NAND2_X1 port map( A1 => din(1), A2 => n70, ZN => n102);
   U59 : OAI21_X1 port map( B1 => net108877, B2 => n72, A => n98, ZN => n28);
   U60 : NAND2_X1 port map( A1 => din(4), A2 => n71, ZN => n98);
   U61 : OAI21_X1 port map( B1 => net108878, B2 => n72, A => n97, ZN => n27);
   U62 : NAND2_X1 port map( A1 => din(5), A2 => n71, ZN => n97);
   U63 : OAI21_X1 port map( B1 => net108873, B2 => n72, A => n103, ZN => n32);
   U64 : NAND2_X1 port map( A1 => din(0), A2 => n70, ZN => n103);
   U65 : OAI21_X1 port map( B1 => net108879, B2 => n72, A => n96, ZN => n26);
   U66 : NAND2_X1 port map( A1 => din(6), A2 => n71, ZN => n96);
   U67 : OAI21_X1 port map( B1 => net108876, B2 => n72, A => n99, ZN => n29);
   U68 : NAND2_X1 port map( A1 => din(3), A2 => n70, ZN => n99);
   U69 : OAI21_X1 port map( B1 => net108875, B2 => n72, A => n101, ZN => n30);
   U70 : NAND2_X1 port map( A1 => din(2), A2 => n70, ZN => n101);
   U71 : OR2_X1 port map( A1 => net108901, A2 => n71, ZN => n68);
   U72 : NAND2_X1 port map( A1 => n104, A2 => n68, ZN => n4);
   U73 : BUF_X1 port map( A => en, Z => n71);
   U74 : NAND2_X1 port map( A1 => din(28), A2 => n70, ZN => n104);
   U75 : NAND2_X1 port map( A1 => din(30), A2 => n70, ZN => n89);
   U76 : NAND2_X1 port map( A1 => din(29), A2 => n71, ZN => n100);
   U77 : NAND2_X1 port map( A1 => din(31), A2 => n69, ZN => n78);
   U78 : CLKBUF_X1 port map( A => en, Z => n74);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE32_9 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0);  
         dout : out std_logic_vector (31 downto 0));

end Mux_DATA_SIZE32_9;

architecture SYN_mux_arch of Mux_DATA_SIZE32_9 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal net134080, net134078, net134076, net134074, net134072, net134070, 
      net134068, net134066, net139420, net139419, net153543, n1, n2, n4, n5, n6
      , n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n35, n36 : 
      std_logic;

begin
   
   syn103 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => 
                           dout(0));
   U1 : BUF_X2 port map( A => net139419, Z => net139420);
   U2 : INV_X1 port map( A => n2, ZN => n1);
   U3 : BUF_X1 port map( A => sel, Z => n2);
   U4 : CLKBUF_X1 port map( A => n2, Z => net134076);
   U5 : INV_X1 port map( A => n2, ZN => net139419);
   U6 : INV_X1 port map( A => n1, ZN => net153543);
   U7 : CLKBUF_X1 port map( A => net153543, Z => net134070);
   U8 : CLKBUF_X1 port map( A => net134072, Z => net134074);
   U9 : CLKBUF_X1 port map( A => net134078, Z => net134080);
   U10 : CLKBUF_X1 port map( A => net134070, Z => net134078);
   U11 : INV_X1 port map( A => n7, ZN => dout(11));
   U12 : INV_X1 port map( A => n15, ZN => dout(19));
   U13 : INV_X1 port map( A => n21, ZN => dout(24));
   U14 : INV_X1 port map( A => n17, ZN => dout(20));
   U15 : INV_X1 port map( A => n22, ZN => dout(25));
   U16 : INV_X1 port map( A => n23, ZN => dout(26));
   U17 : INV_X1 port map( A => n18, ZN => dout(21));
   U18 : INV_X1 port map( A => n19, ZN => dout(22));
   U19 : INV_X1 port map( A => n26, ZN => dout(2));
   U20 : INV_X1 port map( A => n20, ZN => dout(23));
   U21 : INV_X1 port map( A => n6, ZN => dout(10));
   U22 : INV_X1 port map( A => n11, ZN => dout(15));
   U23 : INV_X1 port map( A => n8, ZN => dout(12));
   U24 : INV_X1 port map( A => n28, ZN => dout(31));
   U25 : INV_X1 port map( A => n35, ZN => dout(8));
   U26 : INV_X1 port map( A => n12, ZN => dout(16));
   U27 : INV_X1 port map( A => n29, ZN => dout(3));
   U28 : INV_X1 port map( A => n30, ZN => dout(4));
   U29 : INV_X1 port map( A => n13, ZN => dout(17));
   U30 : INV_X1 port map( A => n36, ZN => dout(9));
   U31 : INV_X1 port map( A => n14, ZN => dout(18));
   U32 : INV_X1 port map( A => n33, ZN => dout(7));
   U33 : INV_X1 port map( A => n32, ZN => dout(6));
   U34 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => dout(29));
   U35 : CLKBUF_X1 port map( A => net153543, Z => net134068);
   U36 : INV_X1 port map( A => net134076, ZN => net134066);
   U37 : NAND2_X1 port map( A1 => din0(29), A2 => net134066, ZN => n4);
   U38 : NAND2_X1 port map( A1 => din1(29), A2 => net134072, ZN => n5);
   U39 : INV_X1 port map( A => n27, ZN => dout(30));
   U40 : INV_X1 port map( A => n9, ZN => dout(13));
   U41 : INV_X1 port map( A => n10, ZN => dout(14));
   U42 : INV_X1 port map( A => n24, ZN => dout(27));
   U43 : AOI22_X1 port map( A1 => din0(27), A2 => net139420, B1 => din1(27), B2
                           => net134072, ZN => n24);
   U44 : AOI22_X1 port map( A1 => din0(26), A2 => net139420, B1 => din1(26), B2
                           => net134072, ZN => n23);
   U45 : AOI22_X1 port map( A1 => din0(25), A2 => net139420, B1 => din1(25), B2
                           => net134074, ZN => n22);
   U46 : AOI22_X1 port map( A1 => din0(23), A2 => net139420, B1 => din1(23), B2
                           => net134078, ZN => n20);
   U47 : AOI22_X1 port map( A1 => din0(22), A2 => net139420, B1 => din1(22), B2
                           => net134078, ZN => n19);
   U48 : AOI22_X1 port map( A1 => din0(21), A2 => net139420, B1 => din1(21), B2
                           => net134074, ZN => n18);
   U49 : AOI22_X1 port map( A1 => din0(7), A2 => net139420, B1 => din1(7), B2 
                           => net134068, ZN => n33);
   U50 : AOI22_X1 port map( A1 => din0(6), A2 => net139420, B1 => din1(6), B2 
                           => net134068, ZN => n32);
   U51 : AOI22_X1 port map( A1 => din0(3), A2 => net139420, B1 => din1(3), B2 
                           => net153543, ZN => n29);
   U52 : AOI22_X1 port map( A1 => din0(2), A2 => n1, B1 => din1(2), B2 => 
                           net134076, ZN => n26);
   U53 : INV_X1 port map( A => n16, ZN => dout(1));
   U54 : AOI22_X1 port map( A1 => din0(31), A2 => net134066, B1 => din1(31), B2
                           => net134070, ZN => n28);
   U55 : AOI22_X1 port map( A1 => din0(30), A2 => net134066, B1 => din1(30), B2
                           => net134078, ZN => n27);
   U56 : AOI22_X1 port map( A1 => din0(24), A2 => net134066, B1 => din1(24), B2
                           => net134074, ZN => n21);
   U57 : AOI22_X1 port map( A1 => din0(20), A2 => net134066, B1 => din1(20), B2
                           => net134078, ZN => n17);
   U58 : AOI22_X1 port map( A1 => din0(9), A2 => net134066, B1 => net134074, B2
                           => din1(9), ZN => n36);
   U59 : AOI22_X1 port map( A1 => din0(8), A2 => net134066, B1 => din1(8), B2 
                           => net134068, ZN => n35);
   U60 : AOI22_X1 port map( A1 => din0(4), A2 => net134066, B1 => din1(4), B2 
                           => net153543, ZN => n30);
   U61 : INV_X1 port map( A => n31, ZN => dout(5));
   U62 : AOI22_X1 port map( A1 => din0(5), A2 => net134066, B1 => din1(5), B2 
                           => net134068, ZN => n31);
   U63 : AOI22_X1 port map( A1 => din0(28), A2 => net134066, B1 => din1(28), B2
                           => net134072, ZN => n25);
   U64 : INV_X1 port map( A => n25, ZN => dout(28));
   U65 : CLKBUF_X1 port map( A => net153543, Z => net134072);
   U66 : AOI22_X1 port map( A1 => din0(19), A2 => net139420, B1 => din1(19), B2
                           => net134074, ZN => n15);
   U67 : AOI22_X1 port map( A1 => din0(15), A2 => net139420, B1 => din1(15), B2
                           => net134080, ZN => n11);
   U68 : AOI22_X1 port map( A1 => din0(18), A2 => net134066, B1 => din1(18), B2
                           => net134078, ZN => n14);
   U69 : AOI22_X1 port map( A1 => din0(16), A2 => net139420, B1 => din1(16), B2
                           => net134074, ZN => n12);
   U70 : AOI22_X1 port map( A1 => din0(14), A2 => net139420, B1 => din1(14), B2
                           => net134080, ZN => n10);
   U71 : AOI22_X1 port map( A1 => din0(17), A2 => net139420, B1 => din1(17), B2
                           => net134078, ZN => n13);
   U72 : AOI22_X1 port map( A1 => din0(13), A2 => net139420, B1 => din1(13), B2
                           => net134080, ZN => n9);
   U73 : AOI22_X1 port map( A1 => din0(12), A2 => net134066, B1 => din1(12), B2
                           => net134080, ZN => n8);
   U74 : AOI22_X1 port map( A1 => din0(11), A2 => net139420, B1 => din1(11), B2
                           => net134072, ZN => n7);
   U75 : AOI22_X1 port map( A1 => din0(10), A2 => net134066, B1 => din1(10), B2
                           => net134074, ZN => n6);
   U76 : AOI22_X1 port map( A1 => din0(1), A2 => net139419, B1 => din1(1), B2 
                           => n2, ZN => n16);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE32_8 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0);  
         dout : out std_logic_vector (31 downto 0));

end Mux_DATA_SIZE32_8;

architecture SYN_mux_arch of Mux_DATA_SIZE32_8 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n14, ZN => n4);
   U2 : INV_X1 port map( A => n14, ZN => n5);
   U3 : BUF_X1 port map( A => n3, Z => n14);
   U4 : BUF_X1 port map( A => n1, Z => n6);
   U5 : BUF_X1 port map( A => n3, Z => n12);
   U6 : BUF_X1 port map( A => n2, Z => n11);
   U7 : BUF_X1 port map( A => n2, Z => n9);
   U8 : BUF_X1 port map( A => n2, Z => n10);
   U9 : BUF_X1 port map( A => n1, Z => n7);
   U10 : BUF_X1 port map( A => n3, Z => n13);
   U11 : BUF_X1 port map( A => n1, Z => n8);
   U12 : INV_X1 port map( A => n48, ZN => dout(29));
   U13 : INV_X1 port map( A => n50, ZN => dout(30));
   U14 : AOI22_X1 port map( A1 => din0(30), A2 => n5, B1 => din1(30), B2 => n10
                           , ZN => n50);
   U15 : INV_X1 port map( A => n47, ZN => dout(28));
   U16 : INV_X1 port map( A => n31, ZN => dout(24));
   U17 : AOI22_X1 port map( A1 => din0(24), A2 => n5, B1 => din1(24), B2 => n9,
                           ZN => n31);
   U18 : INV_X1 port map( A => n32, ZN => dout(25));
   U19 : AOI22_X1 port map( A1 => din0(25), A2 => n5, B1 => din1(25), B2 => n9,
                           ZN => n32);
   U20 : INV_X1 port map( A => n33, ZN => dout(26));
   U21 : AOI22_X1 port map( A1 => din0(26), A2 => n5, B1 => din1(26), B2 => n8,
                           ZN => n33);
   U22 : INV_X1 port map( A => n35, ZN => dout(27));
   U23 : AOI22_X1 port map( A1 => din0(27), A2 => n5, B1 => din1(27), B2 => n8,
                           ZN => n35);
   U24 : INV_X1 port map( A => n15, ZN => dout(0));
   U25 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => n13, 
                           ZN => n15);
   U26 : INV_X1 port map( A => n26, ZN => dout(1));
   U27 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => n10, 
                           ZN => n26);
   U28 : INV_X1 port map( A => n49, ZN => dout(2));
   U29 : AOI22_X1 port map( A1 => din0(2), A2 => n5, B1 => din1(2), B2 => n7, 
                           ZN => n49);
   U30 : INV_X1 port map( A => n52, ZN => dout(3));
   U31 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => din1(3), B2 => n7, 
                           ZN => n52);
   U32 : INV_X1 port map( A => n53, ZN => dout(4));
   U33 : AOI22_X1 port map( A1 => din0(4), A2 => n5, B1 => din1(4), B2 => n7, 
                           ZN => n53);
   U34 : INV_X1 port map( A => n55, ZN => dout(6));
   U35 : AOI22_X1 port map( A1 => din0(6), A2 => n5, B1 => din1(6), B2 => n6, 
                           ZN => n55);
   U36 : INV_X1 port map( A => n56, ZN => dout(7));
   U37 : AOI22_X1 port map( A1 => din0(7), A2 => n5, B1 => din1(7), B2 => n6, 
                           ZN => n56);
   U38 : INV_X1 port map( A => n57, ZN => dout(8));
   U39 : AOI22_X1 port map( A1 => din0(8), A2 => n4, B1 => din1(8), B2 => n6, 
                           ZN => n57);
   U40 : INV_X1 port map( A => n58, ZN => dout(9));
   U41 : AOI22_X1 port map( A1 => din0(9), A2 => n4, B1 => n13, B2 => din1(9), 
                           ZN => n58);
   U42 : INV_X1 port map( A => n16, ZN => dout(10));
   U43 : AOI22_X1 port map( A1 => din0(10), A2 => n4, B1 => din1(10), B2 => n13
                           , ZN => n16);
   U44 : INV_X1 port map( A => n17, ZN => dout(11));
   U45 : AOI22_X1 port map( A1 => din0(11), A2 => n4, B1 => din1(11), B2 => n13
                           , ZN => n17);
   U46 : INV_X1 port map( A => n18, ZN => dout(12));
   U47 : AOI22_X1 port map( A1 => din0(12), A2 => n4, B1 => din1(12), B2 => n12
                           , ZN => n18);
   U48 : INV_X1 port map( A => n19, ZN => dout(13));
   U49 : AOI22_X1 port map( A1 => din0(13), A2 => n4, B1 => din1(13), B2 => n12
                           , ZN => n19);
   U50 : INV_X1 port map( A => n20, ZN => dout(14));
   U51 : AOI22_X1 port map( A1 => din0(14), A2 => n4, B1 => din1(14), B2 => n12
                           , ZN => n20);
   U52 : INV_X1 port map( A => n21, ZN => dout(15));
   U53 : AOI22_X1 port map( A1 => din0(15), A2 => n4, B1 => din1(15), B2 => n12
                           , ZN => n21);
   U54 : INV_X1 port map( A => n22, ZN => dout(16));
   U55 : AOI22_X1 port map( A1 => din0(16), A2 => n4, B1 => din1(16), B2 => n11
                           , ZN => n22);
   U56 : INV_X1 port map( A => n23, ZN => dout(17));
   U57 : AOI22_X1 port map( A1 => din0(17), A2 => n4, B1 => din1(17), B2 => n11
                           , ZN => n23);
   U58 : INV_X1 port map( A => n24, ZN => dout(18));
   U59 : AOI22_X1 port map( A1 => din0(18), A2 => n4, B1 => din1(18), B2 => n11
                           , ZN => n24);
   U60 : INV_X1 port map( A => n25, ZN => dout(19));
   U61 : AOI22_X1 port map( A1 => din0(19), A2 => n4, B1 => din1(19), B2 => n11
                           , ZN => n25);
   U62 : INV_X1 port map( A => n27, ZN => dout(20));
   U63 : AOI22_X1 port map( A1 => din0(20), A2 => n5, B1 => din1(20), B2 => n10
                           , ZN => n27);
   U64 : INV_X1 port map( A => n28, ZN => dout(21));
   U65 : AOI22_X1 port map( A1 => din0(21), A2 => n5, B1 => din1(21), B2 => n10
                           , ZN => n28);
   U66 : INV_X1 port map( A => n29, ZN => dout(22));
   U67 : AOI22_X1 port map( A1 => din0(22), A2 => n5, B1 => din1(22), B2 => n9,
                           ZN => n29);
   U68 : INV_X1 port map( A => n51, ZN => dout(31));
   U69 : AOI22_X1 port map( A1 => din0(31), A2 => n4, B1 => din1(31), B2 => n7,
                           ZN => n51);
   U70 : INV_X1 port map( A => n30, ZN => dout(23));
   U71 : AOI22_X1 port map( A1 => din0(23), A2 => n5, B1 => din1(23), B2 => n9,
                           ZN => n30);
   U72 : INV_X1 port map( A => n54, ZN => dout(5));
   U73 : AOI22_X1 port map( A1 => din0(5), A2 => n5, B1 => din1(5), B2 => n6, 
                           ZN => n54);
   U74 : AOI22_X1 port map( A1 => din0(29), A2 => n5, B1 => din1(29), B2 => n8,
                           ZN => n48);
   U75 : AOI22_X1 port map( A1 => din0(28), A2 => n5, B1 => din1(28), B2 => n8,
                           ZN => n47);
   U76 : CLKBUF_X1 port map( A => sel, Z => n3);
   U77 : CLKBUF_X1 port map( A => sel, Z => n2);
   U78 : CLKBUF_X1 port map( A => sel, Z => n1);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE32_7 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0);  
         dout : out std_logic_vector (31 downto 0));

end Mux_DATA_SIZE32_7;

architecture SYN_mux_arch of Mux_DATA_SIZE32_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33 : std_logic;

begin
   
   U1 : AOI21_X1 port map( B1 => din1(0), B2 => sel, A => din0(0), ZN => n1);
   U2 : INV_X1 port map( A => n27, ZN => dout(4));
   U3 : INV_X1 port map( A => sel, ZN => n32);
   U4 : INV_X1 port map( A => n26, ZN => dout(3));
   U5 : INV_X1 port map( A => n23, ZN => dout(2));
   U6 : INV_X1 port map( A => n12, ZN => dout(1));
   U7 : INV_X1 port map( A => n10, ZN => dout(18));
   U8 : INV_X1 port map( A => n8, ZN => dout(16));
   U9 : INV_X1 port map( A => n11, ZN => dout(19));
   U10 : INV_X1 port map( A => n4, ZN => dout(12));
   U11 : INV_X1 port map( A => n30, ZN => dout(7));
   U12 : AOI22_X1 port map( A1 => din0(7), A2 => n32, B1 => din1(7), B2 => sel,
                           ZN => n30);
   U13 : INV_X1 port map( A => n2, ZN => dout(10));
   U14 : INV_X1 port map( A => n22, ZN => dout(29));
   U15 : AOI22_X1 port map( A1 => din0(29), A2 => n32, B1 => din1(29), B2 => 
                           sel, ZN => n22);
   U16 : INV_X1 port map( A => n33, ZN => dout(9));
   U17 : AOI22_X1 port map( A1 => din0(9), A2 => n32, B1 => sel, B2 => din1(9),
                           ZN => n33);
   U18 : INV_X1 port map( A => n18, ZN => dout(25));
   U19 : AOI22_X1 port map( A1 => din0(25), A2 => n32, B1 => din1(25), B2 => 
                           sel, ZN => n18);
   U20 : INV_X1 port map( A => n16, ZN => dout(23));
   U21 : AOI22_X1 port map( A1 => din0(23), A2 => n32, B1 => din1(23), B2 => 
                           sel, ZN => n16);
   U22 : INV_X1 port map( A => n20, ZN => dout(27));
   U23 : AOI22_X1 port map( A1 => din0(27), A2 => n32, B1 => din1(27), B2 => 
                           sel, ZN => n20);
   U24 : INV_X1 port map( A => n19, ZN => dout(26));
   U25 : AOI22_X1 port map( A1 => din0(26), A2 => n32, B1 => din1(26), B2 => 
                           sel, ZN => n19);
   U26 : INV_X1 port map( A => n7, ZN => dout(15));
   U27 : AOI22_X1 port map( A1 => din0(3), A2 => n32, B1 => din1(3), B2 => sel,
                           ZN => n26);
   U28 : INV_X1 port map( A => n14, ZN => dout(21));
   U29 : AOI22_X1 port map( A1 => din0(21), A2 => n32, B1 => din1(21), B2 => 
                           sel, ZN => n14);
   U30 : INV_X1 port map( A => n3, ZN => dout(11));
   U31 : INV_X1 port map( A => n29, ZN => dout(6));
   U32 : AOI22_X1 port map( A1 => din0(6), A2 => n32, B1 => din1(6), B2 => sel,
                           ZN => n29);
   U33 : INV_X1 port map( A => n9, ZN => dout(17));
   U34 : INV_X1 port map( A => n6, ZN => dout(14));
   U35 : INV_X1 port map( A => n17, ZN => dout(24));
   U36 : AOI22_X1 port map( A1 => din0(24), A2 => n32, B1 => din1(24), B2 => 
                           sel, ZN => n17);
   U37 : INV_X1 port map( A => n31, ZN => dout(8));
   U38 : AOI22_X1 port map( A1 => din0(8), A2 => n32, B1 => din1(8), B2 => sel,
                           ZN => n31);
   U39 : INV_X1 port map( A => n13, ZN => dout(20));
   U40 : AOI22_X1 port map( A1 => din0(20), A2 => n32, B1 => din1(20), B2 => 
                           sel, ZN => n13);
   U41 : INV_X1 port map( A => n21, ZN => dout(28));
   U42 : AOI22_X1 port map( A1 => din0(28), A2 => n32, B1 => din1(28), B2 => 
                           sel, ZN => n21);
   U43 : INV_X1 port map( A => n15, ZN => dout(22));
   U44 : AOI22_X1 port map( A1 => din0(22), A2 => n32, B1 => din1(22), B2 => 
                           sel, ZN => n15);
   U45 : AOI22_X1 port map( A1 => din0(2), A2 => n32, B1 => din1(2), B2 => sel,
                           ZN => n23);
   U46 : AOI22_X1 port map( A1 => din0(1), A2 => n32, B1 => din1(1), B2 => sel,
                           ZN => n12);
   U47 : INV_X1 port map( A => n28, ZN => dout(5));
   U48 : AOI22_X1 port map( A1 => din0(5), A2 => n32, B1 => din1(5), B2 => sel,
                           ZN => n28);
   U49 : AOI22_X1 port map( A1 => din0(4), A2 => n32, B1 => din1(4), B2 => sel,
                           ZN => n27);
   U50 : INV_X1 port map( A => n24, ZN => dout(30));
   U51 : AOI22_X1 port map( A1 => din0(30), A2 => n32, B1 => din1(30), B2 => 
                           sel, ZN => n24);
   U52 : INV_X1 port map( A => n25, ZN => dout(31));
   U53 : AOI22_X1 port map( A1 => din0(31), A2 => n32, B1 => din1(31), B2 => 
                           sel, ZN => n25);
   U54 : AOI21_X1 port map( B1 => din1(18), B2 => sel, A => din0(18), ZN => n10
                           );
   U55 : AOI21_X1 port map( B1 => din1(19), B2 => sel, A => din0(19), ZN => n11
                           );
   U56 : AOI21_X1 port map( B1 => din1(17), B2 => sel, A => din0(17), ZN => n9)
                           ;
   U57 : AOI21_X1 port map( B1 => din1(15), B2 => sel, A => din0(15), ZN => n7)
                           ;
   U58 : AOI21_X1 port map( B1 => din1(14), B2 => sel, A => din0(14), ZN => n6)
                           ;
   U59 : AOI21_X1 port map( B1 => din1(13), B2 => sel, A => din0(13), ZN => n5)
                           ;
   U60 : AOI21_X1 port map( B1 => din1(12), B2 => sel, A => din0(12), ZN => n4)
                           ;
   U61 : AOI21_X1 port map( B1 => din1(10), B2 => sel, A => din0(10), ZN => n2)
                           ;
   U62 : AOI21_X1 port map( B1 => din1(11), B2 => sel, A => din0(11), ZN => n3)
                           ;
   U63 : AOI21_X1 port map( B1 => din1(16), B2 => sel, A => din0(16), ZN => n8)
                           ;
   U64 : INV_X1 port map( A => n5, ZN => dout(13));
   U65 : INV_X1 port map( A => n1, ZN => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE32_6 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0);  
         dout : out std_logic_vector (31 downto 0));

end Mux_DATA_SIZE32_6;

architecture SYN_mux_arch of Mux_DATA_SIZE32_6 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n35 : std_logic;

begin
   
   U1 : INV_X1 port map( A => sel, ZN => n33);
   U2 : AND2_X1 port map( A1 => din1(17), A2 => sel, ZN => n2);
   U3 : OR2_X1 port map( A1 => n2, A2 => din0(17), ZN => dout(17));
   U4 : INV_X1 port map( A => n26, ZN => dout(31));
   U5 : INV_X1 port map( A => n6, ZN => dout(12));
   U6 : INV_X1 port map( A => n19, ZN => dout(25));
   U7 : AOI22_X1 port map( A1 => din0(25), A2 => n33, B1 => din1(25), B2 => sel
                           , ZN => n19);
   U8 : INV_X1 port map( A => n20, ZN => dout(26));
   U9 : AOI22_X1 port map( A1 => din0(26), A2 => n33, B1 => din1(26), B2 => sel
                           , ZN => n20);
   U10 : INV_X1 port map( A => n18, ZN => dout(24));
   U11 : AOI22_X1 port map( A1 => din0(24), A2 => n33, B1 => din1(24), B2 => 
                           sel, ZN => n18);
   U12 : INV_X1 port map( A => n35, ZN => dout(9));
   U13 : AOI22_X1 port map( A1 => din0(9), A2 => n33, B1 => sel, B2 => din1(9),
                           ZN => n35);
   U14 : INV_X1 port map( A => n31, ZN => dout(7));
   U15 : AOI22_X1 port map( A1 => din0(7), A2 => n33, B1 => din1(7), B2 => sel,
                           ZN => n31);
   U16 : INV_X1 port map( A => n30, ZN => dout(6));
   U17 : AOI22_X1 port map( A1 => din0(6), A2 => n33, B1 => din1(6), B2 => sel,
                           ZN => n30);
   U18 : INV_X1 port map( A => n29, ZN => dout(5));
   U19 : AOI22_X1 port map( A1 => din0(5), A2 => n33, B1 => din1(5), B2 => sel,
                           ZN => n29);
   U20 : INV_X1 port map( A => n27, ZN => dout(3));
   U21 : AOI22_X1 port map( A1 => din0(3), A2 => n33, B1 => din1(3), B2 => sel,
                           ZN => n27);
   U22 : INV_X1 port map( A => n28, ZN => dout(4));
   U23 : AOI22_X1 port map( A1 => din0(4), A2 => n33, B1 => din1(4), B2 => sel,
                           ZN => n28);
   U24 : INV_X1 port map( A => n24, ZN => dout(2));
   U25 : AOI22_X1 port map( A1 => din0(2), A2 => n33, B1 => din1(2), B2 => sel,
                           ZN => n24);
   U26 : INV_X1 port map( A => n13, ZN => dout(1));
   U27 : AOI22_X1 port map( A1 => din0(1), A2 => n33, B1 => din1(1), B2 => sel,
                           ZN => n13);
   U28 : INV_X1 port map( A => n15, ZN => dout(21));
   U29 : AOI22_X1 port map( A1 => din0(21), A2 => n33, B1 => din1(21), B2 => 
                           sel, ZN => n15);
   U30 : INV_X1 port map( A => n14, ZN => dout(20));
   U31 : AOI22_X1 port map( A1 => din0(20), A2 => n33, B1 => din1(20), B2 => 
                           sel, ZN => n14);
   U32 : INV_X1 port map( A => n16, ZN => dout(22));
   U33 : AOI22_X1 port map( A1 => din0(22), A2 => n33, B1 => din1(22), B2 => 
                           sel, ZN => n16);
   U34 : INV_X1 port map( A => n17, ZN => dout(23));
   U35 : AOI22_X1 port map( A1 => din0(23), A2 => n33, B1 => din1(23), B2 => 
                           sel, ZN => n17);
   U36 : INV_X1 port map( A => n32, ZN => dout(8));
   U37 : AOI22_X1 port map( A1 => din0(8), A2 => n33, B1 => din1(8), B2 => sel,
                           ZN => n32);
   U38 : INV_X1 port map( A => n11, ZN => dout(18));
   U39 : INV_X1 port map( A => n8, ZN => dout(14));
   U40 : INV_X1 port map( A => n4, ZN => dout(10));
   U41 : INV_X1 port map( A => n5, ZN => dout(11));
   U42 : INV_X1 port map( A => n3, ZN => dout(0));
   U43 : INV_X1 port map( A => n10, ZN => dout(16));
   U44 : INV_X1 port map( A => n12, ZN => dout(19));
   U45 : INV_X1 port map( A => n9, ZN => dout(15));
   U46 : AOI22_X1 port map( A1 => din0(27), A2 => n33, B1 => din1(27), B2 => 
                           sel, ZN => n21);
   U47 : AOI22_X1 port map( A1 => din0(31), A2 => n33, B1 => din1(31), B2 => 
                           sel, ZN => n26);
   U48 : AOI21_X1 port map( B1 => din1(0), B2 => sel, A => din0(0), ZN => n3);
   U49 : AOI21_X1 port map( B1 => din1(10), B2 => sel, A => din0(10), ZN => n4)
                           ;
   U50 : AOI21_X1 port map( B1 => din1(11), B2 => sel, A => din0(11), ZN => n5)
                           ;
   U51 : AOI21_X1 port map( B1 => din1(12), B2 => sel, A => din0(12), ZN => n6)
                           ;
   U52 : AOI21_X1 port map( B1 => din1(13), B2 => sel, A => din0(13), ZN => n7)
                           ;
   U53 : AOI21_X1 port map( B1 => din1(14), B2 => sel, A => din0(14), ZN => n8)
                           ;
   U54 : AOI21_X1 port map( B1 => din1(15), B2 => sel, A => din0(15), ZN => n9)
                           ;
   U55 : AOI21_X1 port map( B1 => din1(16), B2 => sel, A => din0(16), ZN => n10
                           );
   U56 : AOI21_X1 port map( B1 => din1(18), B2 => sel, A => din0(18), ZN => n11
                           );
   U57 : AOI21_X1 port map( B1 => din1(19), B2 => sel, A => din0(19), ZN => n12
                           );
   U58 : AOI22_X1 port map( A1 => din0(29), A2 => n33, B1 => din1(29), B2 => 
                           sel, ZN => n23);
   U59 : AOI22_X1 port map( A1 => din0(30), A2 => n33, B1 => din1(30), B2 => 
                           sel, ZN => n25);
   U60 : INV_X1 port map( A => n25, ZN => dout(30));
   U61 : INV_X1 port map( A => n23, ZN => dout(29));
   U62 : INV_X1 port map( A => n7, ZN => dout(13));
   U63 : INV_X1 port map( A => n21, ZN => dout(27));
   U64 : INV_X1 port map( A => n22, ZN => dout(28));
   U65 : AOI22_X1 port map( A1 => din0(28), A2 => n33, B1 => din1(28), B2 => 
                           sel, ZN => n22);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE32_5 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0);  
         dout : out std_logic_vector (31 downto 0));

end Mux_DATA_SIZE32_5;

architecture SYN_mux_arch of Mux_DATA_SIZE32_5 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n14, ZN => n4);
   U2 : INV_X1 port map( A => n14, ZN => n5);
   U3 : BUF_X1 port map( A => n1, Z => n6);
   U4 : BUF_X1 port map( A => n3, Z => n12);
   U5 : BUF_X1 port map( A => n2, Z => n11);
   U6 : BUF_X1 port map( A => n2, Z => n9);
   U7 : BUF_X1 port map( A => n1, Z => n8);
   U8 : BUF_X1 port map( A => n2, Z => n10);
   U9 : BUF_X1 port map( A => n1, Z => n7);
   U10 : BUF_X1 port map( A => n3, Z => n14);
   U11 : BUF_X1 port map( A => n3, Z => n13);
   U12 : INV_X1 port map( A => n58, ZN => dout(9));
   U13 : AOI22_X1 port map( A1 => din0(9), A2 => n4, B1 => n13, B2 => din1(9), 
                           ZN => n58);
   U14 : INV_X1 port map( A => n26, ZN => dout(1));
   U15 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => n10, 
                           ZN => n26);
   U16 : INV_X1 port map( A => n15, ZN => dout(0));
   U17 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => n13, 
                           ZN => n15);
   U18 : INV_X1 port map( A => n49, ZN => dout(2));
   U19 : AOI22_X1 port map( A1 => din0(2), A2 => n5, B1 => din1(2), B2 => n7, 
                           ZN => n49);
   U20 : INV_X1 port map( A => n54, ZN => dout(5));
   U21 : AOI22_X1 port map( A1 => din0(5), A2 => n5, B1 => din1(5), B2 => n6, 
                           ZN => n54);
   U22 : INV_X1 port map( A => n57, ZN => dout(8));
   U23 : AOI22_X1 port map( A1 => din0(8), A2 => n4, B1 => din1(8), B2 => n6, 
                           ZN => n57);
   U24 : INV_X1 port map( A => n16, ZN => dout(10));
   U25 : AOI22_X1 port map( A1 => din0(10), A2 => n4, B1 => din1(10), B2 => n13
                           , ZN => n16);
   U26 : INV_X1 port map( A => n20, ZN => dout(14));
   U27 : AOI22_X1 port map( A1 => din0(14), A2 => n4, B1 => din1(14), B2 => n12
                           , ZN => n20);
   U28 : INV_X1 port map( A => n52, ZN => dout(3));
   U29 : AOI22_X1 port map( A1 => din0(3), A2 => n5, B1 => din1(3), B2 => n7, 
                           ZN => n52);
   U30 : INV_X1 port map( A => n19, ZN => dout(13));
   U31 : AOI22_X1 port map( A1 => din0(13), A2 => n4, B1 => din1(13), B2 => n12
                           , ZN => n19);
   U32 : INV_X1 port map( A => n56, ZN => dout(7));
   U33 : AOI22_X1 port map( A1 => din0(7), A2 => n4, B1 => din1(7), B2 => n6, 
                           ZN => n56);
   U34 : INV_X1 port map( A => n21, ZN => dout(15));
   U35 : AOI22_X1 port map( A1 => din0(15), A2 => n4, B1 => din1(15), B2 => n12
                           , ZN => n21);
   U36 : INV_X1 port map( A => n17, ZN => dout(11));
   U37 : AOI22_X1 port map( A1 => din0(11), A2 => n4, B1 => din1(11), B2 => n13
                           , ZN => n17);
   U38 : INV_X1 port map( A => n55, ZN => dout(6));
   U39 : AOI22_X1 port map( A1 => din0(6), A2 => n5, B1 => din1(6), B2 => n6, 
                           ZN => n55);
   U40 : INV_X1 port map( A => n53, ZN => dout(4));
   U41 : AOI22_X1 port map( A1 => din0(4), A2 => n4, B1 => din1(4), B2 => n7, 
                           ZN => n53);
   U42 : INV_X1 port map( A => n18, ZN => dout(12));
   U43 : AOI22_X1 port map( A1 => din0(12), A2 => n4, B1 => din1(12), B2 => n12
                           , ZN => n18);
   U44 : INV_X1 port map( A => n29, ZN => dout(22));
   U45 : AOI22_X1 port map( A1 => din0(22), A2 => n5, B1 => din1(22), B2 => n9,
                           ZN => n29);
   U46 : INV_X1 port map( A => n30, ZN => dout(23));
   U47 : AOI22_X1 port map( A1 => din0(23), A2 => n5, B1 => din1(23), B2 => n9,
                           ZN => n30);
   U48 : INV_X1 port map( A => n31, ZN => dout(24));
   U49 : AOI22_X1 port map( A1 => din0(24), A2 => n5, B1 => din1(24), B2 => n9,
                           ZN => n31);
   U50 : INV_X1 port map( A => n32, ZN => dout(25));
   U51 : AOI22_X1 port map( A1 => din0(25), A2 => n5, B1 => din1(25), B2 => n9,
                           ZN => n32);
   U52 : INV_X1 port map( A => n33, ZN => dout(26));
   U53 : AOI22_X1 port map( A1 => din0(26), A2 => n5, B1 => din1(26), B2 => n8,
                           ZN => n33);
   U54 : INV_X1 port map( A => n35, ZN => dout(27));
   U55 : AOI22_X1 port map( A1 => din0(27), A2 => n5, B1 => din1(27), B2 => n8,
                           ZN => n35);
   U56 : INV_X1 port map( A => n47, ZN => dout(28));
   U57 : AOI22_X1 port map( A1 => din0(28), A2 => n5, B1 => din1(28), B2 => n8,
                           ZN => n47);
   U58 : INV_X1 port map( A => n48, ZN => dout(29));
   U59 : AOI22_X1 port map( A1 => din0(29), A2 => n5, B1 => din1(29), B2 => n8,
                           ZN => n48);
   U60 : INV_X1 port map( A => n22, ZN => dout(16));
   U61 : AOI22_X1 port map( A1 => din0(16), A2 => n4, B1 => din1(16), B2 => n11
                           , ZN => n22);
   U62 : INV_X1 port map( A => n23, ZN => dout(17));
   U63 : AOI22_X1 port map( A1 => din0(17), A2 => n4, B1 => din1(17), B2 => n11
                           , ZN => n23);
   U64 : INV_X1 port map( A => n24, ZN => dout(18));
   U65 : AOI22_X1 port map( A1 => din0(18), A2 => n4, B1 => din1(18), B2 => n11
                           , ZN => n24);
   U66 : INV_X1 port map( A => n25, ZN => dout(19));
   U67 : AOI22_X1 port map( A1 => din0(19), A2 => n4, B1 => din1(19), B2 => n11
                           , ZN => n25);
   U68 : INV_X1 port map( A => n27, ZN => dout(20));
   U69 : AOI22_X1 port map( A1 => din0(20), A2 => n5, B1 => din1(20), B2 => n10
                           , ZN => n27);
   U70 : INV_X1 port map( A => n28, ZN => dout(21));
   U71 : AOI22_X1 port map( A1 => din0(21), A2 => n5, B1 => din1(21), B2 => n10
                           , ZN => n28);
   U72 : INV_X1 port map( A => n50, ZN => dout(30));
   U73 : AOI22_X1 port map( A1 => din0(30), A2 => n5, B1 => din1(30), B2 => n10
                           , ZN => n50);
   U74 : INV_X1 port map( A => n51, ZN => dout(31));
   U75 : AOI22_X1 port map( A1 => din0(31), A2 => n5, B1 => din1(31), B2 => n7,
                           ZN => n51);
   U76 : BUF_X1 port map( A => sel, Z => n3);
   U77 : BUF_X1 port map( A => sel, Z => n2);
   U78 : BUF_X1 port map( A => sel, Z => n1);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE32_4 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0);  
         dout : out std_logic_vector (31 downto 0));

end Mux_DATA_SIZE32_4;

architecture SYN_mux_arch of Mux_DATA_SIZE32_4 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n14, ZN => n4);
   U2 : INV_X1 port map( A => n14, ZN => n5);
   U3 : BUF_X1 port map( A => n1, Z => n6);
   U4 : BUF_X1 port map( A => n3, Z => n12);
   U5 : BUF_X1 port map( A => n2, Z => n11);
   U6 : BUF_X1 port map( A => n2, Z => n9);
   U7 : BUF_X1 port map( A => n1, Z => n8);
   U8 : BUF_X1 port map( A => n2, Z => n10);
   U9 : BUF_X1 port map( A => n1, Z => n7);
   U10 : BUF_X1 port map( A => n3, Z => n14);
   U11 : BUF_X1 port map( A => n3, Z => n13);
   U12 : INV_X1 port map( A => n29, ZN => dout(22));
   U13 : AOI22_X1 port map( A1 => din0(22), A2 => n5, B1 => din1(22), B2 => n9,
                           ZN => n29);
   U14 : INV_X1 port map( A => n30, ZN => dout(23));
   U15 : AOI22_X1 port map( A1 => din0(23), A2 => n5, B1 => din1(23), B2 => n9,
                           ZN => n30);
   U16 : INV_X1 port map( A => n31, ZN => dout(24));
   U17 : AOI22_X1 port map( A1 => din0(24), A2 => n5, B1 => din1(24), B2 => n9,
                           ZN => n31);
   U18 : INV_X1 port map( A => n32, ZN => dout(25));
   U19 : AOI22_X1 port map( A1 => din0(25), A2 => n5, B1 => din1(25), B2 => n9,
                           ZN => n32);
   U20 : INV_X1 port map( A => n33, ZN => dout(26));
   U21 : AOI22_X1 port map( A1 => din0(26), A2 => n5, B1 => din1(26), B2 => n8,
                           ZN => n33);
   U22 : INV_X1 port map( A => n35, ZN => dout(27));
   U23 : AOI22_X1 port map( A1 => din0(27), A2 => n5, B1 => din1(27), B2 => n8,
                           ZN => n35);
   U24 : INV_X1 port map( A => n47, ZN => dout(28));
   U25 : AOI22_X1 port map( A1 => din0(28), A2 => n5, B1 => din1(28), B2 => n8,
                           ZN => n47);
   U26 : INV_X1 port map( A => n48, ZN => dout(29));
   U27 : AOI22_X1 port map( A1 => din0(29), A2 => n5, B1 => din1(29), B2 => n8,
                           ZN => n48);
   U28 : INV_X1 port map( A => n15, ZN => dout(0));
   U29 : AOI22_X1 port map( A1 => din0(0), A2 => n4, B1 => din1(0), B2 => n13, 
                           ZN => n15);
   U30 : INV_X1 port map( A => n26, ZN => dout(1));
   U31 : AOI22_X1 port map( A1 => din0(1), A2 => n4, B1 => din1(1), B2 => n10, 
                           ZN => n26);
   U32 : INV_X1 port map( A => n49, ZN => dout(2));
   U33 : AOI22_X1 port map( A1 => din0(2), A2 => n5, B1 => din1(2), B2 => n7, 
                           ZN => n49);
   U34 : INV_X1 port map( A => n52, ZN => dout(3));
   U35 : AOI22_X1 port map( A1 => din0(3), A2 => n4, B1 => din1(3), B2 => n7, 
                           ZN => n52);
   U36 : INV_X1 port map( A => n53, ZN => dout(4));
   U37 : AOI22_X1 port map( A1 => din0(4), A2 => n5, B1 => din1(4), B2 => n7, 
                           ZN => n53);
   U38 : INV_X1 port map( A => n54, ZN => dout(5));
   U39 : AOI22_X1 port map( A1 => din0(5), A2 => n4, B1 => din1(5), B2 => n6, 
                           ZN => n54);
   U40 : INV_X1 port map( A => n55, ZN => dout(6));
   U41 : AOI22_X1 port map( A1 => din0(6), A2 => n5, B1 => din1(6), B2 => n6, 
                           ZN => n55);
   U42 : INV_X1 port map( A => n56, ZN => dout(7));
   U43 : AOI22_X1 port map( A1 => din0(7), A2 => n4, B1 => din1(7), B2 => n6, 
                           ZN => n56);
   U44 : INV_X1 port map( A => n57, ZN => dout(8));
   U45 : AOI22_X1 port map( A1 => din0(8), A2 => n5, B1 => din1(8), B2 => n6, 
                           ZN => n57);
   U46 : INV_X1 port map( A => n58, ZN => dout(9));
   U47 : AOI22_X1 port map( A1 => din0(9), A2 => n4, B1 => n13, B2 => din1(9), 
                           ZN => n58);
   U48 : INV_X1 port map( A => n16, ZN => dout(10));
   U49 : AOI22_X1 port map( A1 => din0(10), A2 => n4, B1 => din1(10), B2 => n13
                           , ZN => n16);
   U50 : INV_X1 port map( A => n17, ZN => dout(11));
   U51 : AOI22_X1 port map( A1 => din0(11), A2 => n4, B1 => din1(11), B2 => n13
                           , ZN => n17);
   U52 : INV_X1 port map( A => n18, ZN => dout(12));
   U53 : AOI22_X1 port map( A1 => din0(12), A2 => n4, B1 => din1(12), B2 => n12
                           , ZN => n18);
   U54 : INV_X1 port map( A => n19, ZN => dout(13));
   U55 : AOI22_X1 port map( A1 => din0(13), A2 => n4, B1 => din1(13), B2 => n12
                           , ZN => n19);
   U56 : INV_X1 port map( A => n20, ZN => dout(14));
   U57 : AOI22_X1 port map( A1 => din0(14), A2 => n4, B1 => din1(14), B2 => n12
                           , ZN => n20);
   U58 : INV_X1 port map( A => n21, ZN => dout(15));
   U59 : AOI22_X1 port map( A1 => din0(15), A2 => n4, B1 => din1(15), B2 => n12
                           , ZN => n21);
   U60 : INV_X1 port map( A => n22, ZN => dout(16));
   U61 : AOI22_X1 port map( A1 => din0(16), A2 => n4, B1 => din1(16), B2 => n11
                           , ZN => n22);
   U62 : INV_X1 port map( A => n23, ZN => dout(17));
   U63 : AOI22_X1 port map( A1 => din0(17), A2 => n4, B1 => din1(17), B2 => n11
                           , ZN => n23);
   U64 : INV_X1 port map( A => n24, ZN => dout(18));
   U65 : AOI22_X1 port map( A1 => din0(18), A2 => n4, B1 => din1(18), B2 => n11
                           , ZN => n24);
   U66 : INV_X1 port map( A => n25, ZN => dout(19));
   U67 : AOI22_X1 port map( A1 => din0(19), A2 => n4, B1 => din1(19), B2 => n11
                           , ZN => n25);
   U68 : INV_X1 port map( A => n27, ZN => dout(20));
   U69 : AOI22_X1 port map( A1 => din0(20), A2 => n5, B1 => din1(20), B2 => n10
                           , ZN => n27);
   U70 : INV_X1 port map( A => n28, ZN => dout(21));
   U71 : AOI22_X1 port map( A1 => din0(21), A2 => n5, B1 => din1(21), B2 => n10
                           , ZN => n28);
   U72 : INV_X1 port map( A => n50, ZN => dout(30));
   U73 : AOI22_X1 port map( A1 => din0(30), A2 => n5, B1 => din1(30), B2 => n10
                           , ZN => n50);
   U74 : INV_X1 port map( A => n51, ZN => dout(31));
   U75 : AOI22_X1 port map( A1 => din0(31), A2 => n5, B1 => din1(31), B2 => n7,
                           ZN => n51);
   U76 : BUF_X1 port map( A => sel, Z => n3);
   U77 : BUF_X1 port map( A => sel, Z => n2);
   U78 : BUF_X1 port map( A => sel, Z => n1);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE32_2 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0);  
         dout : out std_logic_vector (31 downto 0));

end Mux_DATA_SIZE32_2;

architecture SYN_mux_arch of Mux_DATA_SIZE32_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33 : std_logic;

begin
   
   U1 : INV_X1 port map( A => sel, ZN => n32);
   U2 : INV_X1 port map( A => n12, ZN => dout(1));
   U3 : AOI22_X1 port map( A1 => din0(1), A2 => n32, B1 => din1(1), B2 => sel, 
                           ZN => n12);
   U4 : INV_X1 port map( A => n23, ZN => dout(2));
   U5 : AOI22_X1 port map( A1 => din0(2), A2 => n32, B1 => din1(2), B2 => sel, 
                           ZN => n23);
   U6 : INV_X1 port map( A => n26, ZN => dout(3));
   U7 : AOI22_X1 port map( A1 => din0(3), A2 => n32, B1 => din1(3), B2 => sel, 
                           ZN => n26);
   U8 : INV_X1 port map( A => n27, ZN => dout(4));
   U9 : AOI22_X1 port map( A1 => din0(4), A2 => n32, B1 => din1(4), B2 => sel, 
                           ZN => n27);
   U10 : INV_X1 port map( A => n28, ZN => dout(5));
   U11 : AOI22_X1 port map( A1 => din0(5), A2 => n32, B1 => din1(5), B2 => sel,
                           ZN => n28);
   U12 : INV_X1 port map( A => n29, ZN => dout(6));
   U13 : AOI22_X1 port map( A1 => din0(6), A2 => n32, B1 => din1(6), B2 => sel,
                           ZN => n29);
   U14 : INV_X1 port map( A => n30, ZN => dout(7));
   U15 : AOI22_X1 port map( A1 => din0(7), A2 => n32, B1 => din1(7), B2 => sel,
                           ZN => n30);
   U16 : INV_X1 port map( A => n31, ZN => dout(8));
   U17 : AOI22_X1 port map( A1 => din0(8), A2 => n32, B1 => din1(8), B2 => sel,
                           ZN => n31);
   U18 : INV_X1 port map( A => n33, ZN => dout(9));
   U19 : AOI22_X1 port map( A1 => din0(9), A2 => n32, B1 => sel, B2 => din1(9),
                           ZN => n33);
   U20 : INV_X1 port map( A => n13, ZN => dout(20));
   U21 : AOI22_X1 port map( A1 => din0(20), A2 => n32, B1 => din1(20), B2 => 
                           sel, ZN => n13);
   U22 : INV_X1 port map( A => n14, ZN => dout(21));
   U23 : AOI22_X1 port map( A1 => din0(21), A2 => n32, B1 => din1(21), B2 => 
                           sel, ZN => n14);
   U24 : INV_X1 port map( A => n15, ZN => dout(22));
   U25 : AOI22_X1 port map( A1 => din0(22), A2 => n32, B1 => din1(22), B2 => 
                           sel, ZN => n15);
   U26 : INV_X1 port map( A => n16, ZN => dout(23));
   U27 : AOI22_X1 port map( A1 => din0(23), A2 => n32, B1 => din1(23), B2 => 
                           sel, ZN => n16);
   U28 : INV_X1 port map( A => n17, ZN => dout(24));
   U29 : AOI22_X1 port map( A1 => din0(24), A2 => n32, B1 => din1(24), B2 => 
                           sel, ZN => n17);
   U30 : INV_X1 port map( A => n18, ZN => dout(25));
   U31 : AOI22_X1 port map( A1 => din0(25), A2 => n32, B1 => din1(25), B2 => 
                           sel, ZN => n18);
   U32 : INV_X1 port map( A => n19, ZN => dout(26));
   U33 : AOI22_X1 port map( A1 => din0(26), A2 => n32, B1 => din1(26), B2 => 
                           sel, ZN => n19);
   U34 : INV_X1 port map( A => n20, ZN => dout(27));
   U35 : AOI22_X1 port map( A1 => din0(27), A2 => n32, B1 => din1(27), B2 => 
                           sel, ZN => n20);
   U36 : INV_X1 port map( A => n21, ZN => dout(28));
   U37 : AOI22_X1 port map( A1 => din0(28), A2 => n32, B1 => din1(28), B2 => 
                           sel, ZN => n21);
   U38 : INV_X1 port map( A => n22, ZN => dout(29));
   U39 : AOI22_X1 port map( A1 => din0(29), A2 => n32, B1 => din1(29), B2 => 
                           sel, ZN => n22);
   U40 : INV_X1 port map( A => n24, ZN => dout(30));
   U41 : AOI22_X1 port map( A1 => din0(30), A2 => n32, B1 => din1(30), B2 => 
                           sel, ZN => n24);
   U42 : INV_X1 port map( A => n25, ZN => dout(31));
   U43 : AOI22_X1 port map( A1 => din0(31), A2 => n32, B1 => din1(31), B2 => 
                           sel, ZN => n25);
   U44 : INV_X1 port map( A => n2, ZN => dout(10));
   U45 : INV_X1 port map( A => n3, ZN => dout(11));
   U46 : INV_X1 port map( A => n4, ZN => dout(12));
   U47 : INV_X1 port map( A => n5, ZN => dout(13));
   U48 : INV_X1 port map( A => n6, ZN => dout(14));
   U49 : INV_X1 port map( A => n7, ZN => dout(15));
   U50 : INV_X1 port map( A => n8, ZN => dout(16));
   U51 : INV_X1 port map( A => n9, ZN => dout(17));
   U52 : INV_X1 port map( A => n10, ZN => dout(18));
   U53 : INV_X1 port map( A => n11, ZN => dout(19));
   U54 : INV_X1 port map( A => n1, ZN => dout(0));
   U55 : AOI21_X1 port map( B1 => din1(0), B2 => sel, A => din0(0), ZN => n1);
   U56 : AOI21_X1 port map( B1 => din1(10), B2 => sel, A => din0(10), ZN => n2)
                           ;
   U57 : AOI21_X1 port map( B1 => din1(11), B2 => sel, A => din0(11), ZN => n3)
                           ;
   U58 : AOI21_X1 port map( B1 => din1(12), B2 => sel, A => din0(12), ZN => n4)
                           ;
   U59 : AOI21_X1 port map( B1 => din1(13), B2 => sel, A => din0(13), ZN => n5)
                           ;
   U60 : AOI21_X1 port map( B1 => din1(14), B2 => sel, A => din0(14), ZN => n6)
                           ;
   U61 : AOI21_X1 port map( B1 => din1(15), B2 => sel, A => din0(15), ZN => n7)
                           ;
   U62 : AOI21_X1 port map( B1 => din1(16), B2 => sel, A => din0(16), ZN => n8)
                           ;
   U63 : AOI21_X1 port map( B1 => din1(17), B2 => sel, A => din0(17), ZN => n9)
                           ;
   U64 : AOI21_X1 port map( B1 => din1(18), B2 => sel, A => din0(18), ZN => n10
                           );
   U65 : AOI21_X1 port map( B1 => din1(19), B2 => sel, A => din0(19), ZN => n11
                           );

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE32_1 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0);  
         dout : out std_logic_vector (31 downto 0));

end Mux_DATA_SIZE32_1;

architecture SYN_mux_arch of Mux_DATA_SIZE32_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n35, n44, n45, n46, n47, n48, n49, n50, n51, n52 : 
      std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => sel, Z => n1);
   U2 : BUF_X2 port map( A => n5, Z => n9);
   U3 : BUF_X2 port map( A => n1, Z => n5);
   U4 : INV_X1 port map( A => sel, ZN => n2);
   U5 : INV_X2 port map( A => n1, ZN => n3);
   U6 : BUF_X1 port map( A => n1, Z => n6);
   U7 : CLKBUF_X1 port map( A => n5, Z => n11);
   U8 : CLKBUF_X1 port map( A => n7, Z => n10);
   U9 : CLKBUF_X1 port map( A => n11, Z => n8);
   U10 : CLKBUF_X1 port map( A => n1, Z => n7);
   U11 : INV_X1 port map( A => n48, ZN => dout(5));
   U12 : AOI22_X1 port map( A1 => din0(5), A2 => n3, B1 => din1(5), B2 => n5, 
                           ZN => n48);
   U13 : INV_X1 port map( A => n13, ZN => dout(10));
   U14 : AOI22_X1 port map( A1 => din0(10), A2 => n4, B1 => din1(10), B2 => n8,
                           ZN => n13);
   U15 : INV_X1 port map( A => n22, ZN => dout(19));
   U16 : INV_X1 port map( A => n21, ZN => dout(18));
   U17 : INV_X1 port map( A => n25, ZN => dout(21));
   U18 : AOI22_X1 port map( A1 => din0(21), A2 => n4, B1 => din1(21), B2 => n9,
                           ZN => n25);
   U19 : INV_X1 port map( A => n14, ZN => dout(11));
   U20 : AOI22_X1 port map( A1 => din0(11), A2 => n3, B1 => din1(11), B2 => n7,
                           ZN => n14);
   U21 : INV_X1 port map( A => n50, ZN => dout(7));
   U22 : AOI22_X1 port map( A1 => din0(7), A2 => n4, B1 => din1(7), B2 => n5, 
                           ZN => n50);
   U23 : INV_X1 port map( A => n16, ZN => dout(13));
   U24 : AOI22_X1 port map( A1 => din0(13), A2 => n4, B1 => din1(13), B2 => n11
                           , ZN => n16);
   U25 : INV_X1 port map( A => n17, ZN => dout(14));
   U26 : INV_X1 port map( A => n19, ZN => dout(16));
   U27 : INV_X1 port map( A => n20, ZN => dout(17));
   U28 : INV_X1 port map( A => n46, ZN => dout(3));
   U29 : AOI22_X1 port map( A1 => din0(3), A2 => n3, B1 => din1(3), B2 => n6, 
                           ZN => n46);
   U30 : INV_X1 port map( A => n23, ZN => dout(1));
   U31 : AOI22_X1 port map( A1 => din0(1), A2 => n3, B1 => din1(1), B2 => n9, 
                           ZN => n23);
   U32 : INV_X1 port map( A => n51, ZN => dout(8));
   U33 : AOI22_X1 port map( A1 => din0(8), A2 => n3, B1 => din1(8), B2 => n5, 
                           ZN => n51);
   U34 : INV_X1 port map( A => n35, ZN => dout(2));
   U35 : AOI22_X1 port map( A1 => din0(2), A2 => n4, B1 => din1(2), B2 => n6, 
                           ZN => n35);
   U36 : INV_X1 port map( A => n15, ZN => dout(12));
   U37 : AOI22_X1 port map( A1 => din0(12), A2 => n3, B1 => din1(12), B2 => n11
                           , ZN => n15);
   U38 : INV_X1 port map( A => n24, ZN => dout(20));
   U39 : AOI22_X1 port map( A1 => din0(20), A2 => n3, B1 => din1(20), B2 => n9,
                           ZN => n24);
   U40 : INV_X1 port map( A => n49, ZN => dout(6));
   U41 : AOI22_X1 port map( A1 => din0(6), A2 => n3, B1 => din1(6), B2 => n5, 
                           ZN => n49);
   U42 : INV_X1 port map( A => n18, ZN => dout(15));
   U43 : INV_X1 port map( A => n52, ZN => dout(9));
   U44 : AOI22_X1 port map( A1 => din0(9), A2 => n4, B1 => n10, B2 => din1(9), 
                           ZN => n52);
   U45 : INV_X1 port map( A => n47, ZN => dout(4));
   U46 : AOI22_X1 port map( A1 => din0(4), A2 => n4, B1 => din1(4), B2 => n6, 
                           ZN => n47);
   U47 : INV_X1 port map( A => n29, ZN => dout(25));
   U48 : AOI22_X1 port map( A1 => din0(25), A2 => n3, B1 => din1(25), B2 => n8,
                           ZN => n29);
   U49 : INV_X1 port map( A => n33, ZN => dout(29));
   U50 : AOI22_X1 port map( A1 => din0(29), A2 => n4, B1 => din1(29), B2 => n7,
                           ZN => n33);
   U51 : INV_X1 port map( A => n31, ZN => dout(27));
   U52 : AOI22_X1 port map( A1 => din0(27), A2 => n4, B1 => din1(27), B2 => n7,
                           ZN => n31);
   U53 : INV_X1 port map( A => n30, ZN => dout(26));
   U54 : AOI22_X1 port map( A1 => din0(26), A2 => n4, B1 => din1(26), B2 => n7,
                           ZN => n30);
   U55 : INV_X1 port map( A => n45, ZN => dout(31));
   U56 : AOI22_X1 port map( A1 => din0(31), A2 => n3, B1 => din1(31), B2 => n6,
                           ZN => n45);
   U57 : INV_X1 port map( A => n44, ZN => dout(30));
   U58 : AOI22_X1 port map( A1 => din0(30), A2 => n3, B1 => din1(30), B2 => n9,
                           ZN => n44);
   U59 : INV_X1 port map( A => n28, ZN => dout(24));
   U60 : AOI22_X1 port map( A1 => din0(24), A2 => n4, B1 => din1(24), B2 => n8,
                           ZN => n28);
   U61 : INV_X1 port map( A => n27, ZN => dout(23));
   U62 : AOI22_X1 port map( A1 => din0(23), A2 => n3, B1 => din1(23), B2 => n8,
                           ZN => n27);
   U63 : INV_X1 port map( A => n26, ZN => dout(22));
   U64 : AOI22_X1 port map( A1 => din0(22), A2 => n4, B1 => din1(22), B2 => n8,
                           ZN => n26);
   U65 : INV_X1 port map( A => n32, ZN => dout(28));
   U66 : AOI22_X1 port map( A1 => din0(28), A2 => n3, B1 => din1(28), B2 => n7,
                           ZN => n32);
   U67 : AOI22_X1 port map( A1 => din0(19), A2 => n3, B1 => din1(19), B2 => n10
                           , ZN => n22);
   U68 : AOI22_X1 port map( A1 => din0(15), A2 => n4, B1 => din1(15), B2 => n11
                           , ZN => n18);
   U69 : AOI22_X1 port map( A1 => din0(18), A2 => n3, B1 => din1(18), B2 => n10
                           , ZN => n21);
   U70 : AOI22_X1 port map( A1 => din0(16), A2 => n4, B1 => din1(16), B2 => n10
                           , ZN => n19);
   U71 : AOI22_X1 port map( A1 => din0(14), A2 => n4, B1 => din1(14), B2 => n11
                           , ZN => n17);
   U72 : AOI22_X1 port map( A1 => din0(17), A2 => n3, B1 => din1(17), B2 => n10
                           , ZN => n20);
   U73 : INV_X1 port map( A => n12, ZN => dout(0));
   U74 : AOI22_X1 port map( A1 => n2, A2 => din0(0), B1 => sel, B2 => din1(0), 
                           ZN => n12);
   U75 : INV_X1 port map( A => n1, ZN => n4);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Adder_DATA_SIZE32_7 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end Adder_DATA_SIZE32_7;

architecture SYN_adder_arch of Adder_DATA_SIZE32_7 is

   component P4Adder_DATA_SIZE32_SPARSITY4_7
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;

begin
   
   ADDER0 : P4Adder_DATA_SIZE32_SPARSITY4_7 port map( cin => cin, a(31) => 
                           a(31), a(30) => a(30), a(29) => a(29), a(28) => 
                           a(28), a(27) => a(27), a(26) => a(26), a(25) => 
                           a(25), a(24) => a(24), a(23) => a(23), a(22) => 
                           a(22), a(21) => a(21), a(20) => a(20), a(19) => 
                           a(19), a(18) => a(18), a(17) => a(17), a(16) => 
                           a(16), a(15) => a(15), a(14) => a(14), a(13) => 
                           a(13), a(12) => a(12), a(11) => a(11), a(10) => 
                           a(10), a(9) => a(9), a(8) => a(8), a(7) => a(7), 
                           a(6) => a(6), a(5) => a(5), a(4) => a(4), a(3) => 
                           a(3), a(2) => a(2), a(1) => a(1), a(0) => a(0), 
                           b(31) => b(31), b(30) => b(30), b(29) => b(29), 
                           b(28) => b(28), b(27) => b(27), b(26) => b(26), 
                           b(25) => b(25), b(24) => b(24), b(23) => b(23), 
                           b(22) => b(22), b(21) => b(21), b(20) => b(20), 
                           b(19) => b(19), b(18) => b(18), b(17) => b(17), 
                           b(16) => b(16), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           s(31) => s(31), s(30) => s(30), s(29) => s(29), 
                           s(28) => s(28), s(27) => s(27), s(26) => s(26), 
                           s(25) => s(25), s(24) => s(24), s(23) => s(23), 
                           s(22) => s(22), s(21) => s(21), s(20) => s(20), 
                           s(19) => s(19), s(18) => s(18), s(17) => s(17), 
                           s(16) => s(16), s(15) => s(15), s(14) => s(14), 
                           s(13) => s(13), s(12) => s(12), s(11) => s(11), 
                           s(10) => s(10), s(9) => s(9), s(8) => s(8), s(7) => 
                           s(7), s(6) => s(6), s(5) => s(5), s(4) => s(4), s(3)
                           => s(3), s(2) => s(2), s(1) => s(1), s(0) => s(0), 
                           cout => cout);

end SYN_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Adder_DATA_SIZE32_6 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end Adder_DATA_SIZE32_6;

architecture SYN_adder_arch of Adder_DATA_SIZE32_6 is

   component P4Adder_DATA_SIZE32_SPARSITY4_6
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;

begin
   
   ADDER0 : P4Adder_DATA_SIZE32_SPARSITY4_6 port map( cin => cin, a(31) => 
                           a(31), a(30) => a(30), a(29) => a(29), a(28) => 
                           a(28), a(27) => a(27), a(26) => a(26), a(25) => 
                           a(25), a(24) => a(24), a(23) => a(23), a(22) => 
                           a(22), a(21) => a(21), a(20) => a(20), a(19) => 
                           a(19), a(18) => a(18), a(17) => a(17), a(16) => 
                           a(16), a(15) => a(15), a(14) => a(14), a(13) => 
                           a(13), a(12) => a(12), a(11) => a(11), a(10) => 
                           a(10), a(9) => a(9), a(8) => a(8), a(7) => a(7), 
                           a(6) => a(6), a(5) => a(5), a(4) => a(4), a(3) => 
                           a(3), a(2) => a(2), a(1) => a(1), a(0) => a(0), 
                           b(31) => b(31), b(30) => b(30), b(29) => b(29), 
                           b(28) => b(28), b(27) => b(27), b(26) => b(26), 
                           b(25) => b(25), b(24) => b(24), b(23) => b(23), 
                           b(22) => b(22), b(21) => b(21), b(20) => b(20), 
                           b(19) => b(19), b(18) => b(18), b(17) => b(17), 
                           b(16) => b(16), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           s(31) => s(31), s(30) => s(30), s(29) => s(29), 
                           s(28) => s(28), s(27) => s(27), s(26) => s(26), 
                           s(25) => s(25), s(24) => s(24), s(23) => s(23), 
                           s(22) => s(22), s(21) => s(21), s(20) => s(20), 
                           s(19) => s(19), s(18) => s(18), s(17) => s(17), 
                           s(16) => s(16), s(15) => s(15), s(14) => s(14), 
                           s(13) => s(13), s(12) => s(12), s(11) => s(11), 
                           s(10) => s(10), s(9) => s(9), s(8) => s(8), s(7) => 
                           s(7), s(6) => s(6), s(5) => s(5), s(4) => s(4), s(3)
                           => s(3), s(2) => s(2), s(1) => s(1), s(0) => s(0), 
                           cout => cout);

end SYN_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Adder_DATA_SIZE32_5 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end Adder_DATA_SIZE32_5;

architecture SYN_adder_arch of Adder_DATA_SIZE32_5 is

   component P4Adder_DATA_SIZE32_SPARSITY4_5
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;

begin
   
   ADDER0 : P4Adder_DATA_SIZE32_SPARSITY4_5 port map( cin => cin, a(31) => 
                           a(31), a(30) => a(30), a(29) => a(29), a(28) => 
                           a(28), a(27) => a(27), a(26) => a(26), a(25) => 
                           a(25), a(24) => a(24), a(23) => a(23), a(22) => 
                           a(22), a(21) => a(21), a(20) => a(20), a(19) => 
                           a(19), a(18) => a(18), a(17) => a(17), a(16) => 
                           a(16), a(15) => a(15), a(14) => a(14), a(13) => 
                           a(13), a(12) => a(12), a(11) => a(11), a(10) => 
                           a(10), a(9) => a(9), a(8) => a(8), a(7) => a(7), 
                           a(6) => a(6), a(5) => a(5), a(4) => a(4), a(3) => 
                           a(3), a(2) => a(2), a(1) => a(1), a(0) => a(0), 
                           b(31) => b(31), b(30) => b(30), b(29) => b(29), 
                           b(28) => b(28), b(27) => b(27), b(26) => b(26), 
                           b(25) => b(25), b(24) => b(24), b(23) => b(23), 
                           b(22) => b(22), b(21) => b(21), b(20) => b(20), 
                           b(19) => b(19), b(18) => b(18), b(17) => b(17), 
                           b(16) => b(16), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           s(31) => s(31), s(30) => s(30), s(29) => s(29), 
                           s(28) => s(28), s(27) => s(27), s(26) => s(26), 
                           s(25) => s(25), s(24) => s(24), s(23) => s(23), 
                           s(22) => s(22), s(21) => s(21), s(20) => s(20), 
                           s(19) => s(19), s(18) => s(18), s(17) => s(17), 
                           s(16) => s(16), s(15) => s(15), s(14) => s(14), 
                           s(13) => s(13), s(12) => s(12), s(11) => s(11), 
                           s(10) => s(10), s(9) => s(9), s(8) => s(8), s(7) => 
                           s(7), s(6) => s(6), s(5) => s(5), s(4) => s(4), s(3)
                           => s(3), s(2) => s(2), s(1) => s(1), s(0) => s(0), 
                           cout => cout);

end SYN_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Adder_DATA_SIZE32_4 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end Adder_DATA_SIZE32_4;

architecture SYN_adder_arch of Adder_DATA_SIZE32_4 is

   component P4Adder_DATA_SIZE32_SPARSITY4_4
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;

begin
   
   ADDER0 : P4Adder_DATA_SIZE32_SPARSITY4_4 port map( cin => cin, a(31) => 
                           a(31), a(30) => a(30), a(29) => a(29), a(28) => 
                           a(28), a(27) => a(27), a(26) => a(26), a(25) => 
                           a(25), a(24) => a(24), a(23) => a(23), a(22) => 
                           a(22), a(21) => a(21), a(20) => a(20), a(19) => 
                           a(19), a(18) => a(18), a(17) => a(17), a(16) => 
                           a(16), a(15) => a(15), a(14) => a(14), a(13) => 
                           a(13), a(12) => a(12), a(11) => a(11), a(10) => 
                           a(10), a(9) => a(9), a(8) => a(8), a(7) => a(7), 
                           a(6) => a(6), a(5) => a(5), a(4) => a(4), a(3) => 
                           a(3), a(2) => a(2), a(1) => a(1), a(0) => a(0), 
                           b(31) => b(31), b(30) => b(30), b(29) => b(29), 
                           b(28) => b(28), b(27) => b(27), b(26) => b(26), 
                           b(25) => b(25), b(24) => b(24), b(23) => b(23), 
                           b(22) => b(22), b(21) => b(21), b(20) => b(20), 
                           b(19) => b(19), b(18) => b(18), b(17) => b(17), 
                           b(16) => b(16), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           s(31) => s(31), s(30) => s(30), s(29) => s(29), 
                           s(28) => s(28), s(27) => s(27), s(26) => s(26), 
                           s(25) => s(25), s(24) => s(24), s(23) => s(23), 
                           s(22) => s(22), s(21) => s(21), s(20) => s(20), 
                           s(19) => s(19), s(18) => s(18), s(17) => s(17), 
                           s(16) => s(16), s(15) => s(15), s(14) => s(14), 
                           s(13) => s(13), s(12) => s(12), s(11) => s(11), 
                           s(10) => s(10), s(9) => s(9), s(8) => s(8), s(7) => 
                           s(7), s(6) => s(6), s(5) => s(5), s(4) => s(4), s(3)
                           => s(3), s(2) => s(2), s(1) => s(1), s(0) => s(0), 
                           cout => cout);

end SYN_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Adder_DATA_SIZE32_3 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end Adder_DATA_SIZE32_3;

architecture SYN_adder_arch of Adder_DATA_SIZE32_3 is

   component P4Adder_DATA_SIZE32_SPARSITY4_3
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;

begin
   
   ADDER0 : P4Adder_DATA_SIZE32_SPARSITY4_3 port map( cin => cin, a(31) => 
                           a(31), a(30) => a(30), a(29) => a(29), a(28) => 
                           a(28), a(27) => a(27), a(26) => a(26), a(25) => 
                           a(25), a(24) => a(24), a(23) => a(23), a(22) => 
                           a(22), a(21) => a(21), a(20) => a(20), a(19) => 
                           a(19), a(18) => a(18), a(17) => a(17), a(16) => 
                           a(16), a(15) => a(15), a(14) => a(14), a(13) => 
                           a(13), a(12) => a(12), a(11) => a(11), a(10) => 
                           a(10), a(9) => a(9), a(8) => a(8), a(7) => a(7), 
                           a(6) => a(6), a(5) => a(5), a(4) => a(4), a(3) => 
                           a(3), a(2) => a(2), a(1) => a(1), a(0) => a(0), 
                           b(31) => b(31), b(30) => b(30), b(29) => b(29), 
                           b(28) => b(28), b(27) => b(27), b(26) => b(26), 
                           b(25) => b(25), b(24) => b(24), b(23) => b(23), 
                           b(22) => b(22), b(21) => b(21), b(20) => b(20), 
                           b(19) => b(19), b(18) => b(18), b(17) => b(17), 
                           b(16) => b(16), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           s(31) => s(31), s(30) => s(30), s(29) => s(29), 
                           s(28) => s(28), s(27) => s(27), s(26) => s(26), 
                           s(25) => s(25), s(24) => s(24), s(23) => s(23), 
                           s(22) => s(22), s(21) => s(21), s(20) => s(20), 
                           s(19) => s(19), s(18) => s(18), s(17) => s(17), 
                           s(16) => s(16), s(15) => s(15), s(14) => s(14), 
                           s(13) => s(13), s(12) => s(12), s(11) => s(11), 
                           s(10) => s(10), s(9) => s(9), s(8) => s(8), s(7) => 
                           s(7), s(6) => s(6), s(5) => s(5), s(4) => s(4), s(3)
                           => s(3), s(2) => s(2), s(1) => s(1), s(0) => s(0), 
                           cout => cout);

end SYN_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Adder_DATA_SIZE32_2 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end Adder_DATA_SIZE32_2;

architecture SYN_adder_arch of Adder_DATA_SIZE32_2 is

   component P4Adder_DATA_SIZE32_SPARSITY4_2
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;

begin
   
   ADDER0 : P4Adder_DATA_SIZE32_SPARSITY4_2 port map( cin => cin, a(31) => 
                           a(31), a(30) => a(30), a(29) => a(29), a(28) => 
                           a(28), a(27) => a(27), a(26) => a(26), a(25) => 
                           a(25), a(24) => a(24), a(23) => a(23), a(22) => 
                           a(22), a(21) => a(21), a(20) => a(20), a(19) => 
                           a(19), a(18) => a(18), a(17) => a(17), a(16) => 
                           a(16), a(15) => a(15), a(14) => a(14), a(13) => 
                           a(13), a(12) => a(12), a(11) => a(11), a(10) => 
                           a(10), a(9) => a(9), a(8) => a(8), a(7) => a(7), 
                           a(6) => a(6), a(5) => a(5), a(4) => a(4), a(3) => 
                           a(3), a(2) => a(2), a(1) => a(1), a(0) => a(0), 
                           b(31) => b(31), b(30) => b(30), b(29) => b(29), 
                           b(28) => b(28), b(27) => b(27), b(26) => b(26), 
                           b(25) => b(25), b(24) => b(24), b(23) => b(23), 
                           b(22) => b(22), b(21) => b(21), b(20) => b(20), 
                           b(19) => b(19), b(18) => b(18), b(17) => b(17), 
                           b(16) => b(16), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           s(31) => s(31), s(30) => s(30), s(29) => s(29), 
                           s(28) => s(28), s(27) => s(27), s(26) => s(26), 
                           s(25) => s(25), s(24) => s(24), s(23) => s(23), 
                           s(22) => s(22), s(21) => s(21), s(20) => s(20), 
                           s(19) => s(19), s(18) => s(18), s(17) => s(17), 
                           s(16) => s(16), s(15) => s(15), s(14) => s(14), 
                           s(13) => s(13), s(12) => s(12), s(11) => s(11), 
                           s(10) => s(10), s(9) => s(9), s(8) => s(8), s(7) => 
                           s(7), s(6) => s(6), s(5) => s(5), s(4) => s(4), s(3)
                           => s(3), s(2) => s(2), s(1) => s(1), s(0) => s(0), 
                           cout => cout);

end SYN_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Adder_DATA_SIZE32_1 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end Adder_DATA_SIZE32_1;

architecture SYN_adder_arch of Adder_DATA_SIZE32_1 is

   component P4Adder_DATA_SIZE32_SPARSITY4_1
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;

begin
   
   ADDER0 : P4Adder_DATA_SIZE32_SPARSITY4_1 port map( cin => cin, a(31) => 
                           a(31), a(30) => a(30), a(29) => a(29), a(28) => 
                           a(28), a(27) => a(27), a(26) => a(26), a(25) => 
                           a(25), a(24) => a(24), a(23) => a(23), a(22) => 
                           a(22), a(21) => a(21), a(20) => a(20), a(19) => 
                           a(19), a(18) => a(18), a(17) => a(17), a(16) => 
                           a(16), a(15) => a(15), a(14) => a(14), a(13) => 
                           a(13), a(12) => a(12), a(11) => a(11), a(10) => 
                           a(10), a(9) => a(9), a(8) => a(8), a(7) => a(7), 
                           a(6) => a(6), a(5) => a(5), a(4) => a(4), a(3) => 
                           a(3), a(2) => a(2), a(1) => a(1), a(0) => a(0), 
                           b(31) => b(31), b(30) => b(30), b(29) => b(29), 
                           b(28) => b(28), b(27) => b(27), b(26) => b(26), 
                           b(25) => b(25), b(24) => b(24), b(23) => b(23), 
                           b(22) => b(22), b(21) => b(21), b(20) => b(20), 
                           b(19) => b(19), b(18) => b(18), b(17) => b(17), 
                           b(16) => b(16), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           s(31) => s(31), s(30) => s(30), s(29) => s(29), 
                           s(28) => s(28), s(27) => s(27), s(26) => s(26), 
                           s(25) => s(25), s(24) => s(24), s(23) => s(23), 
                           s(22) => s(22), s(21) => s(21), s(20) => s(20), 
                           s(19) => s(19), s(18) => s(18), s(17) => s(17), 
                           s(16) => s(16), s(15) => s(15), s(14) => s(14), 
                           s(13) => s(13), s(12) => s(12), s(11) => s(11), 
                           s(10) => s(10), s(9) => s(9), s(8) => s(8), s(7) => 
                           s(7), s(6) => s(6), s(5) => s(5), s(4) => s(4), s(3)
                           => s(3), s(2) => s(2), s(1) => s(1), s(0) => s(0), 
                           cout => cout);

end SYN_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_0 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_0;

architecture SYN_full_adder_arch of FullAdder_0 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n2, n3 : std_logic;

begin
   
   U3 : XOR2_X1 port map( A => ci, B => n2, Z => s);
   U4 : XOR2_X1 port map( A => a, B => b, Z => n2);
   U1 : INV_X1 port map( A => n3, ZN => co);
   U2 : AOI22_X1 port map( A1 => b, A2 => a, B1 => n2, B2 => ci, ZN => n3);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderSumGenerator_DATA_SIZE64_SPARSITY4 is

   port( a, b : in std_logic_vector (63 downto 0);  cin : in std_logic_vector 
         (15 downto 0);  sum : out std_logic_vector (63 downto 0));

end AdderSumGenerator_DATA_SIZE64_SPARSITY4;

architecture SYN_adder_sum_generator_arch of 
   AdderSumGenerator_DATA_SIZE64_SPARSITY4 is

   component AdderCarrySelect_DATA_SIZE4_17
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_18
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_19
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_20
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_21
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_22
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_23
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_24
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_25
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_26
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_27
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_28
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_29
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_30
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_31
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_32
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;

begin
   
   ACSi_0 : AdderCarrySelect_DATA_SIZE4_32 port map( a(3) => a(3), a(2) => a(2)
                           , a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), sel => cin(0), 
                           sum(3) => sum(3), sum(2) => sum(2), sum(1) => sum(1)
                           , sum(0) => sum(0));
   ACSi_1 : AdderCarrySelect_DATA_SIZE4_31 port map( a(3) => a(7), a(2) => a(6)
                           , a(1) => a(5), a(0) => a(4), b(3) => b(7), b(2) => 
                           b(6), b(1) => b(5), b(0) => b(4), sel => cin(1), 
                           sum(3) => sum(7), sum(2) => sum(6), sum(1) => sum(5)
                           , sum(0) => sum(4));
   ACSi_2 : AdderCarrySelect_DATA_SIZE4_30 port map( a(3) => a(11), a(2) => 
                           a(10), a(1) => a(9), a(0) => a(8), b(3) => b(11), 
                           b(2) => b(10), b(1) => b(9), b(0) => b(8), sel => 
                           cin(2), sum(3) => sum(11), sum(2) => sum(10), sum(1)
                           => sum(9), sum(0) => sum(8));
   ACSi_3 : AdderCarrySelect_DATA_SIZE4_29 port map( a(3) => a(15), a(2) => 
                           a(14), a(1) => a(13), a(0) => a(12), b(3) => b(15), 
                           b(2) => b(14), b(1) => b(13), b(0) => b(12), sel => 
                           cin(3), sum(3) => sum(15), sum(2) => sum(14), sum(1)
                           => sum(13), sum(0) => sum(12));
   ACSi_4 : AdderCarrySelect_DATA_SIZE4_28 port map( a(3) => a(19), a(2) => 
                           a(18), a(1) => a(17), a(0) => a(16), b(3) => b(19), 
                           b(2) => b(18), b(1) => b(17), b(0) => b(16), sel => 
                           cin(4), sum(3) => sum(19), sum(2) => sum(18), sum(1)
                           => sum(17), sum(0) => sum(16));
   ACSi_5 : AdderCarrySelect_DATA_SIZE4_27 port map( a(3) => a(23), a(2) => 
                           a(22), a(1) => a(21), a(0) => a(20), b(3) => b(23), 
                           b(2) => b(22), b(1) => b(21), b(0) => b(20), sel => 
                           cin(5), sum(3) => sum(23), sum(2) => sum(22), sum(1)
                           => sum(21), sum(0) => sum(20));
   ACSi_6 : AdderCarrySelect_DATA_SIZE4_26 port map( a(3) => a(27), a(2) => 
                           a(26), a(1) => a(25), a(0) => a(24), b(3) => b(27), 
                           b(2) => b(26), b(1) => b(25), b(0) => b(24), sel => 
                           cin(6), sum(3) => sum(27), sum(2) => sum(26), sum(1)
                           => sum(25), sum(0) => sum(24));
   ACSi_7 : AdderCarrySelect_DATA_SIZE4_25 port map( a(3) => a(31), a(2) => 
                           a(30), a(1) => a(29), a(0) => a(28), b(3) => b(31), 
                           b(2) => b(30), b(1) => b(29), b(0) => b(28), sel => 
                           cin(7), sum(3) => sum(31), sum(2) => sum(30), sum(1)
                           => sum(29), sum(0) => sum(28));
   ACSi_8 : AdderCarrySelect_DATA_SIZE4_24 port map( a(3) => a(35), a(2) => 
                           a(34), a(1) => a(33), a(0) => a(32), b(3) => b(35), 
                           b(2) => b(34), b(1) => b(33), b(0) => b(32), sel => 
                           cin(8), sum(3) => sum(35), sum(2) => sum(34), sum(1)
                           => sum(33), sum(0) => sum(32));
   ACSi_9 : AdderCarrySelect_DATA_SIZE4_23 port map( a(3) => a(39), a(2) => 
                           a(38), a(1) => a(37), a(0) => a(36), b(3) => b(39), 
                           b(2) => b(38), b(1) => b(37), b(0) => b(36), sel => 
                           cin(9), sum(3) => sum(39), sum(2) => sum(38), sum(1)
                           => sum(37), sum(0) => sum(36));
   ACSi_10 : AdderCarrySelect_DATA_SIZE4_22 port map( a(3) => a(43), a(2) => 
                           a(42), a(1) => a(41), a(0) => a(40), b(3) => b(43), 
                           b(2) => b(42), b(1) => b(41), b(0) => b(40), sel => 
                           cin(10), sum(3) => sum(43), sum(2) => sum(42), 
                           sum(1) => sum(41), sum(0) => sum(40));
   ACSi_11 : AdderCarrySelect_DATA_SIZE4_21 port map( a(3) => a(47), a(2) => 
                           a(46), a(1) => a(45), a(0) => a(44), b(3) => b(47), 
                           b(2) => b(46), b(1) => b(45), b(0) => b(44), sel => 
                           cin(11), sum(3) => sum(47), sum(2) => sum(46), 
                           sum(1) => sum(45), sum(0) => sum(44));
   ACSi_12 : AdderCarrySelect_DATA_SIZE4_20 port map( a(3) => a(51), a(2) => 
                           a(50), a(1) => a(49), a(0) => a(48), b(3) => b(51), 
                           b(2) => b(50), b(1) => b(49), b(0) => b(48), sel => 
                           cin(12), sum(3) => sum(51), sum(2) => sum(50), 
                           sum(1) => sum(49), sum(0) => sum(48));
   ACSi_13 : AdderCarrySelect_DATA_SIZE4_19 port map( a(3) => a(55), a(2) => 
                           a(54), a(1) => a(53), a(0) => a(52), b(3) => b(55), 
                           b(2) => b(54), b(1) => b(53), b(0) => b(52), sel => 
                           cin(13), sum(3) => sum(55), sum(2) => sum(54), 
                           sum(1) => sum(53), sum(0) => sum(52));
   ACSi_14 : AdderCarrySelect_DATA_SIZE4_18 port map( a(3) => a(59), a(2) => 
                           a(58), a(1) => a(57), a(0) => a(56), b(3) => b(59), 
                           b(2) => b(58), b(1) => b(57), b(0) => b(56), sel => 
                           cin(14), sum(3) => sum(59), sum(2) => sum(58), 
                           sum(1) => sum(57), sum(0) => sum(56));
   ACSi_15 : AdderCarrySelect_DATA_SIZE4_17 port map( a(3) => a(63), a(2) => 
                           a(62), a(1) => a(61), a(0) => a(60), b(3) => b(63), 
                           b(2) => b(62), b(1) => b(61), b(0) => b(60), sel => 
                           cin(15), sum(3) => sum(63), sum(2) => sum(62), 
                           sum(1) => sum(61), sum(0) => sum(60));

end SYN_adder_sum_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4CarryGenerator_DATA_SIZE64_SPARSITY4 is

   port( a, b : in std_logic_vector (63 downto 0);  cin : in std_logic;  cout :
         out std_logic_vector (15 downto 0));

end P4CarryGenerator_DATA_SIZE64_SPARSITY4;

architecture SYN_p4_carry_generator_arch of 
   P4CarryGenerator_DATA_SIZE64_SPARSITY4 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal cout_15_port, n458, n459, n460, cout_10_port, cout_9_port, 
      cout_8_port, cout_7_port, n461, n462, n463, cout_2_port, n464, 
      cout_0_port, n77, n78, n79, n80, n81, n82, n83, n84, n85, n151, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n246, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, 
      n228, n229, n230, n244, n245, n247, n248, n249, n250, n251, n252, n253, 
      n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, 
      cout_4_port, n266, n267, n268, n269, cout_3_port, n271, cout_12_port, 
      n273, n274, cout_11_port, cout_13_port, cout_5_port, cout_1_port, 
      cout_6_port, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, 
      n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, 
      n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, 
      n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, 
      n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, 
      n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, 
      n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, 
      n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, 
      n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, 
      n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, 
      n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, 
      n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, 
      n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, 
      n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, 
      n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, cout_14_port,
      n457 : std_logic;

begin
   cout <= ( cout_15_port, cout_14_port, cout_13_port, cout_12_port, 
      cout_11_port, cout_10_port, cout_9_port, cout_8_port, cout_7_port, 
      cout_6_port, cout_5_port, cout_4_port, cout_3_port, cout_2_port, 
      cout_1_port, cout_0_port );
   
   U199 : NAND3_X1 port map( A1 => a(32), A2 => n151, A3 => b(32), ZN => n246);
   U1 : AND2_X1 port map( A1 => a(31), A2 => b(31), ZN => n217);
   U2 : AND2_X1 port map( A1 => n402, A2 => n403, ZN => n218);
   U3 : AND2_X1 port map( A1 => n425, A2 => n426, ZN => n219);
   U4 : AND2_X1 port map( A1 => b(19), A2 => a(19), ZN => n220);
   U5 : AND2_X1 port map( A1 => b(39), A2 => a(39), ZN => n221);
   U6 : AND2_X1 port map( A1 => b(43), A2 => a(43), ZN => n222);
   U7 : AND2_X1 port map( A1 => b(51), A2 => a(51), ZN => n223);
   U8 : AND2_X1 port map( A1 => a(5), A2 => b(5), ZN => n224);
   U9 : AND2_X1 port map( A1 => n316, A2 => n317, ZN => n225);
   U10 : AND2_X1 port map( A1 => n349, A2 => n350, ZN => n226);
   U11 : AND2_X1 port map( A1 => n429, A2 => n430, ZN => n227);
   U12 : AND2_X1 port map( A1 => n436, A2 => n437, ZN => n228);
   U13 : AND2_X1 port map( A1 => a(52), A2 => b(52), ZN => n229);
   U14 : AND2_X1 port map( A1 => a(56), A2 => b(56), ZN => n230);
   U15 : AND2_X1 port map( A1 => n441, A2 => n442, ZN => n244);
   U16 : NAND2_X1 port map( A1 => n388, A2 => n389, ZN => n245);
   U17 : OR2_X1 port map( A1 => n374, A2 => n247, ZN => n390);
   U18 : OR2_X1 port map( A1 => n264, A2 => n245, ZN => n247);
   U19 : CLKBUF_X1 port map( A => n374, Z => n248);
   U20 : CLKBUF_X1 port map( A => n431, Z => n249);
   U21 : CLKBUF_X1 port map( A => n414, Z => n250);
   U22 : NAND2_X1 port map( A1 => n390, A2 => n254, ZN => n251);
   U23 : NAND2_X1 port map( A1 => n251, A2 => n252, ZN => n267);
   U24 : OR2_X1 port map( A1 => n253, A2 => n218, ZN => n252);
   U25 : INV_X1 port map( A => n405, ZN => n253);
   U26 : AND2_X1 port map( A1 => n391, A2 => n405, ZN => n254);
   U27 : NAND2_X1 port map( A1 => n431, A2 => n258, ZN => n255);
   U28 : AND2_X1 port map( A1 => n255, A2 => n256, ZN => n458);
   U29 : OR2_X1 port map( A1 => n257, A2 => n228, ZN => n256);
   U30 : INV_X1 port map( A => n439, ZN => n257);
   U31 : AND2_X1 port map( A1 => n227, A2 => n439, ZN => n258);
   U32 : NAND2_X1 port map( A1 => n414, A2 => n262, ZN => n259);
   U33 : AND2_X1 port map( A1 => n259, A2 => n260, ZN => n459);
   U34 : OR2_X1 port map( A1 => n261, A2 => n219, ZN => n260);
   U35 : INV_X1 port map( A => n428, ZN => n261);
   U36 : AND2_X1 port map( A1 => n413, A2 => n428, ZN => n262);
   U37 : NAND2_X1 port map( A1 => n318, A2 => n225, ZN => n323);
   U38 : NAND2_X1 port map( A1 => cout_9_port, A2 => n218, ZN => n404);
   U39 : OR2_X1 port map( A1 => n248, A2 => n264, ZN => n263);
   U40 : OR3_X1 port map( A1 => n377, A2 => n376, A3 => n375, ZN => n264);
   U41 : CLKBUF_X1 port map( A => n462, Z => cout_4_port);
   U42 : NAND2_X1 port map( A1 => n348, A2 => n347, ZN => n462);
   U43 : NAND2_X1 port map( A1 => n351, A2 => n226, ZN => n356);
   U44 : CLKBUF_X1 port map( A => n280, Z => n266);
   U45 : NAND2_X1 port map( A1 => n438, A2 => n228, ZN => n440);
   U46 : NAND2_X1 port map( A1 => n460, A2 => n219, ZN => n427);
   U47 : NAND2_X1 port map( A1 => n249, A2 => n227, ZN => n438);
   U48 : NAND2_X1 port map( A1 => n443, A2 => n244, ZN => n448);
   U49 : OR2_X1 port map( A1 => n369, A2 => n368, ZN => n268);
   U50 : NAND2_X1 port map( A1 => n268, A2 => n367, ZN => n457);
   U51 : AND2_X1 port map( A1 => b(11), A2 => a(11), ZN => n269);
   U52 : NOR2_X1 port map( A1 => n269, A2 => n281, ZN => n280);
   U53 : CLKBUF_X1 port map( A => n463, Z => cout_3_port);
   U54 : OR2_X1 port map( A1 => n315, A2 => n314, ZN => n271);
   U55 : NAND2_X1 port map( A1 => n271, A2 => n313, ZN => n464);
   U56 : NAND2_X1 port map( A1 => n428, A2 => n427, ZN => cout_12_port);
   U57 : INV_X1 port map( A => n248, ZN => cout_7_port);
   U58 : NAND2_X1 port map( A1 => n334, A2 => n333, ZN => n463);
   U59 : CLKBUF_X1 port map( A => cout_14_port, Z => n273);
   U60 : CLKBUF_X1 port map( A => n304, Z => n274);
   U61 : NAND2_X1 port map( A1 => n250, A2 => n413, ZN => cout_11_port);
   U62 : NAND2_X1 port map( A1 => n440, A2 => n439, ZN => cout_13_port);
   U63 : CLKBUF_X1 port map( A => n461, Z => cout_5_port);
   U64 : NAND2_X1 port map( A1 => n250, A2 => n413, ZN => n460);
   U65 : INV_X1 port map( A => n266, ZN => cout_2_port);
   U66 : CLKBUF_X1 port map( A => n464, Z => cout_1_port);
   U67 : CLKBUF_X1 port map( A => n457, Z => cout_6_port);
   U68 : AND3_X1 port map( A1 => n323, A2 => n322, A3 => n321, ZN => n281);
   U69 : NAND2_X1 port map( A1 => n454, A2 => n455, ZN => n151);
   U70 : NAND2_X1 port map( A1 => n391, A2 => n390, ZN => cout_9_port);
   U71 : INV_X1 port map( A => a(34), ZN => n240);
   U72 : AND2_X1 port map( A1 => n392, A2 => n393, ZN => n282);
   U73 : AND2_X1 port map( A1 => n415, A2 => n416, ZN => n283);
   U74 : NAND2_X1 port map( A1 => n381, A2 => n382, ZN => n389);
   U75 : AND2_X1 port map( A1 => n335, A2 => n336, ZN => n284);
   U76 : INV_X1 port map( A => n243, ZN => n241);
   U77 : INV_X1 port map( A => n231, ZN => n233);
   U78 : OAI21_X1 port map( B1 => n78, B2 => n79, A => n80, ZN => cout_15_port)
                           ;
   U79 : AND2_X1 port map( A1 => a(28), A2 => b(28), ZN => n285);
   U80 : AOI21_X1 port map( B1 => n233, B2 => a(37), A => b(37), ZN => n232);
   U81 : AOI21_X1 port map( B1 => n234, B2 => a(36), A => n235, ZN => n231);
   U82 : INV_X1 port map( A => n236, ZN => n235);
   U83 : OAI21_X1 port map( B1 => a(36), B2 => n234, A => b(36), ZN => n236);
   U84 : INV_X1 port map( A => n77, ZN => n234);
   U85 : AOI21_X1 port map( B1 => n237, B2 => a(35), A => n238, ZN => n77);
   U86 : INV_X1 port map( A => n239, ZN => n238);
   U87 : OAI21_X1 port map( B1 => n237, B2 => a(35), A => b(35), ZN => n239);
   U88 : AOI21_X1 port map( B1 => n240, B2 => n241, A => n242, ZN => n237);
   U89 : OAI21_X1 port map( B1 => n454, B2 => n455, A => n246, ZN => n243);
   U90 : AOI21_X1 port map( B1 => n243, B2 => a(34), A => b(34), ZN => n242);
   U91 : AND2_X1 port map( A1 => a(3), A2 => b(3), ZN => n286);
   U92 : NAND2_X1 port map( A1 => n358, A2 => n357, ZN => n461);
   U93 : OR2_X1 port map( A1 => b(39), A2 => a(39), ZN => n385);
   U94 : OR2_X1 port map( A1 => b(43), A2 => a(43), ZN => n403);
   U95 : OR2_X1 port map( A1 => b(51), A2 => a(51), ZN => n426);
   U96 : AND2_X1 port map( A1 => n359, A2 => n360, ZN => n287);
   U97 : OR2_X1 port map( A1 => b(18), A2 => a(18), ZN => n342);
   U98 : OR2_X1 port map( A1 => b(42), A2 => a(42), ZN => n399);
   U99 : OR2_X1 port map( A1 => b(50), A2 => a(50), ZN => n422);
   U100 : OR2_X1 port map( A1 => b(19), A2 => a(19), ZN => n346);
   U101 : OR2_X1 port map( A1 => a(22), A2 => b(22), ZN => n355);
   U102 : AND2_X1 port map( A1 => a(24), A2 => b(24), ZN => n288);
   U103 : AND2_X1 port map( A1 => a(20), A2 => b(20), ZN => n289);
   U104 : AND2_X1 port map( A1 => a(8), A2 => b(8), ZN => n290);
   U105 : OAI22_X1 port map( A1 => a(62), A2 => n82, B1 => b(62), B2 => n83, ZN
                           => n78);
   U106 : AND2_X1 port map( A1 => n82, A2 => a(62), ZN => n83);
   U107 : OAI22_X1 port map( A1 => n453, A2 => n452, B1 => n84, B2 => n85, ZN 
                           => n82);
   U108 : INV_X1 port map( A => a(61), ZN => n84);
   U109 : OAI22_X1 port map( A1 => b(60), A2 => a(60), B1 => b(61), B2 => a(61)
                           , ZN => n452);
   U110 : INV_X1 port map( A => b(61), ZN => n85);
   U111 : OAI21_X1 port map( B1 => n81, B2 => a(63), A => b(63), ZN => n80);
   U112 : INV_X1 port map( A => n78, ZN => n81);
   U113 : INV_X1 port map( A => a(63), ZN => n79);
   U114 : NAND2_X1 port map( A1 => n405, A2 => n404, ZN => cout_10_port);
   U115 : NAND2_X1 port map( A1 => n361, A2 => n287, ZN => n366);
   U116 : OR2_X1 port map( A1 => n451, A2 => n450, ZN => n291);
   U117 : NAND2_X1 port map( A1 => n291, A2 => n449, ZN => cout_14_port);
   U118 : OAI22_X1 port map( A1 => n301, A2 => n286, B1 => b(3), B2 => a(3), ZN
                           => n304);
   U119 : AOI21_X1 port map( B1 => a(60), B2 => b(60), A => n273, ZN => n453);
   U120 : OAI22_X1 port map( A1 => n373, A2 => n217, B1 => b(31), B2 => a(31), 
                           ZN => n374);
   U121 : NOR2_X1 port map( A1 => b(0), A2 => a(0), ZN => n293);
   U122 : AOI21_X1 port map( B1 => b(0), B2 => a(0), A => cin, ZN => n292);
   U123 : INV_X1 port map( A => b(1), ZN => n294);
   U124 : INV_X1 port map( A => a(1), ZN => n295);
   U125 : OAI22_X1 port map( A1 => n292, A2 => n293, B1 => n294, B2 => n295, ZN
                           => n297);
   U126 : NAND2_X1 port map( A1 => n295, A2 => n294, ZN => n296);
   U127 : NAND2_X1 port map( A1 => n297, A2 => n296, ZN => n300);
   U128 : NAND2_X1 port map( A1 => a(2), A2 => b(2), ZN => n299);
   U129 : NOR2_X1 port map( A1 => b(2), A2 => a(2), ZN => n298);
   U130 : AOI21_X1 port map( B1 => n300, B2 => n299, A => n298, ZN => n301);
   U131 : INV_X1 port map( A => n274, ZN => cout_0_port);
   U132 : INV_X1 port map( A => b(7), ZN => n315);
   U133 : INV_X1 port map( A => a(7), ZN => n314);
   U134 : NAND2_X1 port map( A1 => a(4), A2 => b(4), ZN => n303);
   U135 : NOR2_X1 port map( A1 => b(4), A2 => a(4), ZN => n302);
   U136 : AOI21_X1 port map( B1 => n304, B2 => n303, A => n302, ZN => n305);
   U137 : OAI22_X1 port map( A1 => n305, A2 => n224, B1 => b(5), B2 => a(5), ZN
                           => n307);
   U138 : NAND2_X1 port map( A1 => a(6), A2 => b(6), ZN => n306);
   U139 : NAND2_X1 port map( A1 => n307, A2 => n306, ZN => n312);
   U140 : INV_X1 port map( A => a(6), ZN => n309);
   U141 : INV_X1 port map( A => b(6), ZN => n308);
   U142 : NAND2_X1 port map( A1 => n309, A2 => n308, ZN => n311);
   U143 : NAND2_X1 port map( A1 => n314, A2 => n315, ZN => n310);
   U144 : NAND3_X1 port map( A1 => n312, A2 => n311, A3 => n310, ZN => n313);
   U145 : INV_X1 port map( A => b(11), ZN => n325);
   U146 : INV_X1 port map( A => a(11), ZN => n324);
   U147 : OAI222_X1 port map( A1 => n464, A2 => n290, B1 => b(8), B2 => a(8), 
                           C1 => b(9), C2 => a(9), ZN => n318);
   U148 : NAND2_X1 port map( A1 => a(10), A2 => b(10), ZN => n317);
   U149 : NAND2_X1 port map( A1 => a(9), A2 => b(9), ZN => n316);
   U150 : INV_X1 port map( A => a(10), ZN => n320);
   U151 : INV_X1 port map( A => b(10), ZN => n319);
   U152 : NAND2_X1 port map( A1 => n320, A2 => n319, ZN => n322);
   U153 : NAND2_X1 port map( A1 => n324, A2 => n325, ZN => n321);
   U154 : NAND2_X1 port map( A1 => a(12), A2 => b(12), ZN => n328);
   U155 : NOR2_X1 port map( A1 => b(13), A2 => a(13), ZN => n327);
   U156 : NOR2_X1 port map( A1 => b(12), A2 => a(12), ZN => n326);
   U157 : AOI211_X1 port map( C1 => n280, C2 => n328, A => n327, B => n326, ZN 
                           => n332);
   U158 : NAND2_X1 port map( A1 => a(13), A2 => b(13), ZN => n330);
   U159 : NAND2_X1 port map( A1 => a(14), A2 => b(14), ZN => n329);
   U160 : NAND2_X1 port map( A1 => n330, A2 => n329, ZN => n331);
   U161 : OAI222_X1 port map( A1 => n332, A2 => n331, B1 => a(15), B2 => b(15),
                           C1 => b(14), C2 => a(14), ZN => n334);
   U162 : NAND2_X1 port map( A1 => b(15), A2 => a(15), ZN => n333);
   U163 : INV_X1 port map( A => b(17), ZN => n335);
   U164 : INV_X1 port map( A => a(17), ZN => n336);
   U165 : NAND2_X1 port map( A1 => a(16), A2 => b(16), ZN => n337);
   U166 : OAI22_X1 port map( A1 => n284, A2 => n337, B1 => n336, B2 => n335, ZN
                           => n338);
   U167 : NAND2_X1 port map( A1 => n338, A2 => n342, ZN => n340);
   U168 : NAND2_X1 port map( A1 => b(18), A2 => a(18), ZN => n339);
   U169 : NAND2_X1 port map( A1 => n340, A2 => n339, ZN => n341);
   U170 : AOI21_X1 port map( B1 => n341, B2 => n346, A => n220, ZN => n348);
   U171 : INV_X1 port map( A => n342, ZN => n344);
   U172 : NOR2_X1 port map( A1 => b(16), A2 => a(16), ZN => n343);
   U173 : NOR3_X1 port map( A1 => n344, A2 => n343, A3 => n284, ZN => n345);
   U174 : NAND3_X1 port map( A1 => n463, A2 => n346, A3 => n345, ZN => n347);
   U175 : OAI222_X1 port map( A1 => n462, A2 => n289, B1 => b(20), B2 => a(20),
                           C1 => b(21), C2 => a(21), ZN => n351);
   U176 : NAND2_X1 port map( A1 => a(22), A2 => b(22), ZN => n350);
   U177 : NAND2_X1 port map( A1 => a(21), A2 => b(21), ZN => n349);
   U178 : INV_X1 port map( A => b(23), ZN => n353);
   U179 : INV_X1 port map( A => a(23), ZN => n352);
   U180 : NAND2_X1 port map( A1 => n353, A2 => n352, ZN => n354);
   U181 : NAND3_X1 port map( A1 => n356, A2 => n355, A3 => n354, ZN => n358);
   U182 : NAND2_X1 port map( A1 => b(23), A2 => a(23), ZN => n357);
   U183 : INV_X1 port map( A => b(27), ZN => n369);
   U184 : INV_X1 port map( A => a(27), ZN => n368);
   U185 : OAI222_X1 port map( A1 => n461, A2 => n288, B1 => b(24), B2 => a(24),
                           C1 => b(25), C2 => a(25), ZN => n361);
   U186 : NAND2_X1 port map( A1 => a(26), A2 => b(26), ZN => n360);
   U187 : NAND2_X1 port map( A1 => a(25), A2 => b(25), ZN => n359);
   U188 : INV_X1 port map( A => a(26), ZN => n363);
   U189 : INV_X1 port map( A => b(26), ZN => n362);
   U190 : NAND2_X1 port map( A1 => n363, A2 => n362, ZN => n365);
   U191 : NAND2_X1 port map( A1 => n368, A2 => n369, ZN => n364);
   U192 : NAND3_X1 port map( A1 => n366, A2 => n365, A3 => n364, ZN => n367);
   U193 : AOI22_X1 port map( A1 => a(30), A2 => b(30), B1 => a(29), B2 => b(29)
                           , ZN => n372);
   U194 : OAI222_X1 port map( A1 => n457, A2 => n285, B1 => b(28), B2 => a(28),
                           C1 => b(29), C2 => a(29), ZN => n371);
   U195 : NOR2_X1 port map( A1 => b(30), A2 => a(30), ZN => n370);
   U196 : AOI21_X1 port map( B1 => n371, B2 => n372, A => n370, ZN => n373);
   U197 : INV_X1 port map( A => a(33), ZN => n454);
   U198 : INV_X1 port map( A => b(33), ZN => n455);
   U200 : OAI22_X1 port map( A1 => b(32), A2 => a(32), B1 => b(34), B2 => a(34)
                           , ZN => n377);
   U201 : NOR2_X1 port map( A1 => b(35), A2 => a(35), ZN => n376);
   U202 : INV_X1 port map( A => n151, ZN => n375);
   U203 : NAND2_X1 port map( A1 => n77, A2 => n263, ZN => cout_8_port);
   U204 : INV_X1 port map( A => a(37), ZN => n379);
   U205 : INV_X1 port map( A => b(38), ZN => n381);
   U206 : INV_X1 port map( A => a(38), ZN => n382);
   U207 : INV_X1 port map( A => n389, ZN => n378);
   U208 : AOI21_X1 port map( B1 => n231, B2 => n379, A => n378, ZN => n380);
   U209 : INV_X1 port map( A => n380, ZN => n383);
   U210 : OAI22_X1 port map( A1 => n383, A2 => n232, B1 => n382, B2 => n381, ZN
                           => n384);
   U211 : AOI21_X1 port map( B1 => n384, B2 => n385, A => n221, ZN => n391);
   U212 : OAI22_X1 port map( A1 => b(36), A2 => a(36), B1 => a(37), B2 => b(37)
                           , ZN => n387);
   U213 : INV_X1 port map( A => n385, ZN => n386);
   U214 : NOR2_X1 port map( A1 => n387, A2 => n386, ZN => n388);
   U215 : INV_X1 port map( A => b(41), ZN => n392);
   U216 : INV_X1 port map( A => a(41), ZN => n393);
   U217 : NAND2_X1 port map( A1 => a(40), A2 => b(40), ZN => n394);
   U218 : OAI22_X1 port map( A1 => n282, A2 => n394, B1 => n393, B2 => n392, ZN
                           => n395);
   U219 : NAND2_X1 port map( A1 => n395, A2 => n399, ZN => n397);
   U220 : NAND2_X1 port map( A1 => b(42), A2 => a(42), ZN => n396);
   U221 : NAND2_X1 port map( A1 => n397, A2 => n396, ZN => n398);
   U222 : AOI21_X1 port map( B1 => n398, B2 => n403, A => n222, ZN => n405);
   U223 : INV_X1 port map( A => n399, ZN => n401);
   U224 : NOR2_X1 port map( A1 => b(40), A2 => a(40), ZN => n400);
   U225 : NOR3_X1 port map( A1 => n401, A2 => n400, A3 => n282, ZN => n402);
   U226 : NAND2_X1 port map( A1 => a(44), A2 => b(44), ZN => n408);
   U227 : NOR2_X1 port map( A1 => b(45), A2 => a(45), ZN => n407);
   U228 : NOR2_X1 port map( A1 => b(44), A2 => a(44), ZN => n406);
   U229 : AOI211_X1 port map( C1 => n267, C2 => n408, A => n407, B => n406, ZN 
                           => n412);
   U230 : NAND2_X1 port map( A1 => a(45), A2 => b(45), ZN => n410);
   U231 : NAND2_X1 port map( A1 => a(46), A2 => b(46), ZN => n409);
   U232 : NAND2_X1 port map( A1 => n410, A2 => n409, ZN => n411);
   U233 : OAI222_X1 port map( A1 => n412, A2 => n411, B1 => a(47), B2 => b(47),
                           C1 => b(46), C2 => a(46), ZN => n414);
   U234 : NAND2_X1 port map( A1 => b(47), A2 => a(47), ZN => n413);
   U235 : INV_X1 port map( A => b(49), ZN => n415);
   U236 : INV_X1 port map( A => a(49), ZN => n416);
   U237 : NAND2_X1 port map( A1 => a(48), A2 => b(48), ZN => n417);
   U238 : OAI22_X1 port map( A1 => n283, A2 => n417, B1 => n416, B2 => n415, ZN
                           => n418);
   U239 : NAND2_X1 port map( A1 => n418, A2 => n422, ZN => n420);
   U240 : NAND2_X1 port map( A1 => b(50), A2 => a(50), ZN => n419);
   U241 : NAND2_X1 port map( A1 => n420, A2 => n419, ZN => n421);
   U242 : AOI21_X1 port map( B1 => n421, B2 => n426, A => n223, ZN => n428);
   U243 : INV_X1 port map( A => n422, ZN => n424);
   U244 : NOR2_X1 port map( A1 => b(48), A2 => a(48), ZN => n423);
   U245 : NOR3_X1 port map( A1 => n424, A2 => n423, A3 => n283, ZN => n425);
   U246 : OAI222_X1 port map( A1 => n459, A2 => n229, B1 => b(52), B2 => a(52),
                           C1 => b(53), C2 => a(53), ZN => n431);
   U247 : NAND2_X1 port map( A1 => a(54), A2 => b(54), ZN => n430);
   U248 : NAND2_X1 port map( A1 => a(53), A2 => b(53), ZN => n429);
   U249 : INV_X1 port map( A => a(54), ZN => n433);
   U250 : INV_X1 port map( A => b(54), ZN => n432);
   U251 : NAND2_X1 port map( A1 => n433, A2 => n432, ZN => n437);
   U252 : INV_X1 port map( A => b(55), ZN => n435);
   U253 : INV_X1 port map( A => a(55), ZN => n434);
   U254 : NAND2_X1 port map( A1 => n435, A2 => n434, ZN => n436);
   U255 : NAND2_X1 port map( A1 => b(55), A2 => a(55), ZN => n439);
   U256 : INV_X1 port map( A => b(59), ZN => n451);
   U257 : INV_X1 port map( A => a(59), ZN => n450);
   U258 : OAI222_X1 port map( A1 => n230, A2 => n458, B1 => b(56), B2 => a(56),
                           C1 => b(57), C2 => a(57), ZN => n443);
   U259 : NAND2_X1 port map( A1 => a(58), A2 => b(58), ZN => n442);
   U260 : NAND2_X1 port map( A1 => a(57), A2 => b(57), ZN => n441);
   U261 : INV_X1 port map( A => a(58), ZN => n445);
   U262 : INV_X1 port map( A => b(58), ZN => n444);
   U263 : NAND2_X1 port map( A1 => n445, A2 => n444, ZN => n447);
   U264 : NAND2_X1 port map( A1 => n450, A2 => n451, ZN => n446);
   U265 : NAND3_X1 port map( A1 => n448, A2 => n447, A3 => n446, ZN => n449);

end SYN_p4_carry_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderSumGenerator_DATA_SIZE16_SPARSITY4 is

   port( a, b : in std_logic_vector (15 downto 0);  cin : in std_logic_vector 
         (3 downto 0);  sum : out std_logic_vector (15 downto 0));

end AdderSumGenerator_DATA_SIZE16_SPARSITY4;

architecture SYN_adder_sum_generator_arch of 
   AdderSumGenerator_DATA_SIZE16_SPARSITY4 is

   component AdderCarrySelect_DATA_SIZE4_57
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_58
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_59
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_60
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;

begin
   
   ACSi_0 : AdderCarrySelect_DATA_SIZE4_60 port map( a(3) => a(3), a(2) => a(2)
                           , a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), sel => cin(0), 
                           sum(3) => sum(3), sum(2) => sum(2), sum(1) => sum(1)
                           , sum(0) => sum(0));
   ACSi_1 : AdderCarrySelect_DATA_SIZE4_59 port map( a(3) => a(7), a(2) => a(6)
                           , a(1) => a(5), a(0) => a(4), b(3) => b(7), b(2) => 
                           b(6), b(1) => b(5), b(0) => b(4), sel => cin(1), 
                           sum(3) => sum(7), sum(2) => sum(6), sum(1) => sum(5)
                           , sum(0) => sum(4));
   ACSi_2 : AdderCarrySelect_DATA_SIZE4_58 port map( a(3) => a(11), a(2) => 
                           a(10), a(1) => a(9), a(0) => a(8), b(3) => b(11), 
                           b(2) => b(10), b(1) => b(9), b(0) => b(8), sel => 
                           cin(2), sum(3) => sum(11), sum(2) => sum(10), sum(1)
                           => sum(9), sum(0) => sum(8));
   ACSi_3 : AdderCarrySelect_DATA_SIZE4_57 port map( a(3) => a(15), a(2) => 
                           a(14), a(1) => a(13), a(0) => a(12), b(3) => b(15), 
                           b(2) => b(14), b(1) => b(13), b(0) => b(12), sel => 
                           cin(3), sum(3) => sum(15), sum(2) => sum(14), sum(1)
                           => sum(13), sum(0) => sum(12));

end SYN_adder_sum_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4CarryGenerator_DATA_SIZE16_SPARSITY4 is

   port( a, b : in std_logic_vector (15 downto 0);  cin : in std_logic;  cout :
         out std_logic_vector (3 downto 0));

end P4CarryGenerator_DATA_SIZE16_SPARSITY4;

architecture SYN_p4_carry_generator_arch of 
   P4CarryGenerator_DATA_SIZE16_SPARSITY4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal cout_3_port, cout_2_port, cout_1_port, cout_0_port, n19, n21, n22, 
      n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n36, n37, n38
      , n39, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, 
      n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65 : std_logic;

begin
   cout <= ( cout_3_port, cout_2_port, cout_1_port, cout_0_port );
   
   U1 : OAI22_X1 port map( A1 => n33, A2 => n34, B1 => n64, B2 => n36, ZN => 
                           n32);
   U2 : INV_X1 port map( A => b(10), ZN => n36);
   U3 : NOR2_X1 port map( A1 => b(10), A2 => a(10), ZN => n34);
   U4 : AOI21_X1 port map( B1 => b(9), B2 => a(9), A => n37, ZN => n33);
   U5 : INV_X1 port map( A => n27, ZN => n26);
   U6 : OAI222_X1 port map( A1 => a(12), A2 => cout_2_port, B1 => b(12), B2 => 
                           n28, C1 => b(13), C2 => a(13), ZN => n27);
   U7 : AND2_X1 port map( A1 => cout_2_port, A2 => a(12), ZN => n28);
   U8 : OAI22_X1 port map( A1 => a(14), A2 => n23, B1 => b(14), B2 => n24, ZN 
                           => n19);
   U9 : AND2_X1 port map( A1 => n23, A2 => a(14), ZN => n24);
   U10 : INV_X1 port map( A => n25, ZN => n23);
   U11 : AOI21_X1 port map( B1 => a(13), B2 => b(13), A => n26, ZN => n25);
   U12 : INV_X1 port map( A => n42, ZN => cout_1_port);
   U13 : AOI21_X1 port map( B1 => a(7), B2 => b(7), A => n43, ZN => n42);
   U14 : INV_X1 port map( A => n44, ZN => n43);
   U15 : OAI222_X1 port map( A1 => a(6), A2 => n45, B1 => b(6), B2 => n46, C1 
                           => b(7), C2 => a(7), ZN => n44);
   U16 : INV_X1 port map( A => n52, ZN => cout_0_port);
   U17 : OAI22_X1 port map( A1 => a(3), A2 => n53, B1 => b(3), B2 => n54, ZN =>
                           n52);
   U18 : AND2_X1 port map( A1 => n53, A2 => a(3), ZN => n54);
   U19 : INV_X1 port map( A => n55, ZN => n53);
   U20 : OAI22_X1 port map( A1 => a(4), A2 => cout_0_port, B1 => b(4), B2 => 
                           n51, ZN => n50);
   U21 : AND2_X1 port map( A1 => cout_0_port, A2 => a(4), ZN => n51);
   U22 : INV_X1 port map( A => n29, ZN => cout_2_port);
   U23 : AOI21_X1 port map( B1 => a(11), B2 => b(11), A => n30, ZN => n29);
   U24 : INV_X1 port map( A => n31, ZN => n30);
   U25 : OAI21_X1 port map( B1 => a(11), B2 => b(11), A => n32, ZN => n31);
   U26 : OAI22_X1 port map( A1 => a(2), A2 => n56, B1 => b(2), B2 => n57, ZN =>
                           n55);
   U27 : AND2_X1 port map( A1 => n56, A2 => a(2), ZN => n57);
   U28 : INV_X1 port map( A => n58, ZN => n56);
   U29 : OAI22_X1 port map( A1 => a(1), A2 => n59, B1 => b(1), B2 => n60, ZN =>
                           n58);
   U30 : OAI21_X1 port map( B1 => n19, B2 => n65, A => n21, ZN => cout_3_port);
   U31 : AOI22_X1 port map( A1 => n38, A2 => n39, B1 => n63, B2 => n41, ZN => 
                           n37);
   U32 : INV_X1 port map( A => b(9), ZN => n41);
   U33 : NAND2_X1 port map( A1 => a(8), A2 => cout_1_port, ZN => n38);
   U34 : OAI21_X1 port map( B1 => a(8), B2 => cout_1_port, A => b(8), ZN => n39
                           );
   U35 : OAI21_X1 port map( B1 => n22, B2 => a(15), A => b(15), ZN => n21);
   U36 : INV_X1 port map( A => n19, ZN => n22);
   U37 : INV_X1 port map( A => n61, ZN => n59);
   U38 : OAI22_X1 port map( A1 => b(0), A2 => a(0), B1 => cin, B2 => n62, ZN =>
                           n61);
   U39 : AND2_X1 port map( A1 => a(0), A2 => b(0), ZN => n62);
   U40 : INV_X1 port map( A => n47, ZN => n45);
   U41 : OAI22_X1 port map( A1 => a(5), A2 => n48, B1 => b(5), B2 => n49, ZN =>
                           n47);
   U42 : AND2_X1 port map( A1 => n48, A2 => a(5), ZN => n49);
   U43 : INV_X1 port map( A => n50, ZN => n48);
   U44 : AND2_X1 port map( A1 => n59, A2 => a(1), ZN => n60);
   U45 : AND2_X1 port map( A1 => n45, A2 => a(6), ZN => n46);
   U46 : INV_X1 port map( A => a(9), ZN => n63);
   U47 : INV_X1 port map( A => a(10), ZN => n64);
   U48 : INV_X1 port map( A => a(15), ZN => n65);

end SYN_p4_carry_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_0 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_0;

architecture SYN_mux_arch of Mux_DATA_SIZE4_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n6, n7, n8, n9, n10 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n9, ZN => dout(1));
   U2 : AOI22_X1 port map( A1 => din0(1), A2 => n7, B1 => din1(1), B2 => sel, 
                           ZN => n9);
   U3 : INV_X1 port map( A => n10, ZN => dout(0));
   U4 : AOI22_X1 port map( A1 => din0(0), A2 => n7, B1 => din1(0), B2 => sel, 
                           ZN => n10);
   U5 : INV_X1 port map( A => n8, ZN => dout(2));
   U6 : AOI22_X1 port map( A1 => din0(2), A2 => n7, B1 => din1(2), B2 => sel, 
                           ZN => n8);
   U7 : INV_X1 port map( A => n6, ZN => dout(3));
   U8 : AOI22_X1 port map( A1 => din0(3), A2 => n7, B1 => sel, B2 => din1(3), 
                           ZN => n6);
   U9 : INV_X1 port map( A => sel, ZN => n7);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_0 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_0;

architecture SYN_rca_arch of Rca_DATA_SIZE4_0 is

   component FullAdder_669
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_670
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_671
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_0
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_0 port map( ci => ci, a => a(0), b => b(0), s => s(0), co 
                           => carry_1_port);
   FA3_1 : FullAdder_671 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_670 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_669 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4Adder_DATA_SIZE64_SPARSITY4 is

   port( cin : in std_logic;  a, b : in std_logic_vector (63 downto 0);  s : 
         out std_logic_vector (63 downto 0);  cout : out std_logic);

end P4Adder_DATA_SIZE64_SPARSITY4;

architecture SYN_p4_adder_arch of P4Adder_DATA_SIZE64_SPARSITY4 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AdderSumGenerator_DATA_SIZE64_SPARSITY4
      port( a, b : in std_logic_vector (63 downto 0);  cin : in 
            std_logic_vector (15 downto 0);  sum : out std_logic_vector (63 
            downto 0));
   end component;
   
   component P4CarryGenerator_DATA_SIZE64_SPARSITY4
      port( a, b : in std_logic_vector (63 downto 0);  cin : in std_logic;  
            cout : out std_logic_vector (15 downto 0));
   end component;
   
   signal carry_15_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port, 
      carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port, 
      carry_1_port, n1, n2, n3, n4, n5 : std_logic;

begin
   
   CG0 : P4CarryGenerator_DATA_SIZE64_SPARSITY4 port map( a(63) => a(63), a(62)
                           => a(62), a(61) => a(61), a(60) => a(60), a(59) => 
                           a(59), a(58) => a(58), a(57) => a(57), a(56) => 
                           a(56), a(55) => a(55), a(54) => a(54), a(53) => 
                           a(53), a(52) => a(52), a(51) => a(51), a(50) => 
                           a(50), a(49) => a(49), a(48) => a(48), a(47) => 
                           a(47), a(46) => a(46), a(45) => a(45), a(44) => 
                           a(44), a(43) => a(43), a(42) => a(42), a(41) => 
                           a(41), a(40) => a(40), a(39) => a(39), a(38) => 
                           a(38), a(37) => a(37), a(36) => a(36), a(35) => 
                           a(35), a(34) => a(34), a(33) => a(33), a(32) => 
                           a(32), a(31) => a(31), a(30) => a(30), a(29) => 
                           a(29), a(28) => a(28), a(27) => a(27), a(26) => 
                           a(26), a(25) => a(25), a(24) => a(24), a(23) => 
                           a(23), a(22) => a(22), a(21) => a(21), a(20) => 
                           a(20), a(19) => a(19), a(18) => a(18), a(17) => 
                           a(17), a(16) => a(16), a(15) => a(15), a(14) => 
                           a(14), a(13) => a(13), a(12) => a(12), a(11) => 
                           a(11), a(10) => a(10), a(9) => a(9), a(8) => a(8), 
                           a(7) => a(7), a(6) => a(6), a(5) => a(5), a(4) => 
                           a(4), a(3) => a(3), a(2) => a(2), a(1) => a(1), a(0)
                           => a(0), b(63) => b(63), b(62) => b(62), b(61) => 
                           b(61), b(60) => b(60), b(59) => b(59), b(58) => 
                           b(58), b(57) => b(57), b(56) => b(56), b(55) => 
                           b(55), b(54) => b(54), b(53) => b(53), b(52) => 
                           b(52), b(51) => b(51), b(50) => b(50), b(49) => 
                           b(49), b(48) => b(48), b(47) => b(47), b(46) => 
                           b(46), b(45) => b(45), b(44) => b(44), b(43) => 
                           b(43), b(42) => b(42), b(41) => b(41), b(40) => 
                           b(40), b(39) => b(39), b(38) => b(38), b(37) => 
                           b(37), b(36) => b(36), b(35) => b(35), b(34) => 
                           b(34), b(33) => b(33), b(32) => b(32), b(31) => 
                           b(31), b(30) => b(30), b(29) => b(29), b(28) => 
                           b(28), b(27) => b(27), b(26) => b(26), b(25) => 
                           b(25), b(24) => b(24), b(23) => b(23), b(22) => 
                           b(22), b(21) => b(21), b(20) => b(20), b(19) => 
                           b(19), b(18) => b(18), b(17) => b(17), b(16) => 
                           b(16), b(15) => b(15), b(14) => b(14), b(13) => 
                           b(13), b(12) => b(12), b(11) => b(11), b(10) => 
                           b(10), b(9) => b(9), b(8) => b(8), b(7) => b(7), 
                           b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3) => 
                           b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), cin 
                           => cin, cout(15) => cout, cout(14) => carry_15_port,
                           cout(13) => carry_14_port, cout(12) => carry_13_port
                           , cout(11) => carry_12_port, cout(10) => 
                           carry_11_port, cout(9) => carry_10_port, cout(8) => 
                           carry_9_port, cout(7) => carry_8_port, cout(6) => 
                           carry_7_port, cout(5) => carry_6_port, cout(4) => 
                           carry_5_port, cout(3) => carry_4_port, cout(2) => 
                           carry_3_port, cout(1) => carry_2_port, cout(0) => 
                           carry_1_port);
   SG0 : AdderSumGenerator_DATA_SIZE64_SPARSITY4 port map( a(63) => a(63), 
                           a(62) => a(62), a(61) => a(61), a(60) => a(60), 
                           a(59) => a(59), a(58) => a(58), a(57) => a(57), 
                           a(56) => a(56), a(55) => a(55), a(54) => a(54), 
                           a(53) => a(53), a(52) => a(52), a(51) => a(51), 
                           a(50) => a(50), a(49) => a(49), a(48) => a(48), 
                           a(47) => a(47), a(46) => a(46), a(45) => a(45), 
                           a(44) => a(44), a(43) => a(43), a(42) => a(42), 
                           a(41) => a(41), a(40) => a(40), a(39) => a(39), 
                           a(38) => a(38), a(37) => a(37), a(36) => a(36), 
                           a(35) => a(35), a(34) => a(34), a(33) => a(33), 
                           a(32) => a(32), a(31) => a(31), a(30) => a(30), 
                           a(29) => a(29), a(28) => a(28), a(27) => a(27), 
                           a(26) => a(26), a(25) => a(25), a(24) => a(24), 
                           a(23) => a(23), a(22) => a(22), a(21) => a(21), 
                           a(20) => a(20), a(19) => a(19), a(18) => a(18), 
                           a(17) => a(17), a(16) => a(16), a(15) => a(15), 
                           a(14) => a(14), a(13) => a(13), a(12) => a(12), 
                           a(11) => a(11), a(10) => a(10), a(9) => a(9), a(8) 
                           => a(8), a(7) => a(7), a(6) => a(6), a(5) => a(5), 
                           a(4) => a(4), a(3) => a(3), a(2) => a(2), a(1) => 
                           a(1), a(0) => a(0), b(63) => b(63), b(62) => b(62), 
                           b(61) => b(61), b(60) => b(60), b(59) => b(59), 
                           b(58) => b(58), b(57) => b(57), b(56) => b(56), 
                           b(55) => b(55), b(54) => b(54), b(53) => b(53), 
                           b(52) => b(52), b(51) => b(51), b(50) => b(50), 
                           b(49) => b(49), b(48) => b(48), b(47) => b(47), 
                           b(46) => b(46), b(45) => b(45), b(44) => b(44), 
                           b(43) => b(43), b(42) => b(42), b(41) => b(41), 
                           b(40) => b(40), b(39) => b(39), b(38) => b(38), 
                           b(37) => b(37), b(36) => b(36), b(35) => b(35), 
                           b(34) => b(34), b(33) => b(33), b(32) => b(32), 
                           b(31) => b(31), b(30) => b(30), b(29) => b(29), 
                           b(28) => b(28), b(27) => b(27), b(26) => b(26), 
                           b(25) => b(25), b(24) => b(24), b(23) => b(23), 
                           b(22) => b(22), b(21) => b(21), b(20) => b(20), 
                           b(19) => b(19), b(18) => b(18), b(17) => b(17), 
                           b(16) => b(16), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => n1, b(4) => b(4), b(3) 
                           => n4, b(2) => n5, b(1) => n2, b(0) => n3, cin(15) 
                           => carry_15_port, cin(14) => carry_14_port, cin(13) 
                           => carry_13_port, cin(12) => carry_12_port, cin(11) 
                           => carry_11_port, cin(10) => carry_10_port, cin(9) 
                           => carry_9_port, cin(8) => carry_8_port, cin(7) => 
                           carry_7_port, cin(6) => carry_6_port, cin(5) => 
                           carry_5_port, cin(4) => carry_4_port, cin(3) => 
                           carry_3_port, cin(2) => carry_2_port, cin(1) => 
                           carry_1_port, cin(0) => cin, sum(63) => s(63), 
                           sum(62) => s(62), sum(61) => s(61), sum(60) => s(60)
                           , sum(59) => s(59), sum(58) => s(58), sum(57) => 
                           s(57), sum(56) => s(56), sum(55) => s(55), sum(54) 
                           => s(54), sum(53) => s(53), sum(52) => s(52), 
                           sum(51) => s(51), sum(50) => s(50), sum(49) => s(49)
                           , sum(48) => s(48), sum(47) => s(47), sum(46) => 
                           s(46), sum(45) => s(45), sum(44) => s(44), sum(43) 
                           => s(43), sum(42) => s(42), sum(41) => s(41), 
                           sum(40) => s(40), sum(39) => s(39), sum(38) => s(38)
                           , sum(37) => s(37), sum(36) => s(36), sum(35) => 
                           s(35), sum(34) => s(34), sum(33) => s(33), sum(32) 
                           => s(32), sum(31) => s(31), sum(30) => s(30), 
                           sum(29) => s(29), sum(28) => s(28), sum(27) => s(27)
                           , sum(26) => s(26), sum(25) => s(25), sum(24) => 
                           s(24), sum(23) => s(23), sum(22) => s(22), sum(21) 
                           => s(21), sum(20) => s(20), sum(19) => s(19), 
                           sum(18) => s(18), sum(17) => s(17), sum(16) => s(16)
                           , sum(15) => s(15), sum(14) => s(14), sum(13) => 
                           s(13), sum(12) => s(12), sum(11) => s(11), sum(10) 
                           => s(10), sum(9) => s(9), sum(8) => s(8), sum(7) => 
                           s(7), sum(6) => s(6), sum(5) => s(5), sum(4) => s(4)
                           , sum(3) => s(3), sum(2) => s(2), sum(1) => s(1), 
                           sum(0) => s(0));
   U1 : CLKBUF_X1 port map( A => b(5), Z => n1);
   U2 : CLKBUF_X1 port map( A => b(2), Z => n5);
   U3 : CLKBUF_X1 port map( A => b(1), Z => n2);
   U4 : CLKBUF_X1 port map( A => b(0), Z => n3);
   U5 : CLKBUF_X1 port map( A => b(3), Z => n4);

end SYN_p4_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4Adder_DATA_SIZE16_SPARSITY4 is

   port( cin : in std_logic;  a, b : in std_logic_vector (15 downto 0);  s : 
         out std_logic_vector (15 downto 0);  cout : out std_logic);

end P4Adder_DATA_SIZE16_SPARSITY4;

architecture SYN_p4_adder_arch of P4Adder_DATA_SIZE16_SPARSITY4 is

   component AdderSumGenerator_DATA_SIZE16_SPARSITY4
      port( a, b : in std_logic_vector (15 downto 0);  cin : in 
            std_logic_vector (3 downto 0);  sum : out std_logic_vector (15 
            downto 0));
   end component;
   
   component P4CarryGenerator_DATA_SIZE16_SPARSITY4
      port( a, b : in std_logic_vector (15 downto 0);  cin : in std_logic;  
            cout : out std_logic_vector (3 downto 0));
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   CG0 : P4CarryGenerator_DATA_SIZE16_SPARSITY4 port map( a(15) => a(15), a(14)
                           => a(14), a(13) => a(13), a(12) => a(12), a(11) => 
                           a(11), a(10) => a(10), a(9) => a(9), a(8) => a(8), 
                           a(7) => a(7), a(6) => a(6), a(5) => a(5), a(4) => 
                           a(4), a(3) => a(3), a(2) => a(2), a(1) => a(1), a(0)
                           => a(0), b(15) => b(15), b(14) => b(14), b(13) => 
                           b(13), b(12) => b(12), b(11) => b(11), b(10) => 
                           b(10), b(9) => b(9), b(8) => b(8), b(7) => b(7), 
                           b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3) => 
                           b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), cin 
                           => cin, cout(3) => cout, cout(2) => carry_3_port, 
                           cout(1) => carry_2_port, cout(0) => carry_1_port);
   SG0 : AdderSumGenerator_DATA_SIZE16_SPARSITY4 port map( a(15) => a(15), 
                           a(14) => a(14), a(13) => a(13), a(12) => a(12), 
                           a(11) => a(11), a(10) => a(10), a(9) => a(9), a(8) 
                           => a(8), a(7) => a(7), a(6) => a(6), a(5) => a(5), 
                           a(4) => a(4), a(3) => a(3), a(2) => a(2), a(1) => 
                           a(1), a(0) => a(0), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           cin(3) => carry_3_port, cin(2) => carry_2_port, 
                           cin(1) => carry_1_port, cin(0) => cin, sum(15) => 
                           s(15), sum(14) => s(14), sum(13) => s(13), sum(12) 
                           => s(12), sum(11) => s(11), sum(10) => s(10), sum(9)
                           => s(9), sum(8) => s(8), sum(7) => s(7), sum(6) => 
                           s(6), sum(5) => s(5), sum(4) => s(4), sum(3) => s(3)
                           , sum(2) => s(2), sum(1) => s(1), sum(0) => s(0));

end SYN_p4_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_0 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_0;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_0 is

   component Mux_DATA_SIZE4_0
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_167
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_0
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_0 port map( ci => X_Logic0_port, a(3) => a(3), a(2) =>
                           a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2)
                           => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_167 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_0 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Adder_DATA_SIZE64 is

   port( cin : in std_logic;  a, b : in std_logic_vector (63 downto 0);  s : 
         out std_logic_vector (63 downto 0);  cout : out std_logic);

end Adder_DATA_SIZE64;

architecture SYN_adder_arch of Adder_DATA_SIZE64 is

   component P4Adder_DATA_SIZE64_SPARSITY4
      port( cin : in std_logic;  a, b : in std_logic_vector (63 downto 0);  s :
            out std_logic_vector (63 downto 0);  cout : out std_logic);
   end component;

begin
   
   ADDER0 : P4Adder_DATA_SIZE64_SPARSITY4 port map( cin => cin, a(63) => a(63),
                           a(62) => a(62), a(61) => a(61), a(60) => a(60), 
                           a(59) => a(59), a(58) => a(58), a(57) => a(57), 
                           a(56) => a(56), a(55) => a(55), a(54) => a(54), 
                           a(53) => a(53), a(52) => a(52), a(51) => a(51), 
                           a(50) => a(50), a(49) => a(49), a(48) => a(48), 
                           a(47) => a(47), a(46) => a(46), a(45) => a(45), 
                           a(44) => a(44), a(43) => a(43), a(42) => a(42), 
                           a(41) => a(41), a(40) => a(40), a(39) => a(39), 
                           a(38) => a(38), a(37) => a(37), a(36) => a(36), 
                           a(35) => a(35), a(34) => a(34), a(33) => a(33), 
                           a(32) => a(32), a(31) => a(31), a(30) => a(30), 
                           a(29) => a(29), a(28) => a(28), a(27) => a(27), 
                           a(26) => a(26), a(25) => a(25), a(24) => a(24), 
                           a(23) => a(23), a(22) => a(22), a(21) => a(21), 
                           a(20) => a(20), a(19) => a(19), a(18) => a(18), 
                           a(17) => a(17), a(16) => a(16), a(15) => a(15), 
                           a(14) => a(14), a(13) => a(13), a(12) => a(12), 
                           a(11) => a(11), a(10) => a(10), a(9) => a(9), a(8) 
                           => a(8), a(7) => a(7), a(6) => a(6), a(5) => a(5), 
                           a(4) => a(4), a(3) => a(3), a(2) => a(2), a(1) => 
                           a(1), a(0) => a(0), b(63) => b(63), b(62) => b(62), 
                           b(61) => b(61), b(60) => b(60), b(59) => b(59), 
                           b(58) => b(58), b(57) => b(57), b(56) => b(56), 
                           b(55) => b(55), b(54) => b(54), b(53) => b(53), 
                           b(52) => b(52), b(51) => b(51), b(50) => b(50), 
                           b(49) => b(49), b(48) => b(48), b(47) => b(47), 
                           b(46) => b(46), b(45) => b(45), b(44) => b(44), 
                           b(43) => b(43), b(42) => b(42), b(41) => b(41), 
                           b(40) => b(40), b(39) => b(39), b(38) => b(38), 
                           b(37) => b(37), b(36) => b(36), b(35) => b(35), 
                           b(34) => b(34), b(33) => b(33), b(32) => b(32), 
                           b(31) => b(31), b(30) => b(30), b(29) => b(29), 
                           b(28) => b(28), b(27) => b(27), b(26) => b(26), 
                           b(25) => b(25), b(24) => b(24), b(23) => b(23), 
                           b(22) => b(22), b(21) => b(21), b(20) => b(20), 
                           b(19) => b(19), b(18) => b(18), b(17) => b(17), 
                           b(16) => b(16), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           s(63) => s(63), s(62) => s(62), s(61) => s(61), 
                           s(60) => s(60), s(59) => s(59), s(58) => s(58), 
                           s(57) => s(57), s(56) => s(56), s(55) => s(55), 
                           s(54) => s(54), s(53) => s(53), s(52) => s(52), 
                           s(51) => s(51), s(50) => s(50), s(49) => s(49), 
                           s(48) => s(48), s(47) => s(47), s(46) => s(46), 
                           s(45) => s(45), s(44) => s(44), s(43) => s(43), 
                           s(42) => s(42), s(41) => s(41), s(40) => s(40), 
                           s(39) => s(39), s(38) => s(38), s(37) => s(37), 
                           s(36) => s(36), s(35) => s(35), s(34) => s(34), 
                           s(33) => s(33), s(32) => s(32), s(31) => s(31), 
                           s(30) => s(30), s(29) => s(29), s(28) => s(28), 
                           s(27) => s(27), s(26) => s(26), s(25) => s(25), 
                           s(24) => s(24), s(23) => s(23), s(22) => s(22), 
                           s(21) => s(21), s(20) => s(20), s(19) => s(19), 
                           s(18) => s(18), s(17) => s(17), s(16) => s(16), 
                           s(15) => s(15), s(14) => s(14), s(13) => s(13), 
                           s(12) => s(12), s(11) => s(11), s(10) => s(10), s(9)
                           => s(9), s(8) => s(8), s(7) => s(7), s(6) => s(6), 
                           s(5) => s(5), s(4) => s(4), s(3) => s(3), s(2) => 
                           s(2), s(1) => s(1), s(0) => s(0), cout => cout);

end SYN_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity BoothMul_DATA_SIZE16_STAGE10_DW01_inc_0 is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end BoothMul_DATA_SIZE16_STAGE10_DW01_inc_0;

architecture SYN_rpl of BoothMul_DATA_SIZE16_STAGE10_DW01_inc_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port : std_logic;

begin
   
   U1_1_30 : HA_X1 port map( A => A(30), B => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_1_29 : HA_X1 port map( A => A(29), B => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_1_28 : HA_X1 port map( A => A(28), B => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_1_27 : HA_X1 port map( A => A(27), B => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_1_26 : HA_X1 port map( A => A(26), B => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_1_25 : HA_X1 port map( A => A(25), B => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_1_24 : HA_X1 port map( A => A(24), B => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_1_23 : HA_X1 port map( A => A(23), B => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_1_22 : HA_X1 port map( A => A(22), B => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_1_21 : HA_X1 port map( A => A(21), B => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_1_20 : HA_X1 port map( A => A(20), B => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_1_19 : HA_X1 port map( A => A(19), B => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_1_18 : HA_X1 port map( A => A(18), B => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_1_17 : HA_X1 port map( A => A(17), B => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_1_16 : HA_X1 port map( A => A(16), B => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_1_15 : HA_X1 port map( A => A(15), B => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : XOR2_X1 port map( A => carry_31_port, B => A(31), Z => SUM(31));
   U2 : INV_X1 port map( A => A(0), ZN => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity BoothEncoder is

   port( din : in std_logic_vector (2 downto 0);  sel : out std_logic_vector (2
         downto 0));

end BoothEncoder;

architecture SYN_booth_encoder_arch of BoothEncoder is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n8, n9, n10 : std_logic;

begin
   
   U10 : NAND3_X1 port map( A1 => din(0), A2 => n7, A3 => din(1), ZN => n8);
   U3 : INV_X1 port map( A => din(0), ZN => n9);
   U4 : NAND2_X1 port map( A1 => din(2), A2 => n4, ZN => n10);
   U5 : OAI21_X1 port map( B1 => n6, B2 => din(1), A => n8, ZN => sel(0));
   U6 : OAI221_X1 port map( B1 => din(1), B2 => n4, C1 => din(2), C2 => n5, A 
                           => n10, ZN => sel(2));
   U7 : INV_X1 port map( A => din(1), ZN => n5);
   U8 : OAI21_X1 port map( B1 => din(1), B2 => n7, A => n10, ZN => sel(1));
   U9 : INV_X1 port map( A => din(2), ZN => n7);
   U11 : INV_X1 port map( A => din(0), ZN => n4);
   U12 : NAND2_X1 port map( A1 => din(2), A2 => n9, ZN => n6);

end SYN_booth_encoder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Adder_DATA_SIZE16 is

   port( cin : in std_logic;  a, b : in std_logic_vector (15 downto 0);  s : 
         out std_logic_vector (15 downto 0);  cout : out std_logic);

end Adder_DATA_SIZE16;

architecture SYN_adder_arch of Adder_DATA_SIZE16 is

   component P4Adder_DATA_SIZE16_SPARSITY4
      port( cin : in std_logic;  a, b : in std_logic_vector (15 downto 0);  s :
            out std_logic_vector (15 downto 0);  cout : out std_logic);
   end component;

begin
   
   ADDER0 : P4Adder_DATA_SIZE16_SPARSITY4 port map( cin => cin, a(15) => a(15),
                           a(14) => a(14), a(13) => a(13), a(12) => a(12), 
                           a(11) => a(11), a(10) => a(10), a(9) => a(9), a(8) 
                           => a(8), a(7) => a(7), a(6) => a(6), a(5) => a(5), 
                           a(4) => a(4), a(3) => a(3), a(2) => a(2), a(1) => 
                           a(1), a(0) => a(0), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           s(15) => s(15), s(14) => s(14), s(13) => s(13), 
                           s(12) => s(12), s(11) => s(11), s(10) => s(10), s(9)
                           => s(9), s(8) => s(8), s(7) => s(7), s(6) => s(6), 
                           s(5) => s(5), s(4) => s(4), s(3) => s(3), s(2) => 
                           s(2), s(1) => s(1), s(0) => s(0), cout => cout);

end SYN_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Shifter_DATA_SIZE32_DW_rbsh_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end Shifter_DATA_SIZE32_DW_rbsh_0;

architecture SYN_mx2 of Shifter_DATA_SIZE32_DW_rbsh_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal MR_int_1_31_port, MR_int_1_30_port, MR_int_1_29_port, 
      MR_int_1_28_port, MR_int_1_27_port, MR_int_1_26_port, MR_int_1_25_port, 
      MR_int_1_24_port, MR_int_1_23_port, MR_int_1_22_port, MR_int_1_21_port, 
      MR_int_1_20_port, MR_int_1_19_port, MR_int_1_18_port, MR_int_1_17_port, 
      MR_int_1_16_port, MR_int_1_15_port, MR_int_1_14_port, MR_int_1_13_port, 
      MR_int_1_12_port, MR_int_1_11_port, MR_int_1_10_port, MR_int_1_9_port, 
      MR_int_1_8_port, MR_int_1_7_port, MR_int_1_6_port, MR_int_1_5_port, 
      MR_int_1_4_port, MR_int_1_3_port, MR_int_1_2_port, MR_int_1_1_port, 
      MR_int_1_0_port, MR_int_2_31_port, MR_int_2_30_port, MR_int_2_29_port, 
      MR_int_2_28_port, MR_int_2_27_port, MR_int_2_26_port, MR_int_2_25_port, 
      MR_int_2_24_port, MR_int_2_23_port, MR_int_2_22_port, MR_int_2_21_port, 
      MR_int_2_20_port, MR_int_2_19_port, MR_int_2_18_port, MR_int_2_17_port, 
      MR_int_2_16_port, MR_int_2_15_port, MR_int_2_14_port, MR_int_2_13_port, 
      MR_int_2_12_port, MR_int_2_11_port, MR_int_2_10_port, MR_int_2_9_port, 
      MR_int_2_8_port, MR_int_2_7_port, MR_int_2_6_port, MR_int_2_5_port, 
      MR_int_2_4_port, MR_int_2_3_port, MR_int_2_2_port, MR_int_2_1_port, 
      MR_int_2_0_port, MR_int_3_31_port, MR_int_3_30_port, MR_int_3_29_port, 
      MR_int_3_28_port, MR_int_3_27_port, MR_int_3_26_port, MR_int_3_25_port, 
      MR_int_3_24_port, MR_int_3_23_port, MR_int_3_22_port, MR_int_3_21_port, 
      MR_int_3_20_port, MR_int_3_19_port, MR_int_3_18_port, MR_int_3_17_port, 
      MR_int_3_16_port, MR_int_3_15_port, MR_int_3_14_port, MR_int_3_13_port, 
      MR_int_3_12_port, MR_int_3_11_port, MR_int_3_10_port, MR_int_3_9_port, 
      MR_int_3_8_port, MR_int_3_7_port, MR_int_3_6_port, MR_int_3_5_port, 
      MR_int_3_4_port, MR_int_3_3_port, MR_int_3_2_port, MR_int_3_1_port, 
      MR_int_3_0_port, MR_int_4_31_port, MR_int_4_30_port, MR_int_4_29_port, 
      MR_int_4_28_port, MR_int_4_27_port, MR_int_4_26_port, MR_int_4_25_port, 
      MR_int_4_24_port, MR_int_4_23_port, MR_int_4_22_port, MR_int_4_21_port, 
      MR_int_4_20_port, MR_int_4_19_port, MR_int_4_18_port, MR_int_4_17_port, 
      MR_int_4_16_port, MR_int_4_15_port, MR_int_4_14_port, MR_int_4_13_port, 
      MR_int_4_12_port, MR_int_4_11_port, MR_int_4_10_port, MR_int_4_9_port, 
      MR_int_4_8_port, MR_int_4_7_port, MR_int_4_6_port, MR_int_4_5_port, 
      MR_int_4_4_port, MR_int_4_3_port, MR_int_4_2_port, MR_int_4_1_port, 
      MR_int_4_0_port, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, 
      n16, n17, n18 : std_logic;

begin
   
   M1_4_31 : MUX2_X1 port map( A => MR_int_4_31_port, B => MR_int_4_15_port, S 
                           => n18, Z => B(31));
   M1_4_30 : MUX2_X1 port map( A => MR_int_4_30_port, B => MR_int_4_14_port, S 
                           => n18, Z => B(30));
   M1_4_29 : MUX2_X1 port map( A => MR_int_4_29_port, B => MR_int_4_13_port, S 
                           => n18, Z => B(29));
   M1_4_28 : MUX2_X1 port map( A => MR_int_4_28_port, B => MR_int_4_12_port, S 
                           => n18, Z => B(28));
   M1_4_27 : MUX2_X1 port map( A => MR_int_4_27_port, B => MR_int_4_11_port, S 
                           => n18, Z => B(27));
   M1_4_26 : MUX2_X1 port map( A => MR_int_4_26_port, B => MR_int_4_10_port, S 
                           => n18, Z => B(26));
   M1_4_25 : MUX2_X1 port map( A => MR_int_4_25_port, B => MR_int_4_9_port, S 
                           => n18, Z => B(25));
   M1_4_24 : MUX2_X1 port map( A => MR_int_4_24_port, B => MR_int_4_8_port, S 
                           => n18, Z => B(24));
   M1_4_23 : MUX2_X1 port map( A => MR_int_4_23_port, B => MR_int_4_7_port, S 
                           => n17, Z => B(23));
   M1_4_22 : MUX2_X1 port map( A => MR_int_4_22_port, B => MR_int_4_6_port, S 
                           => n17, Z => B(22));
   M1_4_21 : MUX2_X1 port map( A => MR_int_4_21_port, B => MR_int_4_5_port, S 
                           => n17, Z => B(21));
   M1_4_20 : MUX2_X1 port map( A => MR_int_4_20_port, B => MR_int_4_4_port, S 
                           => n17, Z => B(20));
   M1_4_19 : MUX2_X1 port map( A => MR_int_4_19_port, B => MR_int_4_3_port, S 
                           => n17, Z => B(19));
   M1_4_18 : MUX2_X1 port map( A => MR_int_4_18_port, B => MR_int_4_2_port, S 
                           => n17, Z => B(18));
   M1_4_17 : MUX2_X1 port map( A => MR_int_4_17_port, B => MR_int_4_1_port, S 
                           => n17, Z => B(17));
   M1_4_16 : MUX2_X1 port map( A => MR_int_4_16_port, B => MR_int_4_0_port, S 
                           => n17, Z => B(16));
   M1_4_15 : MUX2_X1 port map( A => MR_int_4_15_port, B => MR_int_4_31_port, S 
                           => n17, Z => B(15));
   M1_4_14 : MUX2_X1 port map( A => MR_int_4_14_port, B => MR_int_4_30_port, S 
                           => n17, Z => B(14));
   M1_4_13 : MUX2_X1 port map( A => MR_int_4_13_port, B => MR_int_4_29_port, S 
                           => n17, Z => B(13));
   M1_4_12 : MUX2_X1 port map( A => MR_int_4_12_port, B => MR_int_4_28_port, S 
                           => n17, Z => B(12));
   M1_4_11 : MUX2_X1 port map( A => MR_int_4_11_port, B => MR_int_4_27_port, S 
                           => n16, Z => B(11));
   M1_4_10 : MUX2_X1 port map( A => MR_int_4_10_port, B => MR_int_4_26_port, S 
                           => n16, Z => B(10));
   M1_4_9 : MUX2_X1 port map( A => MR_int_4_9_port, B => MR_int_4_25_port, S =>
                           n16, Z => B(9));
   M1_4_8 : MUX2_X1 port map( A => MR_int_4_8_port, B => MR_int_4_24_port, S =>
                           n16, Z => B(8));
   M1_4_7 : MUX2_X1 port map( A => MR_int_4_7_port, B => MR_int_4_23_port, S =>
                           n16, Z => B(7));
   M1_4_6 : MUX2_X1 port map( A => MR_int_4_6_port, B => MR_int_4_22_port, S =>
                           n16, Z => B(6));
   M1_4_5 : MUX2_X1 port map( A => MR_int_4_5_port, B => MR_int_4_21_port, S =>
                           n16, Z => B(5));
   M1_4_4 : MUX2_X1 port map( A => MR_int_4_4_port, B => MR_int_4_20_port, S =>
                           n16, Z => B(4));
   M1_4_3 : MUX2_X1 port map( A => MR_int_4_3_port, B => MR_int_4_19_port, S =>
                           n16, Z => B(3));
   M1_4_2 : MUX2_X1 port map( A => MR_int_4_2_port, B => MR_int_4_18_port, S =>
                           n16, Z => B(2));
   M1_4_1 : MUX2_X1 port map( A => MR_int_4_1_port, B => MR_int_4_17_port, S =>
                           n16, Z => B(1));
   M1_4_0 : MUX2_X1 port map( A => MR_int_4_0_port, B => MR_int_4_16_port, S =>
                           n16, Z => B(0));
   M1_3_31_0 : MUX2_X1 port map( A => MR_int_3_31_port, B => MR_int_3_7_port, S
                           => n15, Z => MR_int_4_31_port);
   M1_3_30_0 : MUX2_X1 port map( A => MR_int_3_30_port, B => MR_int_3_6_port, S
                           => n15, Z => MR_int_4_30_port);
   M1_3_29_0 : MUX2_X1 port map( A => MR_int_3_29_port, B => MR_int_3_5_port, S
                           => n15, Z => MR_int_4_29_port);
   M1_3_28_0 : MUX2_X1 port map( A => MR_int_3_28_port, B => MR_int_3_4_port, S
                           => n15, Z => MR_int_4_28_port);
   M1_3_27_0 : MUX2_X1 port map( A => MR_int_3_27_port, B => MR_int_3_3_port, S
                           => n15, Z => MR_int_4_27_port);
   M1_3_26_0 : MUX2_X1 port map( A => MR_int_3_26_port, B => MR_int_3_2_port, S
                           => n15, Z => MR_int_4_26_port);
   M1_3_25_0 : MUX2_X1 port map( A => MR_int_3_25_port, B => MR_int_3_1_port, S
                           => n15, Z => MR_int_4_25_port);
   M1_3_24_0 : MUX2_X1 port map( A => MR_int_3_24_port, B => MR_int_3_0_port, S
                           => n15, Z => MR_int_4_24_port);
   M1_3_23_0 : MUX2_X1 port map( A => MR_int_3_23_port, B => MR_int_3_31_port, 
                           S => n14, Z => MR_int_4_23_port);
   M1_3_22_0 : MUX2_X1 port map( A => MR_int_3_22_port, B => MR_int_3_30_port, 
                           S => n14, Z => MR_int_4_22_port);
   M1_3_21_0 : MUX2_X1 port map( A => MR_int_3_21_port, B => MR_int_3_29_port, 
                           S => n14, Z => MR_int_4_21_port);
   M1_3_20_0 : MUX2_X1 port map( A => MR_int_3_20_port, B => MR_int_3_28_port, 
                           S => n14, Z => MR_int_4_20_port);
   M1_3_19_0 : MUX2_X1 port map( A => MR_int_3_19_port, B => MR_int_3_27_port, 
                           S => n14, Z => MR_int_4_19_port);
   M1_3_18_0 : MUX2_X1 port map( A => MR_int_3_18_port, B => MR_int_3_26_port, 
                           S => n14, Z => MR_int_4_18_port);
   M1_3_17_0 : MUX2_X1 port map( A => MR_int_3_17_port, B => MR_int_3_25_port, 
                           S => n14, Z => MR_int_4_17_port);
   M1_3_16_0 : MUX2_X1 port map( A => MR_int_3_16_port, B => MR_int_3_24_port, 
                           S => n14, Z => MR_int_4_16_port);
   M1_3_15_0 : MUX2_X1 port map( A => MR_int_3_15_port, B => MR_int_3_23_port, 
                           S => n14, Z => MR_int_4_15_port);
   M1_3_14_0 : MUX2_X1 port map( A => MR_int_3_14_port, B => MR_int_3_22_port, 
                           S => n14, Z => MR_int_4_14_port);
   M1_3_13_0 : MUX2_X1 port map( A => MR_int_3_13_port, B => MR_int_3_21_port, 
                           S => n14, Z => MR_int_4_13_port);
   M1_3_12_0 : MUX2_X1 port map( A => MR_int_3_12_port, B => MR_int_3_20_port, 
                           S => n14, Z => MR_int_4_12_port);
   M1_3_11_0 : MUX2_X1 port map( A => MR_int_3_11_port, B => MR_int_3_19_port, 
                           S => n13, Z => MR_int_4_11_port);
   M1_3_10_0 : MUX2_X1 port map( A => MR_int_3_10_port, B => MR_int_3_18_port, 
                           S => n13, Z => MR_int_4_10_port);
   M1_3_9_0 : MUX2_X1 port map( A => MR_int_3_9_port, B => MR_int_3_17_port, S 
                           => n13, Z => MR_int_4_9_port);
   M1_3_8_0 : MUX2_X1 port map( A => MR_int_3_8_port, B => MR_int_3_16_port, S 
                           => n13, Z => MR_int_4_8_port);
   M1_3_7 : MUX2_X1 port map( A => MR_int_3_7_port, B => MR_int_3_15_port, S =>
                           n13, Z => MR_int_4_7_port);
   M1_3_6 : MUX2_X1 port map( A => MR_int_3_6_port, B => MR_int_3_14_port, S =>
                           n13, Z => MR_int_4_6_port);
   M1_3_5 : MUX2_X1 port map( A => MR_int_3_5_port, B => MR_int_3_13_port, S =>
                           n13, Z => MR_int_4_5_port);
   M1_3_4 : MUX2_X1 port map( A => MR_int_3_4_port, B => MR_int_3_12_port, S =>
                           n13, Z => MR_int_4_4_port);
   M1_3_3 : MUX2_X1 port map( A => MR_int_3_3_port, B => MR_int_3_11_port, S =>
                           n13, Z => MR_int_4_3_port);
   M1_3_2 : MUX2_X1 port map( A => MR_int_3_2_port, B => MR_int_3_10_port, S =>
                           n13, Z => MR_int_4_2_port);
   M1_3_1 : MUX2_X1 port map( A => MR_int_3_1_port, B => MR_int_3_9_port, S => 
                           n13, Z => MR_int_4_1_port);
   M1_3_0 : MUX2_X1 port map( A => MR_int_3_0_port, B => MR_int_3_8_port, S => 
                           n13, Z => MR_int_4_0_port);
   M1_2_31_0 : MUX2_X1 port map( A => MR_int_2_31_port, B => MR_int_2_3_port, S
                           => n12, Z => MR_int_3_31_port);
   M1_2_30_0 : MUX2_X1 port map( A => MR_int_2_30_port, B => MR_int_2_2_port, S
                           => n12, Z => MR_int_3_30_port);
   M1_2_29_0 : MUX2_X1 port map( A => MR_int_2_29_port, B => MR_int_2_1_port, S
                           => n12, Z => MR_int_3_29_port);
   M1_2_28_0 : MUX2_X1 port map( A => MR_int_2_28_port, B => MR_int_2_0_port, S
                           => n12, Z => MR_int_3_28_port);
   M1_2_27_0 : MUX2_X1 port map( A => MR_int_2_27_port, B => MR_int_2_31_port, 
                           S => n12, Z => MR_int_3_27_port);
   M1_2_26_0 : MUX2_X1 port map( A => MR_int_2_26_port, B => MR_int_2_30_port, 
                           S => n12, Z => MR_int_3_26_port);
   M1_2_25_0 : MUX2_X1 port map( A => MR_int_2_25_port, B => MR_int_2_29_port, 
                           S => n12, Z => MR_int_3_25_port);
   M1_2_24_0 : MUX2_X1 port map( A => MR_int_2_24_port, B => MR_int_2_28_port, 
                           S => n12, Z => MR_int_3_24_port);
   M1_2_23_0 : MUX2_X1 port map( A => MR_int_2_23_port, B => MR_int_2_27_port, 
                           S => n11, Z => MR_int_3_23_port);
   M1_2_22_0 : MUX2_X1 port map( A => MR_int_2_22_port, B => MR_int_2_26_port, 
                           S => n11, Z => MR_int_3_22_port);
   M1_2_21_0 : MUX2_X1 port map( A => MR_int_2_21_port, B => MR_int_2_25_port, 
                           S => n11, Z => MR_int_3_21_port);
   M1_2_20_0 : MUX2_X1 port map( A => MR_int_2_20_port, B => MR_int_2_24_port, 
                           S => n11, Z => MR_int_3_20_port);
   M1_2_19_0 : MUX2_X1 port map( A => MR_int_2_19_port, B => MR_int_2_23_port, 
                           S => n11, Z => MR_int_3_19_port);
   M1_2_18_0 : MUX2_X1 port map( A => MR_int_2_18_port, B => MR_int_2_22_port, 
                           S => n11, Z => MR_int_3_18_port);
   M1_2_17_0 : MUX2_X1 port map( A => MR_int_2_17_port, B => MR_int_2_21_port, 
                           S => n11, Z => MR_int_3_17_port);
   M1_2_16_0 : MUX2_X1 port map( A => MR_int_2_16_port, B => MR_int_2_20_port, 
                           S => n11, Z => MR_int_3_16_port);
   M1_2_15_0 : MUX2_X1 port map( A => MR_int_2_15_port, B => MR_int_2_19_port, 
                           S => n11, Z => MR_int_3_15_port);
   M1_2_14_0 : MUX2_X1 port map( A => MR_int_2_14_port, B => MR_int_2_18_port, 
                           S => n11, Z => MR_int_3_14_port);
   M1_2_13_0 : MUX2_X1 port map( A => MR_int_2_13_port, B => MR_int_2_17_port, 
                           S => n11, Z => MR_int_3_13_port);
   M1_2_12_0 : MUX2_X1 port map( A => MR_int_2_12_port, B => MR_int_2_16_port, 
                           S => n11, Z => MR_int_3_12_port);
   M1_2_11_0 : MUX2_X1 port map( A => MR_int_2_11_port, B => MR_int_2_15_port, 
                           S => n10, Z => MR_int_3_11_port);
   M1_2_10_0 : MUX2_X1 port map( A => MR_int_2_10_port, B => MR_int_2_14_port, 
                           S => n10, Z => MR_int_3_10_port);
   M1_2_9_0 : MUX2_X1 port map( A => MR_int_2_9_port, B => MR_int_2_13_port, S 
                           => n10, Z => MR_int_3_9_port);
   M1_2_8_0 : MUX2_X1 port map( A => MR_int_2_8_port, B => MR_int_2_12_port, S 
                           => n10, Z => MR_int_3_8_port);
   M1_2_7_0 : MUX2_X1 port map( A => MR_int_2_7_port, B => MR_int_2_11_port, S 
                           => n10, Z => MR_int_3_7_port);
   M1_2_6_0 : MUX2_X1 port map( A => MR_int_2_6_port, B => MR_int_2_10_port, S 
                           => n10, Z => MR_int_3_6_port);
   M1_2_5_0 : MUX2_X1 port map( A => MR_int_2_5_port, B => MR_int_2_9_port, S 
                           => n10, Z => MR_int_3_5_port);
   M1_2_4_0 : MUX2_X1 port map( A => MR_int_2_4_port, B => MR_int_2_8_port, S 
                           => n10, Z => MR_int_3_4_port);
   M1_2_3 : MUX2_X1 port map( A => MR_int_2_3_port, B => MR_int_2_7_port, S => 
                           n10, Z => MR_int_3_3_port);
   M1_2_2 : MUX2_X1 port map( A => MR_int_2_2_port, B => MR_int_2_6_port, S => 
                           n10, Z => MR_int_3_2_port);
   M1_2_1 : MUX2_X1 port map( A => MR_int_2_1_port, B => MR_int_2_5_port, S => 
                           n10, Z => MR_int_3_1_port);
   M1_2_0 : MUX2_X1 port map( A => MR_int_2_0_port, B => MR_int_2_4_port, S => 
                           n10, Z => MR_int_3_0_port);
   M1_1_31_0 : MUX2_X1 port map( A => MR_int_1_31_port, B => MR_int_1_1_port, S
                           => n9, Z => MR_int_2_31_port);
   M1_1_30_0 : MUX2_X1 port map( A => MR_int_1_30_port, B => MR_int_1_0_port, S
                           => n9, Z => MR_int_2_30_port);
   M1_1_29_0 : MUX2_X1 port map( A => MR_int_1_29_port, B => MR_int_1_31_port, 
                           S => n9, Z => MR_int_2_29_port);
   M1_1_28_0 : MUX2_X1 port map( A => MR_int_1_28_port, B => MR_int_1_30_port, 
                           S => n9, Z => MR_int_2_28_port);
   M1_1_27_0 : MUX2_X1 port map( A => MR_int_1_27_port, B => MR_int_1_29_port, 
                           S => n9, Z => MR_int_2_27_port);
   M1_1_26_0 : MUX2_X1 port map( A => MR_int_1_26_port, B => MR_int_1_28_port, 
                           S => n9, Z => MR_int_2_26_port);
   M1_1_25_0 : MUX2_X1 port map( A => MR_int_1_25_port, B => MR_int_1_27_port, 
                           S => n9, Z => MR_int_2_25_port);
   M1_1_24_0 : MUX2_X1 port map( A => MR_int_1_24_port, B => MR_int_1_26_port, 
                           S => n9, Z => MR_int_2_24_port);
   M1_1_23_0 : MUX2_X1 port map( A => MR_int_1_23_port, B => MR_int_1_25_port, 
                           S => n8, Z => MR_int_2_23_port);
   M1_1_22_0 : MUX2_X1 port map( A => MR_int_1_22_port, B => MR_int_1_24_port, 
                           S => n8, Z => MR_int_2_22_port);
   M1_1_21_0 : MUX2_X1 port map( A => MR_int_1_21_port, B => MR_int_1_23_port, 
                           S => n8, Z => MR_int_2_21_port);
   M1_1_20_0 : MUX2_X1 port map( A => MR_int_1_20_port, B => MR_int_1_22_port, 
                           S => n8, Z => MR_int_2_20_port);
   M1_1_19_0 : MUX2_X1 port map( A => MR_int_1_19_port, B => MR_int_1_21_port, 
                           S => n8, Z => MR_int_2_19_port);
   M1_1_18_0 : MUX2_X1 port map( A => MR_int_1_18_port, B => MR_int_1_20_port, 
                           S => n8, Z => MR_int_2_18_port);
   M1_1_17_0 : MUX2_X1 port map( A => MR_int_1_17_port, B => MR_int_1_19_port, 
                           S => n8, Z => MR_int_2_17_port);
   M1_1_16_0 : MUX2_X1 port map( A => MR_int_1_16_port, B => MR_int_1_18_port, 
                           S => n8, Z => MR_int_2_16_port);
   M1_1_15_0 : MUX2_X1 port map( A => MR_int_1_15_port, B => MR_int_1_17_port, 
                           S => n8, Z => MR_int_2_15_port);
   M1_1_14_0 : MUX2_X1 port map( A => MR_int_1_14_port, B => MR_int_1_16_port, 
                           S => n8, Z => MR_int_2_14_port);
   M1_1_13_0 : MUX2_X1 port map( A => MR_int_1_13_port, B => MR_int_1_15_port, 
                           S => n8, Z => MR_int_2_13_port);
   M1_1_12_0 : MUX2_X1 port map( A => MR_int_1_12_port, B => MR_int_1_14_port, 
                           S => n8, Z => MR_int_2_12_port);
   M1_1_11_0 : MUX2_X1 port map( A => MR_int_1_11_port, B => MR_int_1_13_port, 
                           S => n7, Z => MR_int_2_11_port);
   M1_1_10_0 : MUX2_X1 port map( A => MR_int_1_10_port, B => MR_int_1_12_port, 
                           S => n7, Z => MR_int_2_10_port);
   M1_1_9_0 : MUX2_X1 port map( A => MR_int_1_9_port, B => MR_int_1_11_port, S 
                           => n7, Z => MR_int_2_9_port);
   M1_1_8_0 : MUX2_X1 port map( A => MR_int_1_8_port, B => MR_int_1_10_port, S 
                           => n7, Z => MR_int_2_8_port);
   M1_1_7_0 : MUX2_X1 port map( A => MR_int_1_7_port, B => MR_int_1_9_port, S 
                           => n7, Z => MR_int_2_7_port);
   M1_1_6_0 : MUX2_X1 port map( A => MR_int_1_6_port, B => MR_int_1_8_port, S 
                           => n7, Z => MR_int_2_6_port);
   M1_1_5_0 : MUX2_X1 port map( A => MR_int_1_5_port, B => MR_int_1_7_port, S 
                           => n7, Z => MR_int_2_5_port);
   M1_1_4_0 : MUX2_X1 port map( A => MR_int_1_4_port, B => MR_int_1_6_port, S 
                           => n7, Z => MR_int_2_4_port);
   M1_1_3_0 : MUX2_X1 port map( A => MR_int_1_3_port, B => MR_int_1_5_port, S 
                           => n7, Z => MR_int_2_3_port);
   M1_1_2_0 : MUX2_X1 port map( A => MR_int_1_2_port, B => MR_int_1_4_port, S 
                           => n7, Z => MR_int_2_2_port);
   M1_1_1 : MUX2_X1 port map( A => MR_int_1_1_port, B => MR_int_1_3_port, S => 
                           n7, Z => MR_int_2_1_port);
   M1_1_0 : MUX2_X1 port map( A => MR_int_1_0_port, B => MR_int_1_2_port, S => 
                           n7, Z => MR_int_2_0_port);
   M1_0_31_0 : MUX2_X1 port map( A => A(31), B => A(0), S => n6, Z => 
                           MR_int_1_31_port);
   M1_0_30_0 : MUX2_X1 port map( A => A(30), B => A(31), S => n6, Z => 
                           MR_int_1_30_port);
   M1_0_29_0 : MUX2_X1 port map( A => A(29), B => A(30), S => n6, Z => 
                           MR_int_1_29_port);
   M1_0_28_0 : MUX2_X1 port map( A => A(28), B => A(29), S => n6, Z => 
                           MR_int_1_28_port);
   M1_0_27_0 : MUX2_X1 port map( A => A(27), B => A(28), S => n6, Z => 
                           MR_int_1_27_port);
   M1_0_26_0 : MUX2_X1 port map( A => A(26), B => A(27), S => n6, Z => 
                           MR_int_1_26_port);
   M1_0_25_0 : MUX2_X1 port map( A => A(25), B => A(26), S => n6, Z => 
                           MR_int_1_25_port);
   M1_0_24_0 : MUX2_X1 port map( A => A(24), B => A(25), S => n6, Z => 
                           MR_int_1_24_port);
   M1_0_23_0 : MUX2_X1 port map( A => A(23), B => A(24), S => n5, Z => 
                           MR_int_1_23_port);
   M1_0_22_0 : MUX2_X1 port map( A => A(22), B => A(23), S => n5, Z => 
                           MR_int_1_22_port);
   M1_0_21_0 : MUX2_X1 port map( A => A(21), B => A(22), S => n5, Z => 
                           MR_int_1_21_port);
   M1_0_20_0 : MUX2_X1 port map( A => A(20), B => A(21), S => n5, Z => 
                           MR_int_1_20_port);
   M1_0_19_0 : MUX2_X1 port map( A => A(19), B => A(20), S => n5, Z => 
                           MR_int_1_19_port);
   M1_0_18_0 : MUX2_X1 port map( A => A(18), B => A(19), S => n5, Z => 
                           MR_int_1_18_port);
   M1_0_17_0 : MUX2_X1 port map( A => A(17), B => A(18), S => n5, Z => 
                           MR_int_1_17_port);
   M1_0_16_0 : MUX2_X1 port map( A => A(16), B => A(17), S => n5, Z => 
                           MR_int_1_16_port);
   M1_0_15_0 : MUX2_X1 port map( A => A(15), B => A(16), S => n5, Z => 
                           MR_int_1_15_port);
   M1_0_14_0 : MUX2_X1 port map( A => A(14), B => A(15), S => n5, Z => 
                           MR_int_1_14_port);
   M1_0_13_0 : MUX2_X1 port map( A => A(13), B => A(14), S => n5, Z => 
                           MR_int_1_13_port);
   M1_0_12_0 : MUX2_X1 port map( A => A(12), B => A(13), S => n5, Z => 
                           MR_int_1_12_port);
   M1_0_11_0 : MUX2_X1 port map( A => A(11), B => A(12), S => n4, Z => 
                           MR_int_1_11_port);
   M1_0_10_0 : MUX2_X1 port map( A => A(10), B => A(11), S => n4, Z => 
                           MR_int_1_10_port);
   M1_0_9_0 : MUX2_X1 port map( A => A(9), B => A(10), S => n4, Z => 
                           MR_int_1_9_port);
   M1_0_8_0 : MUX2_X1 port map( A => A(8), B => A(9), S => n4, Z => 
                           MR_int_1_8_port);
   M1_0_7_0 : MUX2_X1 port map( A => A(7), B => A(8), S => n4, Z => 
                           MR_int_1_7_port);
   M1_0_6_0 : MUX2_X1 port map( A => A(6), B => A(7), S => n4, Z => 
                           MR_int_1_6_port);
   M1_0_5_0 : MUX2_X1 port map( A => A(5), B => A(6), S => n4, Z => 
                           MR_int_1_5_port);
   M1_0_4_0 : MUX2_X1 port map( A => A(4), B => A(5), S => n4, Z => 
                           MR_int_1_4_port);
   M1_0_3_0 : MUX2_X1 port map( A => A(3), B => A(4), S => n4, Z => 
                           MR_int_1_3_port);
   M1_0_2_0 : MUX2_X1 port map( A => A(2), B => A(3), S => n4, Z => 
                           MR_int_1_2_port);
   M1_0_1_0 : MUX2_X1 port map( A => A(1), B => A(2), S => n4, Z => 
                           MR_int_1_1_port);
   M1_0_0 : MUX2_X1 port map( A => A(0), B => A(1), S => n4, Z => 
                           MR_int_1_0_port);
   U2 : BUF_X1 port map( A => SH(0), Z => n4);
   U3 : BUF_X1 port map( A => SH(0), Z => n5);
   U4 : BUF_X1 port map( A => SH(1), Z => n7);
   U5 : BUF_X1 port map( A => SH(1), Z => n8);
   U6 : BUF_X1 port map( A => SH(2), Z => n10);
   U7 : BUF_X1 port map( A => SH(2), Z => n11);
   U8 : BUF_X1 port map( A => SH(0), Z => n6);
   U9 : BUF_X1 port map( A => SH(1), Z => n9);
   U10 : BUF_X1 port map( A => SH(2), Z => n12);
   U11 : BUF_X1 port map( A => SH(3), Z => n13);
   U12 : BUF_X1 port map( A => SH(3), Z => n14);
   U13 : BUF_X1 port map( A => SH(4), Z => n16);
   U14 : BUF_X1 port map( A => SH(4), Z => n17);
   U15 : BUF_X1 port map( A => SH(3), Z => n15);
   U16 : BUF_X1 port map( A => SH(4), Z => n18);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Shifter_DATA_SIZE32_DW_lbsh_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end Shifter_DATA_SIZE32_DW_lbsh_0;

architecture SYN_mx2 of Shifter_DATA_SIZE32_DW_lbsh_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal ML_int_1_31_port, ML_int_1_30_port, ML_int_1_29_port, 
      ML_int_1_28_port, ML_int_1_27_port, ML_int_1_26_port, ML_int_1_25_port, 
      ML_int_1_24_port, ML_int_1_23_port, ML_int_1_22_port, ML_int_1_21_port, 
      ML_int_1_20_port, ML_int_1_19_port, ML_int_1_18_port, ML_int_1_17_port, 
      ML_int_1_16_port, ML_int_1_15_port, ML_int_1_14_port, ML_int_1_13_port, 
      ML_int_1_12_port, ML_int_1_11_port, ML_int_1_10_port, ML_int_1_9_port, 
      ML_int_1_8_port, ML_int_1_7_port, ML_int_1_6_port, ML_int_1_5_port, 
      ML_int_1_4_port, ML_int_1_3_port, ML_int_1_2_port, ML_int_1_1_port, 
      ML_int_1_0_port, ML_int_2_31_port, ML_int_2_30_port, ML_int_2_29_port, 
      ML_int_2_28_port, ML_int_2_27_port, ML_int_2_26_port, ML_int_2_25_port, 
      ML_int_2_24_port, ML_int_2_23_port, ML_int_2_22_port, ML_int_2_21_port, 
      ML_int_2_20_port, ML_int_2_19_port, ML_int_2_18_port, ML_int_2_17_port, 
      ML_int_2_16_port, ML_int_2_15_port, ML_int_2_14_port, ML_int_2_13_port, 
      ML_int_2_12_port, ML_int_2_11_port, ML_int_2_10_port, ML_int_2_9_port, 
      ML_int_2_8_port, ML_int_2_7_port, ML_int_2_6_port, ML_int_2_5_port, 
      ML_int_2_4_port, ML_int_2_3_port, ML_int_2_2_port, ML_int_2_1_port, 
      ML_int_2_0_port, ML_int_3_31_port, ML_int_3_30_port, ML_int_3_29_port, 
      ML_int_3_28_port, ML_int_3_27_port, ML_int_3_26_port, ML_int_3_25_port, 
      ML_int_3_24_port, ML_int_3_23_port, ML_int_3_22_port, ML_int_3_21_port, 
      ML_int_3_20_port, ML_int_3_19_port, ML_int_3_18_port, ML_int_3_17_port, 
      ML_int_3_16_port, ML_int_3_15_port, ML_int_3_14_port, ML_int_3_13_port, 
      ML_int_3_12_port, ML_int_3_11_port, ML_int_3_10_port, ML_int_3_9_port, 
      ML_int_3_8_port, ML_int_3_7_port, ML_int_3_6_port, ML_int_3_5_port, 
      ML_int_3_4_port, ML_int_3_3_port, ML_int_3_2_port, ML_int_3_1_port, 
      ML_int_3_0_port, ML_int_4_31_port, ML_int_4_30_port, ML_int_4_29_port, 
      ML_int_4_28_port, ML_int_4_27_port, ML_int_4_26_port, ML_int_4_25_port, 
      ML_int_4_24_port, ML_int_4_23_port, ML_int_4_22_port, ML_int_4_21_port, 
      ML_int_4_20_port, ML_int_4_19_port, ML_int_4_18_port, ML_int_4_17_port, 
      ML_int_4_16_port, ML_int_4_15_port, ML_int_4_14_port, ML_int_4_13_port, 
      ML_int_4_12_port, ML_int_4_11_port, ML_int_4_10_port, ML_int_4_9_port, 
      ML_int_4_8_port, ML_int_4_7_port, ML_int_4_6_port, ML_int_4_5_port, 
      ML_int_4_4_port, ML_int_4_3_port, ML_int_4_2_port, ML_int_4_1_port, 
      ML_int_4_0_port, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, 
      n16, n17, n18 : std_logic;

begin
   
   M1_4_31 : MUX2_X1 port map( A => ML_int_4_31_port, B => ML_int_4_15_port, S 
                           => n18, Z => B(31));
   M1_4_30 : MUX2_X1 port map( A => ML_int_4_30_port, B => ML_int_4_14_port, S 
                           => n18, Z => B(30));
   M1_4_29 : MUX2_X1 port map( A => ML_int_4_29_port, B => ML_int_4_13_port, S 
                           => n18, Z => B(29));
   M1_4_28 : MUX2_X1 port map( A => ML_int_4_28_port, B => ML_int_4_12_port, S 
                           => n18, Z => B(28));
   M1_4_27 : MUX2_X1 port map( A => ML_int_4_27_port, B => ML_int_4_11_port, S 
                           => n18, Z => B(27));
   M1_4_26 : MUX2_X1 port map( A => ML_int_4_26_port, B => ML_int_4_10_port, S 
                           => n18, Z => B(26));
   M1_4_25 : MUX2_X1 port map( A => ML_int_4_25_port, B => ML_int_4_9_port, S 
                           => n18, Z => B(25));
   M1_4_24 : MUX2_X1 port map( A => ML_int_4_24_port, B => ML_int_4_8_port, S 
                           => n18, Z => B(24));
   M1_4_23 : MUX2_X1 port map( A => ML_int_4_23_port, B => ML_int_4_7_port, S 
                           => n17, Z => B(23));
   M1_4_22 : MUX2_X1 port map( A => ML_int_4_22_port, B => ML_int_4_6_port, S 
                           => n17, Z => B(22));
   M1_4_21 : MUX2_X1 port map( A => ML_int_4_21_port, B => ML_int_4_5_port, S 
                           => n17, Z => B(21));
   M1_4_20 : MUX2_X1 port map( A => ML_int_4_20_port, B => ML_int_4_4_port, S 
                           => n17, Z => B(20));
   M1_4_19 : MUX2_X1 port map( A => ML_int_4_19_port, B => ML_int_4_3_port, S 
                           => n17, Z => B(19));
   M1_4_18 : MUX2_X1 port map( A => ML_int_4_18_port, B => ML_int_4_2_port, S 
                           => n17, Z => B(18));
   M1_4_17 : MUX2_X1 port map( A => ML_int_4_17_port, B => ML_int_4_1_port, S 
                           => n17, Z => B(17));
   M1_4_16 : MUX2_X1 port map( A => ML_int_4_16_port, B => ML_int_4_0_port, S 
                           => n17, Z => B(16));
   M0_4_15 : MUX2_X1 port map( A => ML_int_4_15_port, B => ML_int_4_31_port, S 
                           => n17, Z => B(15));
   M0_4_14 : MUX2_X1 port map( A => ML_int_4_14_port, B => ML_int_4_30_port, S 
                           => n17, Z => B(14));
   M0_4_13 : MUX2_X1 port map( A => ML_int_4_13_port, B => ML_int_4_29_port, S 
                           => n17, Z => B(13));
   M0_4_12 : MUX2_X1 port map( A => ML_int_4_12_port, B => ML_int_4_28_port, S 
                           => n17, Z => B(12));
   M0_4_11 : MUX2_X1 port map( A => ML_int_4_11_port, B => ML_int_4_27_port, S 
                           => n16, Z => B(11));
   M0_4_10 : MUX2_X1 port map( A => ML_int_4_10_port, B => ML_int_4_26_port, S 
                           => n16, Z => B(10));
   M0_4_9 : MUX2_X1 port map( A => ML_int_4_9_port, B => ML_int_4_25_port, S =>
                           n16, Z => B(9));
   M0_4_8 : MUX2_X1 port map( A => ML_int_4_8_port, B => ML_int_4_24_port, S =>
                           n16, Z => B(8));
   M0_4_7 : MUX2_X1 port map( A => ML_int_4_7_port, B => ML_int_4_23_port, S =>
                           n16, Z => B(7));
   M0_4_6 : MUX2_X1 port map( A => ML_int_4_6_port, B => ML_int_4_22_port, S =>
                           n16, Z => B(6));
   M0_4_5 : MUX2_X1 port map( A => ML_int_4_5_port, B => ML_int_4_21_port, S =>
                           n16, Z => B(5));
   M0_4_4 : MUX2_X1 port map( A => ML_int_4_4_port, B => ML_int_4_20_port, S =>
                           n16, Z => B(4));
   M0_4_3 : MUX2_X1 port map( A => ML_int_4_3_port, B => ML_int_4_19_port, S =>
                           n16, Z => B(3));
   M0_4_2 : MUX2_X1 port map( A => ML_int_4_2_port, B => ML_int_4_18_port, S =>
                           n16, Z => B(2));
   M0_4_1 : MUX2_X1 port map( A => ML_int_4_1_port, B => ML_int_4_17_port, S =>
                           n16, Z => B(1));
   M0_4_0 : MUX2_X1 port map( A => ML_int_4_0_port, B => ML_int_4_16_port, S =>
                           n16, Z => B(0));
   M1_3_31 : MUX2_X1 port map( A => ML_int_3_31_port, B => ML_int_3_23_port, S 
                           => n15, Z => ML_int_4_31_port);
   M1_3_30 : MUX2_X1 port map( A => ML_int_3_30_port, B => ML_int_3_22_port, S 
                           => n15, Z => ML_int_4_30_port);
   M1_3_29 : MUX2_X1 port map( A => ML_int_3_29_port, B => ML_int_3_21_port, S 
                           => n15, Z => ML_int_4_29_port);
   M1_3_28 : MUX2_X1 port map( A => ML_int_3_28_port, B => ML_int_3_20_port, S 
                           => n15, Z => ML_int_4_28_port);
   M1_3_27 : MUX2_X1 port map( A => ML_int_3_27_port, B => ML_int_3_19_port, S 
                           => n15, Z => ML_int_4_27_port);
   M1_3_26 : MUX2_X1 port map( A => ML_int_3_26_port, B => ML_int_3_18_port, S 
                           => n15, Z => ML_int_4_26_port);
   M1_3_25 : MUX2_X1 port map( A => ML_int_3_25_port, B => ML_int_3_17_port, S 
                           => n15, Z => ML_int_4_25_port);
   M1_3_24 : MUX2_X1 port map( A => ML_int_3_24_port, B => ML_int_3_16_port, S 
                           => n15, Z => ML_int_4_24_port);
   M1_3_23 : MUX2_X1 port map( A => ML_int_3_23_port, B => ML_int_3_15_port, S 
                           => n14, Z => ML_int_4_23_port);
   M1_3_22 : MUX2_X1 port map( A => ML_int_3_22_port, B => ML_int_3_14_port, S 
                           => n14, Z => ML_int_4_22_port);
   M1_3_21 : MUX2_X1 port map( A => ML_int_3_21_port, B => ML_int_3_13_port, S 
                           => n14, Z => ML_int_4_21_port);
   M1_3_20 : MUX2_X1 port map( A => ML_int_3_20_port, B => ML_int_3_12_port, S 
                           => n14, Z => ML_int_4_20_port);
   M1_3_19 : MUX2_X1 port map( A => ML_int_3_19_port, B => ML_int_3_11_port, S 
                           => n14, Z => ML_int_4_19_port);
   M1_3_18 : MUX2_X1 port map( A => ML_int_3_18_port, B => ML_int_3_10_port, S 
                           => n14, Z => ML_int_4_18_port);
   M1_3_17 : MUX2_X1 port map( A => ML_int_3_17_port, B => ML_int_3_9_port, S 
                           => n14, Z => ML_int_4_17_port);
   M1_3_16 : MUX2_X1 port map( A => ML_int_3_16_port, B => ML_int_3_8_port, S 
                           => n14, Z => ML_int_4_16_port);
   M1_3_15 : MUX2_X1 port map( A => ML_int_3_15_port, B => ML_int_3_7_port, S 
                           => n14, Z => ML_int_4_15_port);
   M1_3_14 : MUX2_X1 port map( A => ML_int_3_14_port, B => ML_int_3_6_port, S 
                           => n14, Z => ML_int_4_14_port);
   M1_3_13 : MUX2_X1 port map( A => ML_int_3_13_port, B => ML_int_3_5_port, S 
                           => n14, Z => ML_int_4_13_port);
   M1_3_12 : MUX2_X1 port map( A => ML_int_3_12_port, B => ML_int_3_4_port, S 
                           => n14, Z => ML_int_4_12_port);
   M1_3_11 : MUX2_X1 port map( A => ML_int_3_11_port, B => ML_int_3_3_port, S 
                           => n13, Z => ML_int_4_11_port);
   M1_3_10 : MUX2_X1 port map( A => ML_int_3_10_port, B => ML_int_3_2_port, S 
                           => n13, Z => ML_int_4_10_port);
   M1_3_9 : MUX2_X1 port map( A => ML_int_3_9_port, B => ML_int_3_1_port, S => 
                           n13, Z => ML_int_4_9_port);
   M1_3_8 : MUX2_X1 port map( A => ML_int_3_8_port, B => ML_int_3_0_port, S => 
                           n13, Z => ML_int_4_8_port);
   M0_3_7 : MUX2_X1 port map( A => ML_int_3_7_port, B => ML_int_3_31_port, S =>
                           n13, Z => ML_int_4_7_port);
   M0_3_6 : MUX2_X1 port map( A => ML_int_3_6_port, B => ML_int_3_30_port, S =>
                           n13, Z => ML_int_4_6_port);
   M0_3_5 : MUX2_X1 port map( A => ML_int_3_5_port, B => ML_int_3_29_port, S =>
                           n13, Z => ML_int_4_5_port);
   M0_3_4 : MUX2_X1 port map( A => ML_int_3_4_port, B => ML_int_3_28_port, S =>
                           n13, Z => ML_int_4_4_port);
   M0_3_3 : MUX2_X1 port map( A => ML_int_3_3_port, B => ML_int_3_27_port, S =>
                           n13, Z => ML_int_4_3_port);
   M0_3_2 : MUX2_X1 port map( A => ML_int_3_2_port, B => ML_int_3_26_port, S =>
                           n13, Z => ML_int_4_2_port);
   M0_3_1 : MUX2_X1 port map( A => ML_int_3_1_port, B => ML_int_3_25_port, S =>
                           n13, Z => ML_int_4_1_port);
   M0_3_0 : MUX2_X1 port map( A => ML_int_3_0_port, B => ML_int_3_24_port, S =>
                           n13, Z => ML_int_4_0_port);
   M1_2_31 : MUX2_X1 port map( A => ML_int_2_31_port, B => ML_int_2_27_port, S 
                           => n12, Z => ML_int_3_31_port);
   M1_2_30 : MUX2_X1 port map( A => ML_int_2_30_port, B => ML_int_2_26_port, S 
                           => n12, Z => ML_int_3_30_port);
   M1_2_29 : MUX2_X1 port map( A => ML_int_2_29_port, B => ML_int_2_25_port, S 
                           => n12, Z => ML_int_3_29_port);
   M1_2_28 : MUX2_X1 port map( A => ML_int_2_28_port, B => ML_int_2_24_port, S 
                           => n12, Z => ML_int_3_28_port);
   M1_2_27 : MUX2_X1 port map( A => ML_int_2_27_port, B => ML_int_2_23_port, S 
                           => n12, Z => ML_int_3_27_port);
   M1_2_26 : MUX2_X1 port map( A => ML_int_2_26_port, B => ML_int_2_22_port, S 
                           => n12, Z => ML_int_3_26_port);
   M1_2_25 : MUX2_X1 port map( A => ML_int_2_25_port, B => ML_int_2_21_port, S 
                           => n12, Z => ML_int_3_25_port);
   M1_2_24 : MUX2_X1 port map( A => ML_int_2_24_port, B => ML_int_2_20_port, S 
                           => n12, Z => ML_int_3_24_port);
   M1_2_23 : MUX2_X1 port map( A => ML_int_2_23_port, B => ML_int_2_19_port, S 
                           => n11, Z => ML_int_3_23_port);
   M1_2_22 : MUX2_X1 port map( A => ML_int_2_22_port, B => ML_int_2_18_port, S 
                           => n11, Z => ML_int_3_22_port);
   M1_2_21 : MUX2_X1 port map( A => ML_int_2_21_port, B => ML_int_2_17_port, S 
                           => n11, Z => ML_int_3_21_port);
   M1_2_20 : MUX2_X1 port map( A => ML_int_2_20_port, B => ML_int_2_16_port, S 
                           => n11, Z => ML_int_3_20_port);
   M1_2_19 : MUX2_X1 port map( A => ML_int_2_19_port, B => ML_int_2_15_port, S 
                           => n11, Z => ML_int_3_19_port);
   M1_2_18 : MUX2_X1 port map( A => ML_int_2_18_port, B => ML_int_2_14_port, S 
                           => n11, Z => ML_int_3_18_port);
   M1_2_17 : MUX2_X1 port map( A => ML_int_2_17_port, B => ML_int_2_13_port, S 
                           => n11, Z => ML_int_3_17_port);
   M1_2_16 : MUX2_X1 port map( A => ML_int_2_16_port, B => ML_int_2_12_port, S 
                           => n11, Z => ML_int_3_16_port);
   M1_2_15 : MUX2_X1 port map( A => ML_int_2_15_port, B => ML_int_2_11_port, S 
                           => n11, Z => ML_int_3_15_port);
   M1_2_14 : MUX2_X1 port map( A => ML_int_2_14_port, B => ML_int_2_10_port, S 
                           => n11, Z => ML_int_3_14_port);
   M1_2_13 : MUX2_X1 port map( A => ML_int_2_13_port, B => ML_int_2_9_port, S 
                           => n11, Z => ML_int_3_13_port);
   M1_2_12 : MUX2_X1 port map( A => ML_int_2_12_port, B => ML_int_2_8_port, S 
                           => n11, Z => ML_int_3_12_port);
   M1_2_11 : MUX2_X1 port map( A => ML_int_2_11_port, B => ML_int_2_7_port, S 
                           => n10, Z => ML_int_3_11_port);
   M1_2_10 : MUX2_X1 port map( A => ML_int_2_10_port, B => ML_int_2_6_port, S 
                           => n10, Z => ML_int_3_10_port);
   M1_2_9 : MUX2_X1 port map( A => ML_int_2_9_port, B => ML_int_2_5_port, S => 
                           n10, Z => ML_int_3_9_port);
   M1_2_8 : MUX2_X1 port map( A => ML_int_2_8_port, B => ML_int_2_4_port, S => 
                           n10, Z => ML_int_3_8_port);
   M1_2_7 : MUX2_X1 port map( A => ML_int_2_7_port, B => ML_int_2_3_port, S => 
                           n10, Z => ML_int_3_7_port);
   M1_2_6 : MUX2_X1 port map( A => ML_int_2_6_port, B => ML_int_2_2_port, S => 
                           n10, Z => ML_int_3_6_port);
   M1_2_5 : MUX2_X1 port map( A => ML_int_2_5_port, B => ML_int_2_1_port, S => 
                           n10, Z => ML_int_3_5_port);
   M1_2_4 : MUX2_X1 port map( A => ML_int_2_4_port, B => ML_int_2_0_port, S => 
                           n10, Z => ML_int_3_4_port);
   M0_2_3 : MUX2_X1 port map( A => ML_int_2_3_port, B => ML_int_2_31_port, S =>
                           n10, Z => ML_int_3_3_port);
   M0_2_2 : MUX2_X1 port map( A => ML_int_2_2_port, B => ML_int_2_30_port, S =>
                           n10, Z => ML_int_3_2_port);
   M0_2_1 : MUX2_X1 port map( A => ML_int_2_1_port, B => ML_int_2_29_port, S =>
                           n10, Z => ML_int_3_1_port);
   M0_2_0 : MUX2_X1 port map( A => ML_int_2_0_port, B => ML_int_2_28_port, S =>
                           n10, Z => ML_int_3_0_port);
   M1_1_31 : MUX2_X1 port map( A => ML_int_1_31_port, B => ML_int_1_29_port, S 
                           => n9, Z => ML_int_2_31_port);
   M1_1_30 : MUX2_X1 port map( A => ML_int_1_30_port, B => ML_int_1_28_port, S 
                           => n9, Z => ML_int_2_30_port);
   M1_1_29 : MUX2_X1 port map( A => ML_int_1_29_port, B => ML_int_1_27_port, S 
                           => n9, Z => ML_int_2_29_port);
   M1_1_28 : MUX2_X1 port map( A => ML_int_1_28_port, B => ML_int_1_26_port, S 
                           => n9, Z => ML_int_2_28_port);
   M1_1_27 : MUX2_X1 port map( A => ML_int_1_27_port, B => ML_int_1_25_port, S 
                           => n9, Z => ML_int_2_27_port);
   M1_1_26 : MUX2_X1 port map( A => ML_int_1_26_port, B => ML_int_1_24_port, S 
                           => n9, Z => ML_int_2_26_port);
   M1_1_25 : MUX2_X1 port map( A => ML_int_1_25_port, B => ML_int_1_23_port, S 
                           => n9, Z => ML_int_2_25_port);
   M1_1_24 : MUX2_X1 port map( A => ML_int_1_24_port, B => ML_int_1_22_port, S 
                           => n9, Z => ML_int_2_24_port);
   M1_1_23 : MUX2_X1 port map( A => ML_int_1_23_port, B => ML_int_1_21_port, S 
                           => n8, Z => ML_int_2_23_port);
   M1_1_22 : MUX2_X1 port map( A => ML_int_1_22_port, B => ML_int_1_20_port, S 
                           => n8, Z => ML_int_2_22_port);
   M1_1_21 : MUX2_X1 port map( A => ML_int_1_21_port, B => ML_int_1_19_port, S 
                           => n8, Z => ML_int_2_21_port);
   M1_1_20 : MUX2_X1 port map( A => ML_int_1_20_port, B => ML_int_1_18_port, S 
                           => n8, Z => ML_int_2_20_port);
   M1_1_19 : MUX2_X1 port map( A => ML_int_1_19_port, B => ML_int_1_17_port, S 
                           => n8, Z => ML_int_2_19_port);
   M1_1_18 : MUX2_X1 port map( A => ML_int_1_18_port, B => ML_int_1_16_port, S 
                           => n8, Z => ML_int_2_18_port);
   M1_1_17 : MUX2_X1 port map( A => ML_int_1_17_port, B => ML_int_1_15_port, S 
                           => n8, Z => ML_int_2_17_port);
   M1_1_16 : MUX2_X1 port map( A => ML_int_1_16_port, B => ML_int_1_14_port, S 
                           => n8, Z => ML_int_2_16_port);
   M1_1_15 : MUX2_X1 port map( A => ML_int_1_15_port, B => ML_int_1_13_port, S 
                           => n8, Z => ML_int_2_15_port);
   M1_1_14 : MUX2_X1 port map( A => ML_int_1_14_port, B => ML_int_1_12_port, S 
                           => n8, Z => ML_int_2_14_port);
   M1_1_13 : MUX2_X1 port map( A => ML_int_1_13_port, B => ML_int_1_11_port, S 
                           => n8, Z => ML_int_2_13_port);
   M1_1_12 : MUX2_X1 port map( A => ML_int_1_12_port, B => ML_int_1_10_port, S 
                           => n8, Z => ML_int_2_12_port);
   M1_1_11 : MUX2_X1 port map( A => ML_int_1_11_port, B => ML_int_1_9_port, S 
                           => n7, Z => ML_int_2_11_port);
   M1_1_10 : MUX2_X1 port map( A => ML_int_1_10_port, B => ML_int_1_8_port, S 
                           => n7, Z => ML_int_2_10_port);
   M1_1_9 : MUX2_X1 port map( A => ML_int_1_9_port, B => ML_int_1_7_port, S => 
                           n7, Z => ML_int_2_9_port);
   M1_1_8 : MUX2_X1 port map( A => ML_int_1_8_port, B => ML_int_1_6_port, S => 
                           n7, Z => ML_int_2_8_port);
   M1_1_7 : MUX2_X1 port map( A => ML_int_1_7_port, B => ML_int_1_5_port, S => 
                           n7, Z => ML_int_2_7_port);
   M1_1_6 : MUX2_X1 port map( A => ML_int_1_6_port, B => ML_int_1_4_port, S => 
                           n7, Z => ML_int_2_6_port);
   M1_1_5 : MUX2_X1 port map( A => ML_int_1_5_port, B => ML_int_1_3_port, S => 
                           n7, Z => ML_int_2_5_port);
   M1_1_4 : MUX2_X1 port map( A => ML_int_1_4_port, B => ML_int_1_2_port, S => 
                           n7, Z => ML_int_2_4_port);
   M1_1_3 : MUX2_X1 port map( A => ML_int_1_3_port, B => ML_int_1_1_port, S => 
                           n7, Z => ML_int_2_3_port);
   M1_1_2 : MUX2_X1 port map( A => ML_int_1_2_port, B => ML_int_1_0_port, S => 
                           n7, Z => ML_int_2_2_port);
   M0_1_1 : MUX2_X1 port map( A => ML_int_1_1_port, B => ML_int_1_31_port, S =>
                           n7, Z => ML_int_2_1_port);
   M0_1_0 : MUX2_X1 port map( A => ML_int_1_0_port, B => ML_int_1_30_port, S =>
                           n7, Z => ML_int_2_0_port);
   M1_0_31 : MUX2_X1 port map( A => A(31), B => A(30), S => n6, Z => 
                           ML_int_1_31_port);
   M1_0_30 : MUX2_X1 port map( A => A(30), B => A(29), S => n6, Z => 
                           ML_int_1_30_port);
   M1_0_29 : MUX2_X1 port map( A => A(29), B => A(28), S => n6, Z => 
                           ML_int_1_29_port);
   M1_0_28 : MUX2_X1 port map( A => A(28), B => A(27), S => n6, Z => 
                           ML_int_1_28_port);
   M1_0_27 : MUX2_X1 port map( A => A(27), B => A(26), S => n6, Z => 
                           ML_int_1_27_port);
   M1_0_26 : MUX2_X1 port map( A => A(26), B => A(25), S => n6, Z => 
                           ML_int_1_26_port);
   M1_0_25 : MUX2_X1 port map( A => A(25), B => A(24), S => n6, Z => 
                           ML_int_1_25_port);
   M1_0_24 : MUX2_X1 port map( A => A(24), B => A(23), S => n6, Z => 
                           ML_int_1_24_port);
   M1_0_23 : MUX2_X1 port map( A => A(23), B => A(22), S => n5, Z => 
                           ML_int_1_23_port);
   M1_0_22 : MUX2_X1 port map( A => A(22), B => A(21), S => n5, Z => 
                           ML_int_1_22_port);
   M1_0_21 : MUX2_X1 port map( A => A(21), B => A(20), S => n5, Z => 
                           ML_int_1_21_port);
   M1_0_20 : MUX2_X1 port map( A => A(20), B => A(19), S => n5, Z => 
                           ML_int_1_20_port);
   M1_0_19 : MUX2_X1 port map( A => A(19), B => A(18), S => n5, Z => 
                           ML_int_1_19_port);
   M1_0_18 : MUX2_X1 port map( A => A(18), B => A(17), S => n5, Z => 
                           ML_int_1_18_port);
   M1_0_17 : MUX2_X1 port map( A => A(17), B => A(16), S => n5, Z => 
                           ML_int_1_17_port);
   M1_0_16 : MUX2_X1 port map( A => A(16), B => A(15), S => n5, Z => 
                           ML_int_1_16_port);
   M1_0_15 : MUX2_X1 port map( A => A(15), B => A(14), S => n5, Z => 
                           ML_int_1_15_port);
   M1_0_14 : MUX2_X1 port map( A => A(14), B => A(13), S => n5, Z => 
                           ML_int_1_14_port);
   M1_0_13 : MUX2_X1 port map( A => A(13), B => A(12), S => n5, Z => 
                           ML_int_1_13_port);
   M1_0_12 : MUX2_X1 port map( A => A(12), B => A(11), S => n5, Z => 
                           ML_int_1_12_port);
   M1_0_11 : MUX2_X1 port map( A => A(11), B => A(10), S => n4, Z => 
                           ML_int_1_11_port);
   M1_0_10 : MUX2_X1 port map( A => A(10), B => A(9), S => n4, Z => 
                           ML_int_1_10_port);
   M1_0_9 : MUX2_X1 port map( A => A(9), B => A(8), S => n4, Z => 
                           ML_int_1_9_port);
   M1_0_8 : MUX2_X1 port map( A => A(8), B => A(7), S => n4, Z => 
                           ML_int_1_8_port);
   M1_0_7 : MUX2_X1 port map( A => A(7), B => A(6), S => n4, Z => 
                           ML_int_1_7_port);
   M1_0_6 : MUX2_X1 port map( A => A(6), B => A(5), S => n4, Z => 
                           ML_int_1_6_port);
   M1_0_5 : MUX2_X1 port map( A => A(5), B => A(4), S => n4, Z => 
                           ML_int_1_5_port);
   M1_0_4 : MUX2_X1 port map( A => A(4), B => A(3), S => n4, Z => 
                           ML_int_1_4_port);
   M1_0_3 : MUX2_X1 port map( A => A(3), B => A(2), S => n4, Z => 
                           ML_int_1_3_port);
   M1_0_2 : MUX2_X1 port map( A => A(2), B => A(1), S => n4, Z => 
                           ML_int_1_2_port);
   M1_0_1 : MUX2_X1 port map( A => A(1), B => A(0), S => n4, Z => 
                           ML_int_1_1_port);
   M0_0_0 : MUX2_X1 port map( A => A(0), B => A(31), S => n4, Z => 
                           ML_int_1_0_port);
   U2 : BUF_X1 port map( A => SH(0), Z => n4);
   U3 : BUF_X1 port map( A => SH(0), Z => n5);
   U4 : BUF_X1 port map( A => SH(1), Z => n7);
   U5 : BUF_X1 port map( A => SH(1), Z => n8);
   U6 : BUF_X1 port map( A => SH(2), Z => n10);
   U7 : BUF_X1 port map( A => SH(2), Z => n11);
   U8 : BUF_X1 port map( A => SH(0), Z => n6);
   U9 : BUF_X1 port map( A => SH(1), Z => n9);
   U10 : BUF_X1 port map( A => SH(2), Z => n12);
   U11 : BUF_X1 port map( A => SH(3), Z => n13);
   U12 : BUF_X1 port map( A => SH(3), Z => n14);
   U13 : BUF_X1 port map( A => SH(4), Z => n16);
   U14 : BUF_X1 port map( A => SH(4), Z => n17);
   U15 : BUF_X1 port map( A => SH(3), Z => n15);
   U16 : BUF_X1 port map( A => SH(4), Z => n18);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Shifter_DATA_SIZE32_DW_sra_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end Shifter_DATA_SIZE32_DW_sra_0;

architecture SYN_mx2 of Shifter_DATA_SIZE32_DW_sra_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, B_25_port, 
      B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, B_19_port, 
      B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, B_13_port, 
      B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port, B_6_port, 
      B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, B_0_port, n2, n3, n4, 
      n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20
      , n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, 
      n35, n36, n37, n38, n39, n40, n41, n42, n43, n45, n47, n48, n49, n50, n51
      , n52, n54, n56, n57, n58, n59, n60, n61, n63, n64, n66, n67, n68, n69, 
      n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84
      , n85, n86, n87, n88, n89, n90, n91, n92, n93, n95, n96, n98, n99, n100, 
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n119, n122, n123, n124, n125, n126, n129, n130, n131, 
      n132, n133, n136, n138, n139, n140, n144, n147, n148, n149, n150, n151, 
      n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, 
      n164, n165, n166, n167, n168, n169, n172, n173, n174, n175, n176, n177, 
      n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, 
      n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, 
      n202, n203 : std_logic;

begin
   B <= ( A(31), B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, 
      B_25_port, B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, 
      B_19_port, B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, 
      B_13_port, B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port,
      B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, B_0_port );
   
   U2 : NOR2_X2 port map( A1 => SH(2), A2 => SH(3), ZN => n73);
   U142 : MUX2_X1 port map( A => A(31), B => A(30), S => n51, Z => n84);
   U3 : INV_X1 port map( A => n54, ZN => n48);
   U4 : INV_X1 port map( A => n56, ZN => n49);
   U5 : INV_X1 port map( A => n50, ZN => n43);
   U6 : INV_X1 port map( A => n51, ZN => n45);
   U7 : NAND2_X1 port map( A1 => n181, A2 => A(31), ZN => n58);
   U8 : INV_X1 port map( A => n38, ZN => n6);
   U9 : INV_X1 port map( A => n181, ZN => n177);
   U10 : INV_X1 port map( A => n3, ZN => n41);
   U11 : NOR2_X1 port map( A1 => SH(0), A2 => SH(1), ZN => n51);
   U12 : NOR2_X1 port map( A1 => n173, A2 => SH(1), ZN => n50);
   U13 : NAND2_X1 port map( A1 => SH(0), A2 => SH(1), ZN => n56);
   U14 : NAND2_X1 port map( A1 => SH(1), A2 => n173, ZN => n54);
   U15 : NAND2_X1 port map( A1 => n73, A2 => n177, ZN => n3);
   U16 : AND2_X1 port map( A1 => SH(2), A2 => n159, ZN => n10);
   U17 : AOI221_X1 port map( B1 => n50, B2 => A(7), C1 => n51, C2 => A(6), A =>
                           n64, ZN => n26);
   U18 : OAI22_X1 port map( A1 => n188, A2 => n54, B1 => n189, B2 => n56, ZN =>
                           n64);
   U19 : OAI21_X1 port map( B1 => n174, B2 => n203, A => n100, ZN => n114);
   U20 : NAND2_X1 port map( A1 => n71, A2 => n177, ZN => n38);
   U21 : NOR2_X1 port map( A1 => n100, A2 => n174, ZN => n85);
   U22 : AND2_X1 port map( A1 => n159, A2 => n174, ZN => n8);
   U23 : INV_X1 port map( A => n100, ZN => n74);
   U24 : BUF_X1 port map( A => n175, Z => n178);
   U25 : BUF_X1 port map( A => n175, Z => n179);
   U26 : BUF_X1 port map( A => n176, Z => n180);
   U27 : BUF_X1 port map( A => n176, Z => n181);
   U28 : OAI221_X1 port map( B1 => n26, B2 => n3, C1 => n27, C2 => n177, A => 
                           n28, ZN => B_6_port);
   U29 : AOI222_X1 port map( A1 => n6, A2 => n29, B1 => n8, B2 => n30, C1 => 
                           n10, C2 => n31, ZN => n28);
   U30 : OAI221_X1 port map( B1 => n20, B2 => n3, C1 => n21, C2 => n177, A => 
                           n22, ZN => B_7_port);
   U31 : AOI222_X1 port map( A1 => n6, A2 => n23, B1 => n8, B2 => n24, C1 => 
                           n10, C2 => n25, ZN => n22);
   U32 : OAI221_X1 port map( B1 => n148, B2 => n3, C1 => n69, C2 => n177, A => 
                           n149, ZN => B_10_port);
   U33 : INV_X1 port map( A => n29, ZN => n148);
   U34 : AOI222_X1 port map( A1 => n6, A2 => n30, B1 => n8, B2 => n31, C1 => 
                           n10, C2 => n80, ZN => n149);
   U35 : OAI221_X1 port map( B1 => n132, B2 => n3, C1 => n68, C2 => n177, A => 
                           n133, ZN => B_11_port);
   U36 : INV_X1 port map( A => n23, ZN => n132);
   U37 : AOI222_X1 port map( A1 => n6, A2 => n24, B1 => n8, B2 => n25, C1 => 
                           n10, C2 => n78, ZN => n133);
   U38 : OAI221_X1 port map( B1 => n35, B2 => n38, C1 => n107, C2 => n177, A =>
                           n156, ZN => B_0_port);
   U39 : AOI222_X1 port map( A1 => n10, A2 => n16, B1 => n41, B2 => n157, C1 =>
                           n8, C2 => n19, ZN => n156);
   U40 : OAI221_X1 port map( B1 => n54, B2 => n183, C1 => n56, C2 => n184, A =>
                           n160, ZN => n157);
   U41 : AOI22_X1 port map( A1 => A(1), A2 => n50, B1 => A(0), B2 => n51, ZN =>
                           n160);
   U42 : OAI221_X1 port map( B1 => n32, B2 => n38, C1 => n90, C2 => n177, A => 
                           n91, ZN => B_1_port);
   U43 : AOI222_X1 port map( A1 => n10, A2 => n7, B1 => n41, B2 => n92, C1 => 
                           n8, C2 => n12, ZN => n91);
   U44 : OAI221_X1 port map( B1 => n43, B2 => n183, C1 => n45, C2 => n182, A =>
                           n95, ZN => n92);
   U45 : OAI221_X1 port map( B1 => n26, B2 => n38, C1 => n59, C2 => n177, A => 
                           n60, ZN => B_2_port);
   U46 : AOI222_X1 port map( A1 => n10, A2 => n30, B1 => n41, B2 => n61, C1 => 
                           n8, C2 => n29, ZN => n60);
   U47 : OAI221_X1 port map( B1 => n43, B2 => n184, C1 => n45, C2 => n183, A =>
                           n63, ZN => n61);
   U48 : AOI22_X1 port map( A1 => A(4), A2 => n48, B1 => A(5), B2 => n49, ZN =>
                           n63);
   U49 : OAI221_X1 port map( B1 => n20, B2 => n38, C1 => n39, C2 => n177, A => 
                           n40, ZN => B_3_port);
   U50 : AOI222_X1 port map( A1 => n10, A2 => n24, B1 => n41, B2 => n42, C1 => 
                           n8, C2 => n23, ZN => n40);
   U51 : OAI221_X1 port map( B1 => n43, B2 => n185, C1 => n45, C2 => n184, A =>
                           n47, ZN => n42);
   U52 : AOI22_X1 port map( A1 => A(5), A2 => n48, B1 => A(6), B2 => n49, ZN =>
                           n47);
   U53 : OAI221_X1 port map( B1 => n43, B2 => n191, C1 => n45, C2 => n190, A =>
                           n155, ZN => n29);
   U54 : AOI22_X1 port map( A1 => A(12), A2 => n48, B1 => A(13), B2 => n49, ZN 
                           => n155);
   U55 : OAI221_X1 port map( B1 => n43, B2 => n201, C1 => n45, C2 => n200, A =>
                           n119, ZN => n72);
   U56 : AOI22_X1 port map( A1 => A(27), A2 => n48, B1 => A(28), B2 => n49, ZN 
                           => n119);
   U57 : OAI221_X1 port map( B1 => n43, B2 => n192, C1 => n45, C2 => n191, A =>
                           n147, ZN => n23);
   U58 : AOI22_X1 port map( A1 => A(13), A2 => n48, B1 => A(14), B2 => n49, ZN 
                           => n147);
   U59 : OAI221_X1 port map( B1 => n43, B2 => n200, C1 => n45, C2 => n199, A =>
                           n164, ZN => n76);
   U60 : AOI22_X1 port map( A1 => A(26), A2 => n48, B1 => A(27), B2 => n49, ZN 
                           => n164);
   U61 : OAI221_X1 port map( B1 => n43, B2 => n190, C1 => n45, C2 => n189, A =>
                           n93, ZN => n12);
   U62 : AOI22_X1 port map( A1 => A(11), A2 => n48, B1 => A(12), B2 => n49, ZN 
                           => n93);
   U63 : OAI221_X1 port map( B1 => n43, B2 => n193, C1 => n45, C2 => n192, A =>
                           n161, ZN => n16);
   U64 : AOI22_X1 port map( A1 => A(14), A2 => n48, B1 => A(15), B2 => n49, ZN 
                           => n161);
   U65 : OAI221_X1 port map( B1 => n43, B2 => n194, C1 => n45, C2 => n193, A =>
                           n129, ZN => n7);
   U66 : AOI22_X1 port map( A1 => A(15), A2 => n48, B1 => A(16), B2 => n49, ZN 
                           => n129);
   U67 : OAI221_X1 port map( B1 => n43, B2 => n196, C1 => n195, C2 => n45, A =>
                           n168, ZN => n18);
   U68 : AOI22_X1 port map( A1 => A(22), A2 => n48, B1 => A(23), B2 => n49, ZN 
                           => n168);
   U69 : OAI221_X1 port map( B1 => n43, B2 => n197, C1 => n45, C2 => n196, A =>
                           n122, ZN => n11);
   U70 : AOI22_X1 port map( A1 => A(23), A2 => n48, B1 => A(24), B2 => n49, ZN 
                           => n122);
   U71 : OAI221_X1 port map( B1 => n43, B2 => n198, C1 => n45, C2 => n197, A =>
                           n150, ZN => n80);
   U72 : AOI22_X1 port map( A1 => A(24), A2 => n48, B1 => A(25), B2 => n49, ZN 
                           => n150);
   U73 : OAI221_X1 port map( B1 => n43, B2 => n199, C1 => n45, C2 => n198, A =>
                           n136, ZN => n78);
   U74 : AOI22_X1 port map( A1 => A(25), A2 => n48, B1 => A(26), B2 => n49, ZN 
                           => n136);
   U75 : OAI21_X1 port map( B1 => n178, B2 => n107, A => n58, ZN => B_16_port);
   U76 : OAI21_X1 port map( B1 => n178, B2 => n90, A => n58, ZN => B_17_port);
   U77 : OAI21_X1 port map( B1 => n178, B2 => n59, A => n58, ZN => B_18_port);
   U78 : OAI21_X1 port map( B1 => n179, B2 => n39, A => n58, ZN => B_19_port);
   U79 : OAI21_X1 port map( B1 => n178, B2 => n36, A => n58, ZN => B_20_port);
   U80 : OAI21_X1 port map( B1 => n178, B2 => n33, A => n58, ZN => B_21_port);
   U81 : OAI21_X1 port map( B1 => n179, B2 => n27, A => n58, ZN => B_22_port);
   U82 : OAI21_X1 port map( B1 => n179, B2 => n21, A => n58, ZN => B_23_port);
   U83 : OAI21_X1 port map( B1 => n179, B2 => n14, A => n58, ZN => B_24_port);
   U84 : NOR2_X1 port map( A1 => n174, A2 => SH(3), ZN => n71);
   U85 : AOI221_X1 port map( B1 => n50, B2 => A(8), C1 => n51, C2 => A(7), A =>
                           n52, ZN => n20);
   U86 : OAI22_X1 port map( A1 => n189, A2 => n54, B1 => n190, B2 => n56, ZN =>
                           n52);
   U87 : AOI221_X1 port map( B1 => n50, B2 => A(5), C1 => n51, C2 => A(4), A =>
                           n169, ZN => n35);
   U88 : OAI22_X1 port map( A1 => n186, A2 => n54, B1 => n187, B2 => n56, ZN =>
                           n169);
   U89 : AOI221_X1 port map( B1 => n50, B2 => A(6), C1 => n51, C2 => A(5), A =>
                           n96, ZN => n32);
   U90 : OAI22_X1 port map( A1 => n187, A2 => n54, B1 => n188, B2 => n56, ZN =>
                           n96);
   U91 : OAI221_X1 port map( B1 => n43, B2 => n189, C1 => n45, C2 => n188, A =>
                           n158, ZN => n19);
   U92 : AOI22_X1 port map( A1 => A(10), A2 => n48, B1 => A(11), B2 => n49, ZN 
                           => n158);
   U93 : AND2_X1 port map( A1 => SH(3), A2 => n174, ZN => n83);
   U94 : AOI22_X1 port map( A1 => A(3), A2 => n48, B1 => A(4), B2 => n49, ZN =>
                           n95);
   U95 : NAND2_X1 port map( A1 => A(31), A2 => SH(3), ZN => n100);
   U96 : OAI21_X1 port map( B1 => n179, B2 => n4, A => n58, ZN => B_25_port);
   U97 : OAI21_X1 port map( B1 => n180, B2 => n69, A => n58, ZN => B_26_port);
   U98 : OAI21_X1 port map( B1 => n180, B2 => n68, A => n58, ZN => B_27_port);
   U99 : OAI21_X1 port map( B1 => n180, B2 => n67, A => n58, ZN => B_28_port);
   U100 : OAI21_X1 port map( B1 => n180, B2 => n66, A => n58, ZN => B_29_port);
   U101 : OAI21_X1 port map( B1 => n180, B2 => n57, A => n58, ZN => B_30_port);
   U102 : INV_X1 port map( A => n109, ZN => n24);
   U103 : AND2_X1 port map( A1 => SH(2), A2 => SH(3), ZN => n104);
   U104 : AND2_X1 port map( A1 => SH(3), A2 => n177, ZN => n159);
   U105 : BUF_X1 port map( A => SH(4), Z => n176);
   U106 : BUF_X1 port map( A => SH(4), Z => n175);
   U107 : INV_X1 port map( A => A(7), ZN => n187);
   U108 : AOI221_X1 port map( B1 => n77, B2 => n71, C1 => n78, C2 => n73, A => 
                           n74, ZN => n21);
   U109 : AOI221_X1 port map( B1 => n75, B2 => n71, C1 => n76, C2 => n73, A => 
                           n74, ZN => n14);
   U110 : AOI221_X1 port map( B1 => n72, B2 => n71, C1 => n11, C2 => n73, A => 
                           n86, ZN => n33);
   U111 : INV_X1 port map( A => n87, ZN => n86);
   U112 : AOI21_X1 port map( B1 => n83, B2 => n70, A => n85, ZN => n87);
   U113 : AOI221_X1 port map( B1 => n79, B2 => n71, C1 => n80, C2 => n73, A => 
                           n81, ZN => n27);
   U114 : INV_X1 port map( A => n82, ZN => n81);
   U115 : AOI21_X1 port map( B1 => n83, B2 => n84, A => n85, ZN => n82);
   U116 : OAI221_X1 port map( B1 => n13, B2 => n3, C1 => n14, C2 => n177, A => 
                           n15, ZN => B_8_port);
   U117 : INV_X1 port map( A => n19, ZN => n13);
   U118 : AOI222_X1 port map( A1 => n6, A2 => n16, B1 => n8, B2 => n17, C1 => 
                           n10, C2 => n18, ZN => n15);
   U119 : OAI221_X1 port map( B1 => n32, B2 => n3, C1 => n33, C2 => n177, A => 
                           n34, ZN => B_5_port);
   U120 : AOI222_X1 port map( A1 => n6, A2 => n12, B1 => n8, B2 => n7, C1 => 
                           n10, C2 => n9, ZN => n34);
   U121 : OAI221_X1 port map( B1 => n115, B2 => n3, C1 => n66, C2 => n177, A =>
                           n116, ZN => B_13_port);
   U122 : INV_X1 port map( A => n7, ZN => n115);
   U123 : AOI222_X1 port map( A1 => n6, A2 => n9, B1 => n8, B2 => n11, C1 => 
                           n10, C2 => n72, ZN => n116);
   U124 : OAI221_X1 port map( B1 => n112, B2 => n3, C1 => n57, C2 => n177, A =>
                           n113, ZN => B_14_port);
   U125 : AOI222_X1 port map( A1 => n6, A2 => n31, B1 => n8, B2 => n80, C1 => 
                           n10, C2 => n79, ZN => n113);
   U126 : OAI221_X1 port map( B1 => n35, B2 => n3, C1 => n36, C2 => n177, A => 
                           n37, ZN => B_4_port);
   U127 : AOI222_X1 port map( A1 => n6, A2 => n19, B1 => n8, B2 => n16, C1 => 
                           n10, C2 => n17, ZN => n37);
   U128 : OAI221_X1 port map( B1 => n2, B2 => n3, C1 => n4, C2 => n177, A => n5
                           , ZN => B_9_port);
   U129 : INV_X1 port map( A => n12, ZN => n2);
   U130 : AOI222_X1 port map( A1 => n6, A2 => n7, B1 => n8, B2 => n9, C1 => n10
                           , C2 => n11, ZN => n5);
   U131 : OAI221_X1 port map( B1 => n130, B2 => n3, C1 => n67, C2 => n177, A =>
                           n131, ZN => B_12_port);
   U132 : INV_X1 port map( A => n16, ZN => n130);
   U133 : AOI222_X1 port map( A1 => n6, A2 => n17, B1 => n8, B2 => n18, C1 => 
                           n10, C2 => n76, ZN => n131);
   U134 : OAI221_X1 port map( B1 => n108, B2 => n38, C1 => n109, C2 => n3, A =>
                           n110, ZN => B_15_port);
   U135 : INV_X1 port map( A => n25, ZN => n108);
   U136 : AOI221_X1 port map( B1 => n10, B2 => n77, C1 => n8, C2 => n78, A => 
                           n111, ZN => n110);
   U137 : INV_X1 port map( A => n58, ZN => n111);
   U138 : OAI221_X1 port map( B1 => n138, B2 => n43, C1 => n123, C2 => n45, A 
                           => n151, ZN => n31);
   U139 : AOI22_X1 port map( A1 => A(20), A2 => n48, B1 => A(21), B2 => n49, ZN
                           => n151);
   U140 : OAI221_X1 port map( B1 => n195, B2 => n43, C1 => n138, C2 => n45, A 
                           => n139, ZN => n25);
   U141 : AOI22_X1 port map( A1 => A(21), A2 => n48, B1 => A(22), B2 => n49, ZN
                           => n139);
   U143 : INV_X1 port map( A => n112, ZN => n30);
   U144 : AOI221_X1 port map( B1 => n18, B2 => n71, C1 => n17, C2 => n73, A => 
                           n162, ZN => n107);
   U145 : INV_X1 port map( A => n163, ZN => n162);
   U146 : AOI22_X1 port map( A1 => n104, A2 => n75, B1 => n83, B2 => n76, ZN =>
                           n163);
   U147 : AOI221_X1 port map( B1 => n11, B2 => n71, C1 => n9, C2 => n73, A => 
                           n105, ZN => n90);
   U148 : INV_X1 port map( A => n106, ZN => n105);
   U149 : AOI22_X1 port map( A1 => n104, A2 => n70, B1 => n83, B2 => n72, ZN =>
                           n106);
   U150 : AOI221_X1 port map( B1 => n80, B2 => n71, C1 => n31, C2 => n73, A => 
                           n102, ZN => n59);
   U151 : INV_X1 port map( A => n103, ZN => n102);
   U152 : AOI22_X1 port map( A1 => n104, A2 => n84, B1 => n83, B2 => n79, ZN =>
                           n103);
   U153 : AOI221_X1 port map( B1 => n78, B2 => n71, C1 => n25, C2 => n73, A => 
                           n98, ZN => n39);
   U154 : INV_X1 port map( A => n99, ZN => n98);
   U155 : AOI21_X1 port map( B1 => n83, B2 => n77, A => n85, ZN => n99);
   U156 : AOI221_X1 port map( B1 => n76, B2 => n71, C1 => n18, C2 => n73, A => 
                           n88, ZN => n36);
   U157 : INV_X1 port map( A => n89, ZN => n88);
   U158 : AOI21_X1 port map( B1 => n83, B2 => n75, A => n85, ZN => n89);
   U159 : AOI221_X1 port map( B1 => n70, B2 => n71, C1 => n72, C2 => n73, A => 
                           n74, ZN => n4);
   U160 : AOI221_X1 port map( B1 => n84, B2 => n71, C1 => n79, C2 => n73, A => 
                           n74, ZN => n69);
   U161 : AOI221_X1 port map( B1 => n50, B2 => A(16), C1 => n51, C2 => A(15), A
                           => n140, ZN => n109);
   U162 : OAI22_X1 port map( A1 => n124, A2 => n54, B1 => n123, B2 => n56, ZN 
                           => n140);
   U163 : AOI21_X1 port map( B1 => n77, B2 => n73, A => n114, ZN => n68);
   U164 : AOI21_X1 port map( B1 => n75, B2 => n73, A => n114, ZN => n67);
   U165 : AOI21_X1 port map( B1 => n70, B2 => n73, A => n114, ZN => n66);
   U166 : AOI21_X1 port map( B1 => n84, B2 => n73, A => n114, ZN => n57);
   U167 : AOI221_X1 port map( B1 => n50, B2 => A(15), C1 => n51, C2 => A(14), A
                           => n152, ZN => n112);
   U168 : INV_X1 port map( A => n153, ZN => n152);
   U169 : AOI22_X1 port map( A1 => A(16), A2 => n48, B1 => A(17), B2 => n49, ZN
                           => n153);
   U170 : OAI221_X1 port map( B1 => n43, B2 => n123, C1 => n45, C2 => n124, A 
                           => n125, ZN => n9);
   U171 : AOI22_X1 port map( A1 => A(19), A2 => n48, B1 => A(20), B2 => n49, ZN
                           => n125);
   U172 : OAI221_X1 port map( B1 => n43, B2 => n202, C1 => n45, C2 => n201, A 
                           => n154, ZN => n79);
   U173 : AOI22_X1 port map( A1 => A(28), A2 => n48, B1 => A(29), B2 => n49, ZN
                           => n154);
   U174 : OAI221_X1 port map( B1 => n43, B2 => n172, C1 => n45, C2 => n202, A 
                           => n144, ZN => n77);
   U175 : AOI22_X1 port map( A1 => A(29), A2 => n48, B1 => A(30), B2 => n49, ZN
                           => n144);
   U176 : OAI221_X1 port map( B1 => n43, B2 => n165, C1 => n45, C2 => n172, A 
                           => n166, ZN => n75);
   U177 : INV_X1 port map( A => A(29), ZN => n165);
   U178 : AOI22_X1 port map( A1 => A(30), A2 => n48, B1 => A(31), B2 => n49, ZN
                           => n166);
   U179 : OAI221_X1 port map( B1 => n54, B2 => n123, C1 => n138, C2 => n56, A 
                           => n167, ZN => n17);
   U180 : AOI22_X1 port map( A1 => A(17), A2 => n50, B1 => A(16), B2 => n51, ZN
                           => n167);
   U181 : INV_X1 port map( A => n126, ZN => n70);
   U182 : AOI222_X1 port map( A1 => n51, A2 => A(29), B1 => n50, B2 => A(30), 
                           C1 => SH(1), C2 => A(31), ZN => n126);
   U183 : INV_X1 port map( A => A(18), ZN => n123);
   U184 : INV_X1 port map( A => A(19), ZN => n138);
   U185 : INV_X1 port map( A => A(17), ZN => n124);
   U186 : INV_X1 port map( A => A(28), ZN => n172);
   U187 : INV_X1 port map( A => SH(0), ZN => n173);
   U188 : INV_X1 port map( A => SH(2), ZN => n174);
   U189 : INV_X1 port map( A => A(1), ZN => n182);
   U190 : INV_X1 port map( A => A(2), ZN => n183);
   U191 : INV_X1 port map( A => A(3), ZN => n184);
   U192 : INV_X1 port map( A => A(4), ZN => n185);
   U193 : INV_X1 port map( A => A(6), ZN => n186);
   U194 : INV_X1 port map( A => A(8), ZN => n188);
   U195 : INV_X1 port map( A => A(9), ZN => n189);
   U196 : INV_X1 port map( A => A(10), ZN => n190);
   U197 : INV_X1 port map( A => A(11), ZN => n191);
   U198 : INV_X1 port map( A => A(12), ZN => n192);
   U199 : INV_X1 port map( A => A(13), ZN => n193);
   U200 : INV_X1 port map( A => A(14), ZN => n194);
   U201 : INV_X1 port map( A => A(20), ZN => n195);
   U202 : INV_X1 port map( A => A(21), ZN => n196);
   U203 : INV_X1 port map( A => A(22), ZN => n197);
   U204 : INV_X1 port map( A => A(23), ZN => n198);
   U205 : INV_X1 port map( A => A(24), ZN => n199);
   U206 : INV_X1 port map( A => A(25), ZN => n200);
   U207 : INV_X1 port map( A => A(26), ZN => n201);
   U208 : INV_X1 port map( A => A(27), ZN => n202);
   U209 : INV_X1 port map( A => A(31), ZN => n203);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Shifter_DATA_SIZE32_DW_rash_0 is

   port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH : 
         in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out 
         std_logic_vector (31 downto 0));

end Shifter_DATA_SIZE32_DW_rash_0;

architecture SYN_mx2 of Shifter_DATA_SIZE32_DW_rash_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, 
      n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31
      , n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n46, 
      n48, n49, n50, n51, n52, n53, n55, n57, n58, n59, n60, n61, n62, n63, n65
      , n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97
      , n98, n99, n100, n101, n102, n103, n104, n105, n108, n109, n111, n114, 
      n117, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n131, 
      n132, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, 
      n146, n147, n150, n152, n154, n155, n156, n157, n158, n160, n161, n163, 
      n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, 
      n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199 : 
      std_logic;

begin
   
   U3 : NOR2_X2 port map( A1 => SH(0), A2 => SH(1), ZN => n50);
   U4 : NOR2_X2 port map( A1 => n167, A2 => SH(1), ZN => n49);
   U102 : MUX2_X1 port map( A => n75, B => n58, S => SH(2), Z => n89);
   U5 : NOR2_X1 port map( A1 => n168, A2 => n169, ZN => n73);
   U6 : INV_X1 port map( A => n38, ZN => n6);
   U7 : INV_X1 port map( A => n3, ZN => n41);
   U8 : INV_X1 port map( A => n165, ZN => n52);
   U9 : NAND2_X1 port map( A1 => n72, A2 => n177, ZN => n3);
   U10 : NAND2_X1 port map( A1 => n73, A2 => n177, ZN => n38);
   U11 : INV_X1 port map( A => n50, ZN => n57);
   U12 : INV_X1 port map( A => n49, ZN => n55);
   U13 : INV_X1 port map( A => n44, ZN => n51);
   U14 : BUF_X1 port map( A => n46, Z => n165);
   U15 : INV_X1 port map( A => n12, ZN => n37);
   U16 : INV_X1 port map( A => n2, ZN => n33);
   U17 : INV_X1 port map( A => n174, ZN => n177);
   U18 : NOR2_X1 port map( A1 => n177, A2 => n124, ZN => n99);
   U19 : AND2_X1 port map( A1 => n147, A2 => n168, ZN => n8);
   U20 : INV_X1 port map( A => n124, ZN => n72);
   U21 : NOR3_X1 port map( A1 => n69, A2 => n171, A3 => n169, ZN => B(27));
   U22 : BUF_X1 port map( A => n46, Z => n164);
   U23 : BUF_X1 port map( A => n46, Z => n166);
   U24 : AND2_X1 port map( A1 => n41, A2 => n58, ZN => B(31));
   U25 : NAND2_X1 port map( A1 => SH(1), A2 => SH(0), ZN => n44);
   U26 : AOI221_X1 port map( B1 => n51, B2 => A(11), C1 => n52, C2 => A(10), A 
                           => n146, ZN => n12);
   U27 : OAI22_X1 port map( A1 => n185, A2 => n55, B1 => n184, B2 => n57, ZN =>
                           n146);
   U28 : AOI221_X1 port map( B1 => n51, B2 => A(12), C1 => n52, C2 => A(11), A 
                           => n83, ZN => n2);
   U29 : OAI22_X1 port map( A1 => n186, A2 => n55, B1 => n185, B2 => n57, ZN =>
                           n83);
   U30 : NOR2_X1 port map( A1 => n199, A2 => n57, ZN => n58);
   U31 : NAND2_X1 port map( A1 => SH(1), A2 => n167, ZN => n46);
   U32 : NOR2_X1 port map( A1 => n173, A2 => n39, ZN => B(19));
   U33 : NOR2_X1 port map( A1 => n174, A2 => n60, ZN => B(18));
   U34 : INV_X1 port map( A => n63, ZN => n27);
   U35 : INV_X1 port map( A => n43, ZN => n21);
   U36 : INV_X1 port map( A => n89, ZN => n69);
   U37 : AND2_X1 port map( A1 => SH(2), A2 => n147, ZN => n10);
   U38 : NOR2_X1 port map( A1 => n170, A2 => SH(2), ZN => n76);
   U39 : AOI221_X1 port map( B1 => n51, B2 => A(8), C1 => n52, C2 => A(7), A =>
                           n88, ZN => n30);
   U40 : OAI22_X1 port map( A1 => n182, A2 => n55, B1 => n181, B2 => n57, ZN =>
                           n88);
   U41 : AOI221_X1 port map( B1 => n51, B2 => A(9), C1 => n52, C2 => A(8), A =>
                           n66, ZN => n24);
   U42 : OAI22_X1 port map( A1 => n183, A2 => n55, B1 => n182, B2 => n57, ZN =>
                           n66);
   U43 : AOI221_X1 port map( B1 => n51, B2 => A(10), C1 => n52, C2 => A(9), A 
                           => n53, ZN => n18);
   U44 : OAI22_X1 port map( A1 => n184, A2 => n55, B1 => n183, B2 => n57, ZN =>
                           n53);
   U45 : NOR2_X1 port map( A1 => n168, A2 => n170, ZN => n92);
   U46 : NOR2_X1 port map( A1 => n170, A2 => n171, ZN => n147);
   U47 : NAND2_X1 port map( A1 => n168, A2 => n170, ZN => n124);
   U48 : NOR2_X1 port map( A1 => n173, A2 => n31, ZN => B(21));
   U49 : NOR2_X1 port map( A1 => n173, A2 => n25, ZN => B(22));
   U50 : NOR2_X1 port map( A1 => n172, A2 => n19, ZN => B(23));
   U51 : NOR2_X1 port map( A1 => n172, A2 => n4, ZN => B(25));
   U52 : NOR2_X1 port map( A1 => n171, A2 => n70, ZN => B(26));
   U53 : BUF_X1 port map( A => n176, Z => n171);
   U54 : BUF_X1 port map( A => n175, Z => n173);
   U55 : BUF_X1 port map( A => n176, Z => n172);
   U56 : BUF_X1 port map( A => n175, Z => n174);
   U57 : OAI221_X1 port map( B1 => n44, B2 => n198, C1 => n165, C2 => n197, A 
                           => n156, ZN => n74);
   U58 : AOI22_X1 port map( A1 => A(25), A2 => n49, B1 => A(24), B2 => n50, ZN 
                           => n156);
   U59 : OAI221_X1 port map( B1 => n44, B2 => n163, C1 => n164, C2 => n198, A 
                           => n114, ZN => n71);
   U60 : AOI22_X1 port map( A1 => A(26), A2 => n49, B1 => A(25), B2 => n50, ZN 
                           => n114);
   U61 : AOI222_X1 port map( A1 => n23, A2 => n72, B1 => n77, B2 => n73, C1 => 
                           n89, C2 => n169, ZN => n39);
   U62 : AOI221_X1 port map( B1 => n51, B2 => A(13), C1 => n52, C2 => A(12), A 
                           => n143, ZN => n63);
   U63 : OAI22_X1 port map( A1 => n187, A2 => n55, B1 => n186, B2 => n57, ZN =>
                           n143);
   U64 : AOI221_X1 port map( B1 => n51, B2 => A(14), C1 => n52, C2 => A(13), A 
                           => n132, ZN => n43);
   U65 : OAI22_X1 port map( A1 => n188, A2 => n55, B1 => n187, B2 => n57, ZN =>
                           n132);
   U66 : OAI221_X1 port map( B1 => n24, B2 => n3, C1 => n25, C2 => n177, A => 
                           n26, ZN => B(6));
   U67 : AOI222_X1 port map( A1 => n6, A2 => n27, B1 => n8, B2 => n28, C1 => 
                           n10, C2 => n29, ZN => n26);
   U68 : OAI221_X1 port map( B1 => n18, B2 => n3, C1 => n19, C2 => n177, A => 
                           n20, ZN => B(7));
   U69 : AOI222_X1 port map( A1 => n6, A2 => n21, B1 => n8, B2 => n22, C1 => 
                           n10, C2 => n23, ZN => n20);
   U70 : OAI221_X1 port map( B1 => n34, B2 => n38, C1 => n95, C2 => n177, A => 
                           n144, ZN => B(0));
   U71 : AOI222_X1 port map( A1 => n10, A2 => n15, B1 => n41, B2 => n145, C1 =>
                           n8, C2 => n37, ZN => n144);
   U72 : OAI221_X1 port map( B1 => n44, B2 => n179, C1 => n164, C2 => n178, A 
                           => n150, ZN => n145);
   U73 : AOI22_X1 port map( A1 => A(1), A2 => n49, B1 => A(0), B2 => n50, ZN =>
                           n150);
   U74 : OAI221_X1 port map( B1 => n30, B2 => n38, C1 => n80, C2 => n177, A => 
                           n81, ZN => B(1));
   U75 : AOI222_X1 port map( A1 => n10, A2 => n7, B1 => n41, B2 => n82, C1 => 
                           n8, C2 => n33, ZN => n81);
   U76 : OAI221_X1 port map( B1 => n44, B2 => n180, C1 => n166, C2 => n179, A 
                           => n87, ZN => n82);
   U77 : AOI22_X1 port map( A1 => A(2), A2 => n49, B1 => A(1), B2 => n50, ZN =>
                           n87);
   U78 : OAI221_X1 port map( B1 => n24, B2 => n38, C1 => n60, C2 => n177, A => 
                           n61, ZN => B(2));
   U79 : AOI222_X1 port map( A1 => n10, A2 => n28, B1 => n41, B2 => n62, C1 => 
                           n8, C2 => n27, ZN => n61);
   U80 : OAI221_X1 port map( B1 => n44, B2 => n181, C1 => n166, C2 => n180, A 
                           => n65, ZN => n62);
   U81 : AOI22_X1 port map( A1 => A(3), A2 => n49, B1 => A(2), B2 => n50, ZN =>
                           n65);
   U82 : OAI221_X1 port map( B1 => n18, B2 => n38, C1 => n39, C2 => n177, A => 
                           n40, ZN => B(3));
   U83 : AOI222_X1 port map( A1 => n10, A2 => n22, B1 => n41, B2 => n42, C1 => 
                           n8, C2 => n21, ZN => n40);
   U84 : OAI221_X1 port map( B1 => n44, B2 => n182, C1 => n166, C2 => n181, A 
                           => n48, ZN => n42);
   U85 : AOI22_X1 port map( A1 => A(4), A2 => n49, B1 => A(3), B2 => n50, ZN =>
                           n48);
   U86 : OAI221_X1 port map( B1 => n97, B2 => n38, C1 => n43, C2 => n3, A => 
                           n125, ZN => B(11));
   U87 : AOI221_X1 port map( B1 => n10, B2 => n77, C1 => n8, C2 => n23, A => 
                           n126, ZN => n125);
   U88 : NOR3_X1 port map( A1 => n177, A2 => n169, A3 => n69, ZN => n126);
   U89 : OAI221_X1 port map( B1 => n55, B2 => n193, C1 => n192, C2 => n57, A =>
                           n160, ZN => n17);
   U90 : AOI22_X1 port map( A1 => A(23), A2 => n51, B1 => A(22), B2 => n52, ZN 
                           => n160);
   U91 : AOI221_X1 port map( B1 => n79, B2 => n73, C1 => n29, C2 => n72, A => 
                           n90, ZN => n60);
   U92 : INV_X1 port map( A => n91, ZN => n90);
   U93 : AOI22_X1 port map( A1 => n92, A2 => n59, B1 => n76, B2 => n78, ZN => 
                           n91);
   U94 : NOR2_X1 port map( A1 => n172, A2 => n80, ZN => B(17));
   U95 : NOR2_X1 port map( A1 => n171, A2 => n95, ZN => B(16));
   U96 : OAI221_X1 port map( B1 => n44, B2 => n190, C1 => n164, C2 => n189, A 
                           => n152, ZN => n15);
   U97 : AOI22_X1 port map( A1 => A(13), A2 => n49, B1 => A(12), B2 => n50, ZN 
                           => n152);
   U98 : OAI221_X1 port map( B1 => n44, B2 => n195, C1 => n164, C2 => n194, A 
                           => n108, ZN => n11);
   U99 : AOI22_X1 port map( A1 => A(22), A2 => n49, B1 => A(21), B2 => n50, ZN 
                           => n108);
   U100 : OAI221_X1 port map( B1 => n44, B2 => n196, C1 => n166, C2 => n195, A 
                           => n139, ZN => n79);
   U101 : AOI22_X1 port map( A1 => A(23), A2 => n49, B1 => A(22), B2 => n50, ZN
                           => n139);
   U103 : OAI221_X1 port map( B1 => n44, B2 => n197, C1 => n165, C2 => n196, A 
                           => n131, ZN => n77);
   U104 : AOI22_X1 port map( A1 => A(24), A2 => n49, B1 => A(23), B2 => n50, ZN
                           => n131);
   U105 : AOI222_X1 port map( A1 => n71, A2 => n73, B1 => n67, B2 => n76, C1 =>
                           n11, C2 => n72, ZN => n31);
   U106 : AOI222_X1 port map( A1 => n78, A2 => n73, B1 => n59, B2 => n76, C1 =>
                           n79, C2 => n72, ZN => n25);
   U107 : AOI222_X1 port map( A1 => n75, A2 => n73, B1 => n58, B2 => n76, C1 =>
                           n77, C2 => n72, ZN => n19);
   U108 : AOI221_X1 port map( B1 => n51, B2 => A(7), C1 => n52, C2 => A(6), A 
                           => n161, ZN => n34);
   U109 : OAI22_X1 port map( A1 => n181, A2 => n55, B1 => n180, B2 => n57, ZN 
                           => n161);
   U110 : OAI221_X1 port map( B1 => n63, B2 => n3, C1 => n70, C2 => n177, A => 
                           n138, ZN => B(10));
   U111 : AOI222_X1 port map( A1 => n6, A2 => n28, B1 => n8, B2 => n29, C1 => 
                           n10, C2 => n79, ZN => n138);
   U112 : OAI221_X1 port map( B1 => n100, B2 => n38, C1 => n101, C2 => n3, A =>
                           n102, ZN => B(14));
   U113 : INV_X1 port map( A => n28, ZN => n101);
   U114 : INV_X1 port map( A => n29, ZN => n100);
   U115 : AOI222_X1 port map( A1 => n10, A2 => n78, B1 => n99, B2 => n59, C1 =>
                           n8, C2 => n79, ZN => n102);
   U116 : OAI221_X1 port map( B1 => n44, B2 => n191, C1 => n164, C2 => n190, A 
                           => n117, ZN => n7);
   U117 : AOI22_X1 port map( A1 => A(14), A2 => n49, B1 => A(13), B2 => n50, ZN
                           => n117);
   U118 : AOI22_X1 port map( A1 => n71, A2 => n72, B1 => n67, B2 => n73, ZN => 
                           n4);
   U119 : AOI22_X1 port map( A1 => n78, A2 => n72, B1 => n59, B2 => n73, ZN => 
                           n70);
   U120 : INV_X1 port map( A => SH(3), ZN => n170);
   U121 : NOR2_X1 port map( A1 => n173, A2 => n35, ZN => B(20));
   U122 : NOR2_X1 port map( A1 => n172, A2 => n13, ZN => B(24));
   U123 : INV_X1 port map( A => n22, ZN => n97);
   U124 : OAI221_X1 port map( B1 => n96, B2 => n38, C1 => n97, C2 => n3, A => 
                           n98, ZN => B(15));
   U125 : AOI222_X1 port map( A1 => n10, A2 => n75, B1 => n99, B2 => n58, C1 =>
                           n8, C2 => n77, ZN => n98);
   U126 : INV_X1 port map( A => n23, ZN => n96);
   U127 : AND2_X1 port map( A1 => n67, A2 => n41, ZN => B(29));
   U128 : AND2_X1 port map( A1 => n59, A2 => n41, ZN => B(30));
   U129 : BUF_X1 port map( A => SH(4), Z => n175);
   U130 : BUF_X1 port map( A => SH(4), Z => n176);
   U131 : INV_X1 port map( A => A(11), ZN => n187);
   U132 : INV_X1 port map( A => A(8), ZN => n184);
   U133 : INV_X1 port map( A => A(10), ZN => n186);
   U134 : INV_X1 port map( A => A(7), ZN => n183);
   U135 : INV_X1 port map( A => A(9), ZN => n185);
   U136 : OAI222_X1 port map( A1 => n55, A2 => n109, B1 => n164, B2 => n199, C1
                           => n57, C2 => n111, ZN => n67);
   U137 : OAI221_X1 port map( B1 => n44, B2 => n111, C1 => n164, C2 => n163, A 
                           => n142, ZN => n78);
   U138 : AOI22_X1 port map( A1 => A(27), A2 => n49, B1 => A(26), B2 => n50, ZN
                           => n142);
   U139 : OAI22_X1 port map( A1 => n57, A2 => n109, B1 => n55, B2 => n199, ZN 
                           => n59);
   U140 : AOI222_X1 port map( A1 => n74, A2 => n73, B1 => n68, B2 => n76, C1 =>
                           n17, C2 => n72, ZN => n35);
   U141 : AOI221_X1 port map( B1 => n17, B2 => n73, C1 => n16, C2 => n72, A => 
                           n154, ZN => n95);
   U142 : INV_X1 port map( A => n155, ZN => n154);
   U143 : AOI22_X1 port map( A1 => n92, A2 => n68, B1 => n76, B2 => n74, ZN => 
                           n155);
   U144 : AOI221_X1 port map( B1 => n11, B2 => n73, C1 => n9, C2 => n72, A => 
                           n93, ZN => n80);
   U145 : INV_X1 port map( A => n94, ZN => n93);
   U146 : AOI22_X1 port map( A1 => n92, A2 => n67, B1 => n76, B2 => n71, ZN => 
                           n94);
   U147 : OAI221_X1 port map( B1 => n12, B2 => n3, C1 => n13, C2 => n177, A => 
                           n14, ZN => B(8));
   U148 : AOI222_X1 port map( A1 => n6, A2 => n15, B1 => n8, B2 => n16, C1 => 
                           n10, C2 => n17, ZN => n14);
   U149 : OAI221_X1 port map( B1 => n34, B2 => n3, C1 => n35, C2 => n177, A => 
                           n36, ZN => B(4));
   U150 : AOI222_X1 port map( A1 => n6, A2 => n37, B1 => n8, B2 => n15, C1 => 
                           n10, C2 => n16, ZN => n36);
   U151 : OAI221_X1 port map( B1 => n30, B2 => n3, C1 => n31, C2 => n177, A => 
                           n32, ZN => B(5));
   U152 : AOI222_X1 port map( A1 => n6, A2 => n33, B1 => n8, B2 => n7, C1 => 
                           n10, C2 => n9, ZN => n32);
   U153 : OAI221_X1 port map( B1 => n44, B2 => n109, C1 => n165, C2 => n111, A 
                           => n127, ZN => n75);
   U154 : AOI22_X1 port map( A1 => A(28), A2 => n49, B1 => A(27), B2 => n50, ZN
                           => n127);
   U155 : OAI221_X1 port map( B1 => n119, B2 => n55, C1 => n135, C2 => n57, A 
                           => n140, ZN => n29);
   U156 : AOI22_X1 port map( A1 => A(21), A2 => n51, B1 => n52, B2 => A(20), ZN
                           => n140);
   U157 : OAI221_X1 port map( B1 => n192, B2 => n55, C1 => n119, C2 => n57, A 
                           => n128, ZN => n23);
   U158 : AOI22_X1 port map( A1 => A(22), A2 => n51, B1 => A(21), B2 => n52, ZN
                           => n128);
   U159 : INV_X1 port map( A => n121, ZN => B(12));
   U160 : AOI221_X1 port map( B1 => n16, B2 => n6, C1 => n15, C2 => n41, A => 
                           n122, ZN => n121);
   U161 : INV_X1 port map( A => n123, ZN => n122);
   U162 : AOI222_X1 port map( A1 => n10, A2 => n74, B1 => n99, B2 => n68, C1 =>
                           n8, C2 => n17, ZN => n123);
   U163 : OAI221_X1 port map( B1 => n2, B2 => n3, C1 => n4, C2 => n177, A => n5
                           , ZN => B(9));
   U164 : AOI222_X1 port map( A1 => n6, A2 => n7, B1 => n8, B2 => n9, C1 => n10
                           , C2 => n11, ZN => n5);
   U165 : OAI221_X1 port map( B1 => n103, B2 => n38, C1 => n104, C2 => n3, A =>
                           n105, ZN => B(13));
   U166 : INV_X1 port map( A => n7, ZN => n104);
   U167 : INV_X1 port map( A => n9, ZN => n103);
   U168 : AOI222_X1 port map( A1 => n10, A2 => n71, B1 => n99, B2 => n67, C1 =>
                           n8, C2 => n11, ZN => n105);
   U169 : OAI221_X1 port map( B1 => n44, B2 => n136, C1 => n166, C2 => n191, A 
                           => n141, ZN => n28);
   U170 : AOI22_X1 port map( A1 => A(15), A2 => n49, B1 => A(14), B2 => n50, ZN
                           => n141);
   U171 : OAI221_X1 port map( B1 => n44, B2 => n135, C1 => n166, C2 => n136, A 
                           => n137, ZN => n22);
   U172 : AOI22_X1 port map( A1 => A(16), A2 => n49, B1 => A(15), B2 => n50, ZN
                           => n137);
   U173 : AOI22_X1 port map( A1 => n74, A2 => n72, B1 => n68, B2 => n73, ZN => 
                           n13);
   U174 : AND2_X1 port map( A1 => n68, A2 => n41, ZN => B(28));
   U175 : OAI221_X1 port map( B1 => n44, B2 => n199, C1 => n165, C2 => n109, A 
                           => n157, ZN => n68);
   U176 : AOI22_X1 port map( A1 => A(29), A2 => n49, B1 => A(28), B2 => n50, ZN
                           => n157);
   U177 : OAI221_X1 port map( B1 => n44, B2 => n192, C1 => n165, C2 => n119, A 
                           => n120, ZN => n9);
   U178 : AOI22_X1 port map( A1 => A(18), A2 => n49, B1 => A(17), B2 => n50, ZN
                           => n120);
   U179 : OAI221_X1 port map( B1 => n44, B2 => n119, C1 => n165, C2 => n135, A 
                           => n158, ZN => n16);
   U180 : AOI22_X1 port map( A1 => A(17), A2 => n49, B1 => A(16), B2 => n50, ZN
                           => n158);
   U181 : INV_X1 port map( A => A(19), ZN => n119);
   U182 : INV_X1 port map( A => A(30), ZN => n109);
   U183 : INV_X1 port map( A => A(18), ZN => n135);
   U184 : INV_X1 port map( A => A(29), ZN => n111);
   U185 : INV_X1 port map( A => A(17), ZN => n136);
   U186 : INV_X1 port map( A => A(28), ZN => n163);
   U187 : INV_X1 port map( A => SH(0), ZN => n167);
   U188 : INV_X1 port map( A => SH(2), ZN => n168);
   U189 : INV_X1 port map( A => n170, ZN => n169);
   U190 : INV_X1 port map( A => A(2), ZN => n178);
   U191 : INV_X1 port map( A => A(3), ZN => n179);
   U192 : INV_X1 port map( A => A(4), ZN => n180);
   U193 : INV_X1 port map( A => A(5), ZN => n181);
   U194 : INV_X1 port map( A => A(6), ZN => n182);
   U195 : INV_X1 port map( A => A(12), ZN => n188);
   U196 : INV_X1 port map( A => A(14), ZN => n189);
   U197 : INV_X1 port map( A => A(15), ZN => n190);
   U198 : INV_X1 port map( A => A(16), ZN => n191);
   U199 : INV_X1 port map( A => A(20), ZN => n192);
   U200 : INV_X1 port map( A => A(21), ZN => n193);
   U201 : INV_X1 port map( A => A(23), ZN => n194);
   U202 : INV_X1 port map( A => A(24), ZN => n195);
   U203 : INV_X1 port map( A => A(25), ZN => n196);
   U204 : INV_X1 port map( A => A(26), ZN => n197);
   U205 : INV_X1 port map( A => A(27), ZN => n198);
   U206 : INV_X1 port map( A => A(31), ZN => n199);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Shifter_DATA_SIZE32_DW_sla_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end Shifter_DATA_SIZE32_DW_sla_0;

architecture SYN_mx2 of Shifter_DATA_SIZE32_DW_sla_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal B_31_port, B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, 
      B_25_port, B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, 
      B_19_port, B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, 
      B_13_port, B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port,
      B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, n2, n3, n4, 
      n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20
      , n21, n22, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, 
      n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50
      , n51, n52, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, 
      n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80
      , n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, 
      n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n120, 
      n121, n123, n126, n128, n129, n130, n131, n132, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n145, n147, n150, n151, n152, n155, n157, 
      n159, n160, n161, n162, n164, n166, n167, n168, n170, n171, n172, n174, 
      n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, 
      n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, 
      n199, n200, n201 : std_logic;

begin
   B <= ( B_31_port, B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, 
      B_25_port, B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, 
      B_19_port, B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, 
      B_13_port, B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port,
      B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, A(0) );
   
   U2 : NOR2_X2 port map( A1 => SH(2), A2 => SH(3), ZN => n75);
   U142 : MUX2_X1 port map( A => A(1), B => A(0), S => n34, Z => n79);
   U3 : NOR2_X1 port map( A1 => n177, A2 => SH(3), ZN => n73);
   U4 : INV_X1 port map( A => n34, ZN => n26);
   U5 : INV_X1 port map( A => n20, ZN => n37);
   U6 : INV_X1 port map( A => n22, ZN => n38);
   U7 : INV_X1 port map( A => n33, ZN => n25);
   U8 : NAND2_X1 port map( A1 => n175, A2 => n176, ZN => n34);
   U9 : OAI21_X1 port map( B1 => n183, B2 => n5, A => n3, ZN => B_7_port);
   U10 : OAI21_X1 port map( B1 => n183, B2 => n4, A => n3, ZN => B_8_port);
   U11 : OAI21_X1 port map( B1 => n181, B2 => n56, A => n3, ZN => B_11_port);
   U12 : OAI21_X1 port map( B1 => n181, B2 => n48, A => n3, ZN => B_12_port);
   U13 : OAI21_X1 port map( B1 => n182, B2 => n41, A => n3, ZN => B_13_port);
   U14 : OAI21_X1 port map( B1 => n181, B2 => n28, A => n3, ZN => B_14_port);
   U15 : OAI21_X1 port map( B1 => n181, B2 => n12, A => n3, ZN => B_15_port);
   U16 : NAND2_X1 port map( A1 => n184, A2 => A(0), ZN => n3);
   U17 : INV_X1 port map( A => n11, ZN => n58);
   U18 : INV_X1 port map( A => n184, ZN => n180);
   U19 : INV_X1 port map( A => n55, ZN => n16);
   U20 : OAI21_X1 port map( B1 => n182, B2 => n9, A => n3, ZN => B_3_port);
   U21 : OAI21_X1 port map( B1 => n182, B2 => n8, A => n3, ZN => B_4_port);
   U22 : OAI21_X1 port map( B1 => n183, B2 => n7, A => n3, ZN => B_5_port);
   U23 : OAI21_X1 port map( B1 => n183, B2 => n6, A => n3, ZN => B_6_port);
   U24 : OAI21_X1 port map( B1 => n183, B2 => n2, A => n3, ZN => B_9_port);
   U25 : OAI21_X1 port map( B1 => n181, B2 => n63, A => n3, ZN => B_10_port);
   U26 : NAND2_X1 port map( A1 => SH(0), A2 => n176, ZN => n33);
   U27 : NAND2_X1 port map( A1 => SH(0), A2 => SH(1), ZN => n22);
   U28 : AOI221_X1 port map( B1 => n94, B2 => n73, C1 => n95, C2 => n75, A => 
                           n88, ZN => n5);
   U29 : AOI221_X1 port map( B1 => n86, B2 => n73, C1 => n87, C2 => n75, A => 
                           n88, ZN => n4);
   U30 : AOI221_X1 port map( B1 => n74, B2 => n73, C1 => n70, C2 => n75, A => 
                           n141, ZN => n41);
   U31 : INV_X1 port map( A => n142, ZN => n141);
   U32 : AOI22_X1 port map( A1 => n136, A2 => n79, B1 => n78, B2 => n72, ZN => 
                           n142);
   U33 : AOI221_X1 port map( B1 => n92, B2 => n73, C1 => n59, C2 => n75, A => 
                           n134, ZN => n12);
   U34 : INV_X1 port map( A => n135, ZN => n134);
   U35 : AOI22_X1 port map( A1 => n136, A2 => n94, B1 => n78, B2 => n95, ZN => 
                           n135);
   U36 : NAND2_X1 port map( A1 => SH(1), A2 => n175, ZN => n20);
   U37 : OAI221_X1 port map( B1 => n128, B2 => n11, C1 => n112, C2 => n55, A =>
                           n129, ZN => B_16_port);
   U38 : INV_X1 port map( A => n84, ZN => n128);
   U39 : AOI221_X1 port map( B1 => n14, B2 => n86, C1 => n18, C2 => n87, A => 
                           n130, ZN => n129);
   U40 : INV_X1 port map( A => n3, ZN => n130);
   U41 : AOI221_X1 port map( B1 => n99, B2 => n73, C1 => n65, C2 => n75, A => 
                           n138, ZN => n28);
   U42 : INV_X1 port map( A => n139, ZN => n138);
   U43 : AOI22_X1 port map( A1 => n136, A2 => n101, B1 => n78, B2 => n102, ZN 
                           => n139);
   U44 : AOI221_X1 port map( B1 => n95, B2 => n73, C1 => n92, C2 => n75, A => 
                           n160, ZN => n56);
   U45 : INV_X1 port map( A => n161, ZN => n160);
   U46 : AOI21_X1 port map( B1 => n78, B2 => n94, A => n80, ZN => n161);
   U47 : AOI221_X1 port map( B1 => n87, B2 => n73, C1 => n84, C2 => n75, A => 
                           n151, ZN => n48);
   U48 : INV_X1 port map( A => n152, ZN => n151);
   U49 : AOI21_X1 port map( B1 => n78, B2 => n86, A => n80, ZN => n152);
   U50 : INV_X1 port map( A => n112, ZN => n50);
   U51 : INV_X1 port map( A => n60, ZN => n19);
   U52 : OAI222_X1 port map( A1 => n34, A2 => n187, B1 => n186, B2 => n33, C1 
                           => n185, C2 => n176, ZN => n101);
   U53 : NAND2_X1 port map( A1 => n75, A2 => n180, ZN => n55);
   U54 : AND2_X1 port map( A1 => n131, A2 => SH(2), ZN => n14);
   U55 : AOI221_X1 port map( B1 => n79, B2 => n73, C1 => n72, C2 => n75, A => 
                           n88, ZN => n7);
   U56 : AOI221_X1 port map( B1 => n101, B2 => n73, C1 => n102, C2 => n75, A =>
                           n88, ZN => n6);
   U57 : AOI221_X1 port map( B1 => n72, B2 => n73, C1 => n74, C2 => n75, A => 
                           n76, ZN => n2);
   U58 : INV_X1 port map( A => n77, ZN => n76);
   U59 : AOI21_X1 port map( B1 => n78, B2 => n79, A => n80, ZN => n77);
   U60 : AOI221_X1 port map( B1 => n102, B2 => n73, C1 => n99, C2 => n75, A => 
                           n167, ZN => n63);
   U61 : INV_X1 port map( A => n168, ZN => n167);
   U62 : AOI21_X1 port map( B1 => n78, B2 => n101, A => n80, ZN => n168);
   U63 : OAI21_X1 port map( B1 => n185, B2 => n177, A => n107, ZN => n113);
   U64 : NAND2_X1 port map( A1 => n73, A2 => n180, ZN => n11);
   U65 : NOR2_X1 port map( A1 => n177, A2 => n107, ZN => n80);
   U66 : AND2_X1 port map( A1 => n131, A2 => n177, ZN => n18);
   U67 : AOI21_X1 port map( B1 => n79, B2 => n75, A => n113, ZN => n116);
   U68 : AOI21_X1 port map( B1 => n101, B2 => n75, A => n113, ZN => n39);
   U69 : AOI21_X1 port map( B1 => n94, B2 => n75, A => n113, ZN => n9);
   U70 : AOI21_X1 port map( B1 => n86, B2 => n75, A => n113, ZN => n8);
   U71 : INV_X1 port map( A => n107, ZN => n88);
   U72 : BUF_X1 port map( A => n179, Z => n183);
   U73 : BUF_X1 port map( A => n178, Z => n182);
   U74 : BUF_X1 port map( A => n178, Z => n181);
   U75 : BUF_X1 port map( A => n179, Z => n184);
   U76 : OAI221_X1 port map( B1 => n33, B2 => n188, C1 => n34, C2 => n189, A =>
                           n145, ZN => n72);
   U77 : AOI22_X1 port map( A1 => A(3), A2 => n37, B1 => A(2), B2 => n38, ZN =>
                           n145);
   U78 : OAI221_X1 port map( B1 => n33, B2 => n190, C1 => n34, C2 => n191, A =>
                           n166, ZN => n95);
   U79 : AOI22_X1 port map( A1 => A(5), A2 => n37, B1 => A(4), B2 => n38, ZN =>
                           n166);
   U80 : OAI221_X1 port map( B1 => n33, B2 => n192, C1 => n34, C2 => n193, A =>
                           n150, ZN => n74);
   U81 : AOI22_X1 port map( A1 => A(7), A2 => n37, B1 => A(6), B2 => n38, ZN =>
                           n150);
   U82 : OAI221_X1 port map( B1 => n33, B2 => n193, C1 => n34, C2 => n194, A =>
                           n170, ZN => n99);
   U83 : AOI22_X1 port map( A1 => A(8), A2 => n37, B1 => A(7), B2 => n38, ZN =>
                           n170);
   U84 : OAI221_X1 port map( B1 => n33, B2 => n194, C1 => n34, C2 => n195, A =>
                           n164, ZN => n92);
   U85 : AOI22_X1 port map( A1 => A(9), A2 => n37, B1 => A(8), B2 => n38, ZN =>
                           n164);
   U86 : AOI221_X1 port map( B1 => n25, B2 => A(22), C1 => n26, C2 => A(23), A 
                           => n96, ZN => n60);
   U87 : INV_X1 port map( A => n97, ZN => n96);
   U88 : AOI22_X1 port map( A1 => A(21), A2 => n37, B1 => A(20), B2 => n38, ZN 
                           => n97);
   U89 : AOI221_X1 port map( B1 => n25, B2 => A(15), C1 => n26, C2 => A(16), A 
                           => n132, ZN => n112);
   U90 : OAI22_X1 port map( A1 => n198, A2 => n20, B1 => n197, B2 => n22, ZN =>
                           n132);
   U91 : INV_X1 port map( A => n171, ZN => n102);
   U92 : AOI221_X1 port map( B1 => n37, B2 => A(4), C1 => A(3), C2 => n38, A =>
                           n172, ZN => n171);
   U93 : OAI22_X1 port map( A1 => n189, A2 => n33, B1 => n190, B2 => n34, ZN =>
                           n172);
   U94 : OAI221_X1 port map( B1 => n60, B2 => n55, C1 => n5, C2 => n180, A => 
                           n91, ZN => B_23_port);
   U95 : AOI222_X1 port map( A1 => n58, A2 => n15, B1 => n18, B2 => n59, C1 => 
                           n14, C2 => n92, ZN => n91);
   U96 : OAI221_X1 port map( B1 => n47, B2 => n55, C1 => n4, C2 => n180, A => 
                           n83, ZN => B_24_port);
   U97 : AOI222_X1 port map( A1 => n58, A2 => n52, B1 => n18, B2 => n50, C1 => 
                           n14, C2 => n84, ZN => n83);
   U98 : OAI221_X1 port map( B1 => n40, B2 => n55, C1 => n2, C2 => n180, A => 
                           n69, ZN => B_25_port);
   U99 : AOI222_X1 port map( A1 => n58, A2 => n45, B1 => n18, B2 => n43, C1 => 
                           n14, C2 => n70, ZN => n69);
   U100 : OAI221_X1 port map( B1 => n27, B2 => n55, C1 => n63, C2 => n180, A =>
                           n64, ZN => B_26_port);
   U101 : AOI222_X1 port map( A1 => n58, A2 => n32, B1 => n18, B2 => n30, C1 =>
                           n14, C2 => n65, ZN => n64);
   U102 : OAI221_X1 port map( B1 => n10, B2 => n55, C1 => n56, C2 => n180, A =>
                           n57, ZN => B_27_port);
   U103 : AOI222_X1 port map( A1 => n58, A2 => n19, B1 => n18, B2 => n15, C1 =>
                           n14, C2 => n59, ZN => n57);
   U104 : OAI221_X1 port map( B1 => n47, B2 => n11, C1 => n48, C2 => n180, A =>
                           n49, ZN => B_28_port);
   U105 : AOI222_X1 port map( A1 => n14, A2 => n50, B1 => n16, B2 => n51, C1 =>
                           n18, C2 => n52, ZN => n49);
   U106 : OAI221_X1 port map( B1 => n33, B2 => n201, C1 => n34, C2 => n174, A 
                           => n54, ZN => n51);
   U107 : AOI22_X1 port map( A1 => A(26), A2 => n37, B1 => A(25), B2 => n38, ZN
                           => n54);
   U108 : OAI221_X1 port map( B1 => n33, B2 => n197, C1 => n34, C2 => n198, A 
                           => n140, ZN => n65);
   U109 : AOI22_X1 port map( A1 => A(12), A2 => n37, B1 => A(11), B2 => n38, ZN
                           => n140);
   U110 : OAI221_X1 port map( B1 => n33, B2 => n198, C1 => n34, C2 => n199, A 
                           => n137, ZN => n59);
   U111 : AOI22_X1 port map( A1 => A(13), A2 => n37, B1 => A(12), B2 => n38, ZN
                           => n137);
   U112 : OAI221_X1 port map( B1 => n33, B2 => n196, C1 => n34, C2 => n197, A 
                           => n147, ZN => n70);
   U113 : AOI22_X1 port map( A1 => A(11), A2 => n37, B1 => A(10), B2 => n38, ZN
                           => n147);
   U114 : OAI221_X1 port map( B1 => n33, B2 => n191, C1 => n34, C2 => n192, A 
                           => n159, ZN => n87);
   U115 : AOI22_X1 port map( A1 => A(6), A2 => n37, B1 => A(5), B2 => n38, ZN 
                           => n159);
   U116 : OAI221_X1 port map( B1 => n33, B2 => n195, C1 => n34, C2 => n196, A 
                           => n157, ZN => n84);
   U117 : AOI22_X1 port map( A1 => A(10), A2 => n37, B1 => A(9), B2 => n38, ZN 
                           => n157);
   U118 : OAI221_X1 port map( B1 => n20, B2 => n187, C1 => n186, C2 => n22, A 
                           => n155, ZN => n86);
   U119 : AOI22_X1 port map( A1 => n25, A2 => A(3), B1 => A(4), B2 => n26, ZN 
                           => n155);
   U120 : OAI221_X1 port map( B1 => n186, B2 => n20, C1 => n185, C2 => n22, A 
                           => n162, ZN => n94);
   U121 : AOI22_X1 port map( A1 => n25, A2 => A(2), B1 => A(3), B2 => n26, ZN 
                           => n162);
   U122 : OAI21_X1 port map( B1 => n182, B2 => n116, A => n3, ZN => B_1_port);
   U123 : OAI21_X1 port map( B1 => n182, B2 => n39, A => n3, ZN => B_2_port);
   U124 : AOI221_X1 port map( B1 => n25, B2 => A(23), C1 => n26, C2 => A(24), A
                           => n89, ZN => n47);
   U125 : INV_X1 port map( A => n90, ZN => n89);
   U126 : AOI22_X1 port map( A1 => A(22), A2 => n37, B1 => A(21), B2 => n38, ZN
                           => n90);
   U127 : AOI221_X1 port map( B1 => n25, B2 => A(24), C1 => n26, C2 => A(25), A
                           => n81, ZN => n40);
   U128 : INV_X1 port map( A => n82, ZN => n81);
   U129 : AOI22_X1 port map( A1 => A(23), A2 => n37, B1 => A(22), B2 => n38, ZN
                           => n82);
   U130 : AOI221_X1 port map( B1 => n25, B2 => A(25), C1 => n26, C2 => A(26), A
                           => n67, ZN => n27);
   U131 : INV_X1 port map( A => n68, ZN => n67);
   U132 : AOI22_X1 port map( A1 => A(24), A2 => n37, B1 => A(23), B2 => n38, ZN
                           => n68);
   U133 : AOI221_X1 port map( B1 => n25, B2 => A(26), C1 => n26, C2 => A(27), A
                           => n61, ZN => n10);
   U134 : INV_X1 port map( A => n62, ZN => n61);
   U135 : AOI22_X1 port map( A1 => A(25), A2 => n37, B1 => A(24), B2 => n38, ZN
                           => n62);
   U136 : AOI22_X1 port map( A1 => A(28), A2 => n37, B1 => A(27), B2 => n38, ZN
                           => n36);
   U137 : AND2_X1 port map( A1 => SH(3), A2 => n177, ZN => n78);
   U138 : NAND2_X1 port map( A1 => SH(3), A2 => A(0), ZN => n107);
   U139 : AND2_X1 port map( A1 => SH(2), A2 => SH(3), ZN => n136);
   U140 : AND2_X1 port map( A1 => SH(3), A2 => n180, ZN => n131);
   U141 : BUF_X1 port map( A => SH(4), Z => n179);
   U143 : BUF_X1 port map( A => SH(4), Z => n178);
   U144 : INV_X1 port map( A => A(2), ZN => n187);
   U145 : INV_X1 port map( A => A(16), ZN => n200);
   U146 : OAI221_X1 port map( B1 => n100, B2 => n55, C1 => n39, C2 => n180, A 
                           => n120, ZN => B_18_port);
   U147 : AOI222_X1 port map( A1 => n58, A2 => n65, B1 => n18, B2 => n99, C1 =>
                           n14, C2 => n102, ZN => n120);
   U148 : OAI221_X1 port map( B1 => n106, B2 => n55, C1 => n116, C2 => n180, A 
                           => n123, ZN => B_17_port);
   U149 : AOI222_X1 port map( A1 => n58, A2 => n70, B1 => n18, B2 => n74, C1 =>
                           n14, C2 => n72, ZN => n123);
   U150 : OAI221_X1 port map( B1 => n93, B2 => n55, C1 => n9, C2 => n180, A => 
                           n117, ZN => B_19_port);
   U151 : AOI222_X1 port map( A1 => n58, A2 => n59, B1 => n18, B2 => n92, C1 =>
                           n14, C2 => n95, ZN => n117);
   U152 : OAI221_X1 port map( B1 => n85, B2 => n55, C1 => n8, C2 => n180, A => 
                           n111, ZN => B_20_port);
   U153 : AOI222_X1 port map( A1 => n58, A2 => n50, B1 => n18, B2 => n84, C1 =>
                           n14, C2 => n87, ZN => n111);
   U154 : OAI221_X1 port map( B1 => n71, B2 => n55, C1 => n7, C2 => n180, A => 
                           n105, ZN => B_21_port);
   U155 : AOI222_X1 port map( A1 => n58, A2 => n43, B1 => n18, B2 => n70, C1 =>
                           n14, C2 => n74, ZN => n105);
   U156 : OAI221_X1 port map( B1 => n66, B2 => n55, C1 => n6, C2 => n180, A => 
                           n98, ZN => B_22_port);
   U157 : AOI222_X1 port map( A1 => n58, A2 => n30, B1 => n18, B2 => n65, C1 =>
                           n14, C2 => n99, ZN => n98);
   U158 : OAI221_X1 port map( B1 => n40, B2 => n11, C1 => n41, C2 => n180, A =>
                           n42, ZN => B_29_port);
   U159 : AOI222_X1 port map( A1 => n14, A2 => n43, B1 => n16, B2 => n44, C1 =>
                           n18, C2 => n45, ZN => n42);
   U160 : OAI221_X1 port map( B1 => n33, B2 => n174, C1 => n34, C2 => n21, A =>
                           n46, ZN => n44);
   U161 : AOI22_X1 port map( A1 => A(27), A2 => n37, B1 => A(26), B2 => n38, ZN
                           => n46);
   U162 : INV_X1 port map( A => n100, ZN => n30);
   U163 : INV_X1 port map( A => n93, ZN => n15);
   U164 : INV_X1 port map( A => n106, ZN => n43);
   U165 : INV_X1 port map( A => n85, ZN => n52);
   U166 : INV_X1 port map( A => n66, ZN => n32);
   U167 : INV_X1 port map( A => n71, ZN => n45);
   U168 : AOI221_X1 port map( B1 => n25, B2 => A(18), C1 => n26, C2 => A(19), A
                           => n118, ZN => n93);
   U169 : OAI22_X1 port map( A1 => n115, A2 => n20, B1 => n200, B2 => n22, ZN 
                           => n118);
   U170 : AOI221_X1 port map( B1 => n25, B2 => A(16), C1 => n26, C2 => A(17), A
                           => n126, ZN => n106);
   U171 : OAI22_X1 port map( A1 => n199, A2 => n20, B1 => n198, B2 => n22, ZN 
                           => n126);
   U172 : AOI221_X1 port map( B1 => n25, B2 => A(17), C1 => n26, C2 => A(18), A
                           => n121, ZN => n100);
   U173 : OAI22_X1 port map( A1 => n200, A2 => n20, B1 => n199, B2 => n22, ZN 
                           => n121);
   U174 : AOI221_X1 port map( B1 => n25, B2 => A(19), C1 => n26, C2 => A(20), A
                           => n114, ZN => n85);
   U175 : OAI22_X1 port map( A1 => n110, A2 => n20, B1 => n115, B2 => n22, ZN 
                           => n114);
   U176 : AOI221_X1 port map( B1 => n25, B2 => A(20), C1 => n26, C2 => A(21), A
                           => n108, ZN => n71);
   U177 : OAI22_X1 port map( A1 => n109, A2 => n20, B1 => n110, B2 => n22, ZN 
                           => n108);
   U178 : INV_X1 port map( A => A(19), ZN => n109);
   U179 : AOI221_X1 port map( B1 => n25, B2 => A(21), C1 => n26, C2 => A(22), A
                           => n103, ZN => n66);
   U180 : INV_X1 port map( A => n104, ZN => n103);
   U181 : AOI22_X1 port map( A1 => A(20), A2 => n37, B1 => A(19), B2 => n38, ZN
                           => n104);
   U182 : OAI221_X1 port map( B1 => n27, B2 => n11, C1 => n28, C2 => n180, A =>
                           n29, ZN => B_30_port);
   U183 : AOI222_X1 port map( A1 => n14, A2 => n30, B1 => n16, B2 => n31, C1 =>
                           n18, C2 => n32, ZN => n29);
   U184 : OAI221_X1 port map( B1 => n33, B2 => n21, C1 => n34, C2 => n35, A => 
                           n36, ZN => n31);
   U185 : INV_X1 port map( A => A(30), ZN => n35);
   U186 : OAI221_X1 port map( B1 => n10, B2 => n11, C1 => n12, C2 => n180, A =>
                           n13, ZN => B_31_port);
   U187 : AOI222_X1 port map( A1 => n14, A2 => n15, B1 => n16, B2 => n17, C1 =>
                           n18, C2 => n19, ZN => n13);
   U188 : OAI221_X1 port map( B1 => n20, B2 => n21, C1 => n22, C2 => n174, A =>
                           n24, ZN => n17);
   U189 : AOI22_X1 port map( A1 => A(30), A2 => n25, B1 => A(31), B2 => n26, ZN
                           => n24);
   U190 : INV_X1 port map( A => A(29), ZN => n21);
   U191 : INV_X1 port map( A => A(17), ZN => n115);
   U192 : INV_X1 port map( A => A(18), ZN => n110);
   U193 : INV_X1 port map( A => A(28), ZN => n174);
   U194 : INV_X1 port map( A => SH(0), ZN => n175);
   U195 : INV_X1 port map( A => SH(1), ZN => n176);
   U196 : INV_X1 port map( A => SH(2), ZN => n177);
   U197 : INV_X1 port map( A => A(0), ZN => n185);
   U198 : INV_X1 port map( A => A(1), ZN => n186);
   U199 : INV_X1 port map( A => A(4), ZN => n188);
   U200 : INV_X1 port map( A => A(5), ZN => n189);
   U201 : INV_X1 port map( A => A(6), ZN => n190);
   U202 : INV_X1 port map( A => A(7), ZN => n191);
   U203 : INV_X1 port map( A => A(8), ZN => n192);
   U204 : INV_X1 port map( A => A(9), ZN => n193);
   U205 : INV_X1 port map( A => A(10), ZN => n194);
   U206 : INV_X1 port map( A => A(11), ZN => n195);
   U207 : INV_X1 port map( A => A(12), ZN => n196);
   U208 : INV_X1 port map( A => A(13), ZN => n197);
   U209 : INV_X1 port map( A => A(14), ZN => n198);
   U210 : INV_X1 port map( A => A(15), ZN => n199);
   U211 : INV_X1 port map( A => A(27), ZN => n201);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Shifter_DATA_SIZE32_DW01_ash_0 is

   port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH : 
         in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out 
         std_logic_vector (31 downto 0));

end Shifter_DATA_SIZE32_DW01_ash_0;

architecture SYN_mx2 of Shifter_DATA_SIZE32_DW01_ash_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal ML_int_1_31_port, ML_int_1_30_port, ML_int_1_29_port, 
      ML_int_1_28_port, ML_int_1_27_port, ML_int_1_26_port, ML_int_1_25_port, 
      ML_int_1_24_port, ML_int_1_23_port, ML_int_1_22_port, ML_int_1_21_port, 
      ML_int_1_20_port, ML_int_1_19_port, ML_int_1_18_port, ML_int_1_17_port, 
      ML_int_1_16_port, ML_int_1_15_port, ML_int_1_14_port, ML_int_1_13_port, 
      ML_int_1_12_port, ML_int_1_11_port, ML_int_1_10_port, ML_int_1_9_port, 
      ML_int_1_8_port, ML_int_1_7_port, ML_int_1_6_port, ML_int_1_5_port, 
      ML_int_1_4_port, ML_int_1_3_port, ML_int_1_2_port, ML_int_1_1_port, 
      ML_int_1_0_port, ML_int_2_31_port, ML_int_2_30_port, ML_int_2_29_port, 
      ML_int_2_28_port, ML_int_2_27_port, ML_int_2_26_port, ML_int_2_25_port, 
      ML_int_2_24_port, ML_int_2_23_port, ML_int_2_22_port, ML_int_2_21_port, 
      ML_int_2_20_port, ML_int_2_19_port, ML_int_2_18_port, ML_int_2_17_port, 
      ML_int_2_16_port, ML_int_2_15_port, ML_int_2_14_port, ML_int_2_13_port, 
      ML_int_2_12_port, ML_int_2_11_port, ML_int_2_10_port, ML_int_2_9_port, 
      ML_int_2_8_port, ML_int_2_7_port, ML_int_2_6_port, ML_int_2_5_port, 
      ML_int_2_4_port, ML_int_2_3_port, ML_int_2_2_port, ML_int_2_1_port, 
      ML_int_2_0_port, ML_int_3_31_port, ML_int_3_30_port, ML_int_3_29_port, 
      ML_int_3_28_port, ML_int_3_27_port, ML_int_3_26_port, ML_int_3_25_port, 
      ML_int_3_24_port, ML_int_3_23_port, ML_int_3_22_port, ML_int_3_21_port, 
      ML_int_3_20_port, ML_int_3_19_port, ML_int_3_18_port, ML_int_3_17_port, 
      ML_int_3_16_port, ML_int_3_15_port, ML_int_3_14_port, ML_int_3_13_port, 
      ML_int_3_12_port, ML_int_3_11_port, ML_int_3_10_port, ML_int_3_9_port, 
      ML_int_3_8_port, ML_int_3_7_port, ML_int_3_6_port, ML_int_3_5_port, 
      ML_int_3_4_port, ML_int_3_3_port, ML_int_3_2_port, ML_int_3_1_port, 
      ML_int_3_0_port, ML_int_4_31_port, ML_int_4_30_port, ML_int_4_29_port, 
      ML_int_4_28_port, ML_int_4_27_port, ML_int_4_26_port, ML_int_4_25_port, 
      ML_int_4_24_port, ML_int_4_23_port, ML_int_4_22_port, ML_int_4_21_port, 
      ML_int_4_20_port, ML_int_4_19_port, ML_int_4_18_port, ML_int_4_17_port, 
      ML_int_4_16_port, ML_int_4_15_port, ML_int_4_14_port, ML_int_4_13_port, 
      ML_int_4_12_port, ML_int_4_11_port, ML_int_4_10_port, ML_int_4_9_port, 
      ML_int_4_8_port, ML_int_4_7_port, ML_int_4_6_port, ML_int_4_5_port, 
      ML_int_4_4_port, ML_int_4_3_port, ML_int_4_2_port, ML_int_4_1_port, 
      ML_int_4_0_port, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15
      , n16, n17, n18, n19, n20, n21 : std_logic;

begin
   
   M1_4_31 : MUX2_X1 port map( A => ML_int_4_31_port, B => ML_int_4_15_port, S 
                           => n20, Z => B(31));
   M1_4_30 : MUX2_X1 port map( A => ML_int_4_30_port, B => ML_int_4_14_port, S 
                           => n20, Z => B(30));
   M1_4_29 : MUX2_X1 port map( A => ML_int_4_29_port, B => ML_int_4_13_port, S 
                           => n20, Z => B(29));
   M1_4_28 : MUX2_X1 port map( A => ML_int_4_28_port, B => ML_int_4_12_port, S 
                           => n20, Z => B(28));
   M1_4_27 : MUX2_X1 port map( A => ML_int_4_27_port, B => ML_int_4_11_port, S 
                           => n20, Z => B(27));
   M1_4_26 : MUX2_X1 port map( A => ML_int_4_26_port, B => ML_int_4_10_port, S 
                           => SH(4), Z => B(26));
   M1_4_25 : MUX2_X1 port map( A => ML_int_4_25_port, B => ML_int_4_9_port, S 
                           => SH(4), Z => B(25));
   M1_4_24 : MUX2_X1 port map( A => ML_int_4_24_port, B => ML_int_4_8_port, S 
                           => SH(4), Z => B(24));
   M1_4_23 : MUX2_X1 port map( A => ML_int_4_23_port, B => ML_int_4_7_port, S 
                           => SH(4), Z => B(23));
   M1_4_22 : MUX2_X1 port map( A => ML_int_4_22_port, B => ML_int_4_6_port, S 
                           => SH(4), Z => B(22));
   M1_4_21 : MUX2_X1 port map( A => ML_int_4_21_port, B => ML_int_4_5_port, S 
                           => SH(4), Z => B(21));
   M1_4_20 : MUX2_X1 port map( A => ML_int_4_20_port, B => ML_int_4_4_port, S 
                           => SH(4), Z => B(20));
   M1_4_19 : MUX2_X1 port map( A => ML_int_4_19_port, B => ML_int_4_3_port, S 
                           => SH(4), Z => B(19));
   M1_4_18 : MUX2_X1 port map( A => ML_int_4_18_port, B => ML_int_4_2_port, S 
                           => SH(4), Z => B(18));
   M1_4_17 : MUX2_X1 port map( A => ML_int_4_17_port, B => ML_int_4_1_port, S 
                           => SH(4), Z => B(17));
   M1_4_16 : MUX2_X1 port map( A => ML_int_4_16_port, B => ML_int_4_0_port, S 
                           => n20, Z => B(16));
   M1_3_31 : MUX2_X1 port map( A => ML_int_3_31_port, B => ML_int_3_23_port, S 
                           => n18, Z => ML_int_4_31_port);
   M1_3_30 : MUX2_X1 port map( A => ML_int_3_30_port, B => ML_int_3_22_port, S 
                           => n18, Z => ML_int_4_30_port);
   M1_3_29 : MUX2_X1 port map( A => ML_int_3_29_port, B => ML_int_3_21_port, S 
                           => n18, Z => ML_int_4_29_port);
   M1_3_28 : MUX2_X1 port map( A => ML_int_3_28_port, B => ML_int_3_20_port, S 
                           => n18, Z => ML_int_4_28_port);
   M1_3_27 : MUX2_X1 port map( A => ML_int_3_27_port, B => ML_int_3_19_port, S 
                           => n18, Z => ML_int_4_27_port);
   M1_3_26 : MUX2_X1 port map( A => ML_int_3_26_port, B => ML_int_3_18_port, S 
                           => SH(3), Z => ML_int_4_26_port);
   M1_3_25 : MUX2_X1 port map( A => ML_int_3_25_port, B => ML_int_3_17_port, S 
                           => SH(3), Z => ML_int_4_25_port);
   M1_3_24 : MUX2_X1 port map( A => ML_int_3_24_port, B => ML_int_3_16_port, S 
                           => SH(3), Z => ML_int_4_24_port);
   M1_3_23 : MUX2_X1 port map( A => ML_int_3_23_port, B => ML_int_3_15_port, S 
                           => n18, Z => ML_int_4_23_port);
   M1_3_22 : MUX2_X1 port map( A => ML_int_3_22_port, B => ML_int_3_14_port, S 
                           => SH(3), Z => ML_int_4_22_port);
   M1_3_21 : MUX2_X1 port map( A => ML_int_3_21_port, B => ML_int_3_13_port, S 
                           => SH(3), Z => ML_int_4_21_port);
   M1_3_20 : MUX2_X1 port map( A => ML_int_3_20_port, B => ML_int_3_12_port, S 
                           => SH(3), Z => ML_int_4_20_port);
   M1_3_19 : MUX2_X1 port map( A => ML_int_3_19_port, B => ML_int_3_11_port, S 
                           => n18, Z => ML_int_4_19_port);
   M1_3_18 : MUX2_X1 port map( A => ML_int_3_18_port, B => ML_int_3_10_port, S 
                           => n18, Z => ML_int_4_18_port);
   M1_3_17 : MUX2_X1 port map( A => ML_int_3_17_port, B => ML_int_3_9_port, S 
                           => n18, Z => ML_int_4_17_port);
   M1_3_16 : MUX2_X1 port map( A => ML_int_3_16_port, B => ML_int_3_8_port, S 
                           => n18, Z => ML_int_4_16_port);
   M1_3_15 : MUX2_X1 port map( A => ML_int_3_15_port, B => ML_int_3_7_port, S 
                           => n18, Z => ML_int_4_15_port);
   M1_3_14 : MUX2_X1 port map( A => ML_int_3_14_port, B => ML_int_3_6_port, S 
                           => n18, Z => ML_int_4_14_port);
   M1_3_13 : MUX2_X1 port map( A => ML_int_3_13_port, B => ML_int_3_5_port, S 
                           => n18, Z => ML_int_4_13_port);
   M1_3_12 : MUX2_X1 port map( A => ML_int_3_12_port, B => ML_int_3_4_port, S 
                           => n18, Z => ML_int_4_12_port);
   M1_3_11 : MUX2_X1 port map( A => ML_int_3_11_port, B => ML_int_3_3_port, S 
                           => n18, Z => ML_int_4_11_port);
   M1_3_10 : MUX2_X1 port map( A => ML_int_3_10_port, B => ML_int_3_2_port, S 
                           => n18, Z => ML_int_4_10_port);
   M1_3_9 : MUX2_X1 port map( A => ML_int_3_9_port, B => ML_int_3_1_port, S => 
                           n18, Z => ML_int_4_9_port);
   M1_3_8 : MUX2_X1 port map( A => ML_int_3_8_port, B => ML_int_3_0_port, S => 
                           n18, Z => ML_int_4_8_port);
   M1_2_31 : MUX2_X1 port map( A => ML_int_2_31_port, B => ML_int_2_27_port, S 
                           => SH(2), Z => ML_int_3_31_port);
   M1_2_30 : MUX2_X1 port map( A => ML_int_2_30_port, B => ML_int_2_26_port, S 
                           => SH(2), Z => ML_int_3_30_port);
   M1_2_29 : MUX2_X1 port map( A => ML_int_2_29_port, B => ML_int_2_25_port, S 
                           => n16, Z => ML_int_3_29_port);
   M1_2_28 : MUX2_X1 port map( A => ML_int_2_28_port, B => ML_int_2_24_port, S 
                           => SH(2), Z => ML_int_3_28_port);
   M1_2_27 : MUX2_X1 port map( A => ML_int_2_27_port, B => ML_int_2_23_port, S 
                           => n16, Z => ML_int_3_27_port);
   M1_2_26 : MUX2_X1 port map( A => ML_int_2_26_port, B => ML_int_2_22_port, S 
                           => n16, Z => ML_int_3_26_port);
   M1_2_25 : MUX2_X1 port map( A => ML_int_2_25_port, B => ML_int_2_21_port, S 
                           => n16, Z => ML_int_3_25_port);
   M1_2_24 : MUX2_X1 port map( A => ML_int_2_24_port, B => ML_int_2_20_port, S 
                           => n16, Z => ML_int_3_24_port);
   M1_2_23 : MUX2_X1 port map( A => ML_int_2_23_port, B => ML_int_2_19_port, S 
                           => n16, Z => ML_int_3_23_port);
   M1_2_22 : MUX2_X1 port map( A => ML_int_2_22_port, B => ML_int_2_18_port, S 
                           => n16, Z => ML_int_3_22_port);
   M1_2_21 : MUX2_X1 port map( A => ML_int_2_21_port, B => ML_int_2_17_port, S 
                           => n16, Z => ML_int_3_21_port);
   M1_2_20 : MUX2_X1 port map( A => ML_int_2_20_port, B => ML_int_2_16_port, S 
                           => n16, Z => ML_int_3_20_port);
   M1_2_19 : MUX2_X1 port map( A => ML_int_2_19_port, B => ML_int_2_15_port, S 
                           => n16, Z => ML_int_3_19_port);
   M1_2_18 : MUX2_X1 port map( A => ML_int_2_18_port, B => ML_int_2_14_port, S 
                           => n16, Z => ML_int_3_18_port);
   M1_2_17 : MUX2_X1 port map( A => ML_int_2_17_port, B => ML_int_2_13_port, S 
                           => n16, Z => ML_int_3_17_port);
   M1_2_16 : MUX2_X1 port map( A => ML_int_2_16_port, B => ML_int_2_12_port, S 
                           => n16, Z => ML_int_3_16_port);
   M1_2_15 : MUX2_X1 port map( A => ML_int_2_15_port, B => ML_int_2_11_port, S 
                           => n16, Z => ML_int_3_15_port);
   M1_2_14 : MUX2_X1 port map( A => ML_int_2_14_port, B => ML_int_2_10_port, S 
                           => n16, Z => ML_int_3_14_port);
   M1_2_13 : MUX2_X1 port map( A => ML_int_2_13_port, B => ML_int_2_9_port, S 
                           => n16, Z => ML_int_3_13_port);
   M1_2_12 : MUX2_X1 port map( A => ML_int_2_12_port, B => ML_int_2_8_port, S 
                           => n16, Z => ML_int_3_12_port);
   M1_2_11 : MUX2_X1 port map( A => ML_int_2_11_port, B => ML_int_2_7_port, S 
                           => SH(2), Z => ML_int_3_11_port);
   M1_2_10 : MUX2_X1 port map( A => ML_int_2_10_port, B => ML_int_2_6_port, S 
                           => SH(2), Z => ML_int_3_10_port);
   M1_2_9 : MUX2_X1 port map( A => ML_int_2_9_port, B => ML_int_2_5_port, S => 
                           n16, Z => ML_int_3_9_port);
   M1_2_8 : MUX2_X1 port map( A => ML_int_2_8_port, B => ML_int_2_4_port, S => 
                           n16, Z => ML_int_3_8_port);
   M1_2_7 : MUX2_X1 port map( A => ML_int_2_7_port, B => ML_int_2_3_port, S => 
                           n16, Z => ML_int_3_7_port);
   M1_2_6 : MUX2_X1 port map( A => ML_int_2_6_port, B => ML_int_2_2_port, S => 
                           n16, Z => ML_int_3_6_port);
   M1_2_5 : MUX2_X1 port map( A => ML_int_2_5_port, B => ML_int_2_1_port, S => 
                           n16, Z => ML_int_3_5_port);
   M1_2_4 : MUX2_X1 port map( A => ML_int_2_4_port, B => ML_int_2_0_port, S => 
                           n16, Z => ML_int_3_4_port);
   M1_1_31 : MUX2_X1 port map( A => ML_int_1_31_port, B => ML_int_1_29_port, S 
                           => SH(1), Z => ML_int_2_31_port);
   M1_1_30 : MUX2_X1 port map( A => ML_int_1_30_port, B => ML_int_1_28_port, S 
                           => SH(1), Z => ML_int_2_30_port);
   M1_1_29 : MUX2_X1 port map( A => ML_int_1_29_port, B => ML_int_1_27_port, S 
                           => SH(1), Z => ML_int_2_29_port);
   M1_1_28 : MUX2_X1 port map( A => ML_int_1_28_port, B => ML_int_1_26_port, S 
                           => SH(1), Z => ML_int_2_28_port);
   M1_1_27 : MUX2_X1 port map( A => ML_int_1_27_port, B => ML_int_1_25_port, S 
                           => SH(1), Z => ML_int_2_27_port);
   M1_1_26 : MUX2_X1 port map( A => ML_int_1_26_port, B => ML_int_1_24_port, S 
                           => SH(1), Z => ML_int_2_26_port);
   M1_1_25 : MUX2_X1 port map( A => ML_int_1_25_port, B => ML_int_1_23_port, S 
                           => SH(1), Z => ML_int_2_25_port);
   M1_1_24 : MUX2_X1 port map( A => ML_int_1_24_port, B => ML_int_1_22_port, S 
                           => SH(1), Z => ML_int_2_24_port);
   M1_1_23 : MUX2_X1 port map( A => ML_int_1_23_port, B => ML_int_1_21_port, S 
                           => SH(1), Z => ML_int_2_23_port);
   M1_1_22 : MUX2_X1 port map( A => ML_int_1_22_port, B => ML_int_1_20_port, S 
                           => SH(1), Z => ML_int_2_22_port);
   M1_1_21 : MUX2_X1 port map( A => ML_int_1_21_port, B => ML_int_1_19_port, S 
                           => SH(1), Z => ML_int_2_21_port);
   M1_1_20 : MUX2_X1 port map( A => ML_int_1_20_port, B => ML_int_1_18_port, S 
                           => SH(1), Z => ML_int_2_20_port);
   M1_1_19 : MUX2_X1 port map( A => ML_int_1_19_port, B => ML_int_1_17_port, S 
                           => SH(1), Z => ML_int_2_19_port);
   M1_1_18 : MUX2_X1 port map( A => ML_int_1_18_port, B => ML_int_1_16_port, S 
                           => SH(1), Z => ML_int_2_18_port);
   M1_1_17 : MUX2_X1 port map( A => ML_int_1_17_port, B => ML_int_1_15_port, S 
                           => SH(1), Z => ML_int_2_17_port);
   M1_1_16 : MUX2_X1 port map( A => ML_int_1_16_port, B => ML_int_1_14_port, S 
                           => SH(1), Z => ML_int_2_16_port);
   M1_1_15 : MUX2_X1 port map( A => ML_int_1_15_port, B => ML_int_1_13_port, S 
                           => SH(1), Z => ML_int_2_15_port);
   M1_1_14 : MUX2_X1 port map( A => ML_int_1_14_port, B => ML_int_1_12_port, S 
                           => SH(1), Z => ML_int_2_14_port);
   M1_1_13 : MUX2_X1 port map( A => ML_int_1_13_port, B => ML_int_1_11_port, S 
                           => n14, Z => ML_int_2_13_port);
   M1_1_12 : MUX2_X1 port map( A => ML_int_1_12_port, B => ML_int_1_10_port, S 
                           => n14, Z => ML_int_2_12_port);
   M1_1_11 : MUX2_X1 port map( A => ML_int_1_11_port, B => ML_int_1_9_port, S 
                           => n14, Z => ML_int_2_11_port);
   M1_1_10 : MUX2_X1 port map( A => ML_int_1_10_port, B => ML_int_1_8_port, S 
                           => n14, Z => ML_int_2_10_port);
   M1_1_9 : MUX2_X1 port map( A => ML_int_1_9_port, B => ML_int_1_7_port, S => 
                           n14, Z => ML_int_2_9_port);
   M1_1_8 : MUX2_X1 port map( A => ML_int_1_8_port, B => ML_int_1_6_port, S => 
                           n14, Z => ML_int_2_8_port);
   M1_1_7 : MUX2_X1 port map( A => ML_int_1_7_port, B => ML_int_1_5_port, S => 
                           n14, Z => ML_int_2_7_port);
   M1_1_6 : MUX2_X1 port map( A => ML_int_1_6_port, B => ML_int_1_4_port, S => 
                           n14, Z => ML_int_2_6_port);
   M1_1_5 : MUX2_X1 port map( A => ML_int_1_5_port, B => ML_int_1_3_port, S => 
                           n14, Z => ML_int_2_5_port);
   M1_1_4 : MUX2_X1 port map( A => ML_int_1_4_port, B => ML_int_1_2_port, S => 
                           n14, Z => ML_int_2_4_port);
   M1_1_3 : MUX2_X1 port map( A => ML_int_1_3_port, B => ML_int_1_1_port, S => 
                           n14, Z => ML_int_2_3_port);
   M1_1_2 : MUX2_X1 port map( A => ML_int_1_2_port, B => ML_int_1_0_port, S => 
                           n14, Z => ML_int_2_2_port);
   M1_0_31 : MUX2_X1 port map( A => A(31), B => A(30), S => SH(0), Z => 
                           ML_int_1_31_port);
   M1_0_30 : MUX2_X1 port map( A => A(30), B => A(29), S => SH(0), Z => 
                           ML_int_1_30_port);
   M1_0_29 : MUX2_X1 port map( A => A(29), B => A(28), S => SH(0), Z => 
                           ML_int_1_29_port);
   M1_0_28 : MUX2_X1 port map( A => A(28), B => A(27), S => SH(0), Z => 
                           ML_int_1_28_port);
   M1_0_27 : MUX2_X1 port map( A => A(27), B => A(26), S => SH(0), Z => 
                           ML_int_1_27_port);
   M1_0_26 : MUX2_X1 port map( A => A(26), B => A(25), S => SH(0), Z => 
                           ML_int_1_26_port);
   M1_0_25 : MUX2_X1 port map( A => A(25), B => A(24), S => n12, Z => 
                           ML_int_1_25_port);
   M1_0_24 : MUX2_X1 port map( A => A(24), B => A(23), S => n12, Z => 
                           ML_int_1_24_port);
   M1_0_23 : MUX2_X1 port map( A => A(23), B => A(22), S => n12, Z => 
                           ML_int_1_23_port);
   M1_0_22 : MUX2_X1 port map( A => A(22), B => A(21), S => n12, Z => 
                           ML_int_1_22_port);
   M1_0_21 : MUX2_X1 port map( A => A(21), B => A(20), S => n12, Z => 
                           ML_int_1_21_port);
   M1_0_20 : MUX2_X1 port map( A => A(20), B => A(19), S => n12, Z => 
                           ML_int_1_20_port);
   M1_0_19 : MUX2_X1 port map( A => A(19), B => A(18), S => n12, Z => 
                           ML_int_1_19_port);
   M1_0_18 : MUX2_X1 port map( A => A(18), B => A(17), S => n12, Z => 
                           ML_int_1_18_port);
   M1_0_17 : MUX2_X1 port map( A => A(17), B => A(16), S => n12, Z => 
                           ML_int_1_17_port);
   M1_0_16 : MUX2_X1 port map( A => A(16), B => A(15), S => n12, Z => 
                           ML_int_1_16_port);
   M1_0_15 : MUX2_X1 port map( A => A(15), B => A(14), S => n12, Z => 
                           ML_int_1_15_port);
   M1_0_14 : MUX2_X1 port map( A => A(14), B => A(13), S => n12, Z => 
                           ML_int_1_14_port);
   M1_0_13 : MUX2_X1 port map( A => A(13), B => A(12), S => n12, Z => 
                           ML_int_1_13_port);
   M1_0_12 : MUX2_X1 port map( A => A(12), B => A(11), S => n11, Z => 
                           ML_int_1_12_port);
   M1_0_11 : MUX2_X1 port map( A => A(11), B => A(10), S => n11, Z => 
                           ML_int_1_11_port);
   M1_0_10 : MUX2_X1 port map( A => A(10), B => A(9), S => n11, Z => 
                           ML_int_1_10_port);
   M1_0_9 : MUX2_X1 port map( A => A(9), B => A(8), S => n11, Z => 
                           ML_int_1_9_port);
   M1_0_8 : MUX2_X1 port map( A => A(8), B => A(7), S => n11, Z => 
                           ML_int_1_8_port);
   M1_0_7 : MUX2_X1 port map( A => A(7), B => A(6), S => n11, Z => 
                           ML_int_1_7_port);
   M1_0_6 : MUX2_X1 port map( A => A(6), B => A(5), S => n11, Z => 
                           ML_int_1_6_port);
   M1_0_5 : MUX2_X1 port map( A => A(5), B => A(4), S => n11, Z => 
                           ML_int_1_5_port);
   M1_0_4 : MUX2_X1 port map( A => A(4), B => A(3), S => n11, Z => 
                           ML_int_1_4_port);
   M1_0_3 : MUX2_X1 port map( A => A(3), B => A(2), S => n11, Z => 
                           ML_int_1_3_port);
   M1_0_2 : MUX2_X1 port map( A => A(2), B => A(1), S => n11, Z => 
                           ML_int_1_2_port);
   M1_0_1 : MUX2_X1 port map( A => A(1), B => A(0), S => n11, Z => 
                           ML_int_1_1_port);
   U3 : INV_X1 port map( A => n13, ZN => n11);
   U4 : INV_X1 port map( A => n13, ZN => n12);
   U5 : INV_X1 port map( A => n15, ZN => n14);
   U6 : INV_X1 port map( A => n17, ZN => n16);
   U7 : NOR2_X1 port map( A1 => n20, A2 => n9, ZN => B(1));
   U8 : NOR2_X1 port map( A1 => n20, A2 => n8, ZN => B(2));
   U9 : NOR2_X1 port map( A1 => n20, A2 => n7, ZN => B(3));
   U10 : NOR2_X1 port map( A1 => n20, A2 => n5, ZN => B(5));
   U11 : NOR2_X1 port map( A1 => n20, A2 => n3, ZN => B(7));
   U12 : INV_X1 port map( A => n10, ZN => ML_int_4_0_port);
   U13 : AND2_X1 port map( A1 => ML_int_2_2_port, A2 => n17, ZN => 
                           ML_int_3_2_port);
   U14 : AND2_X1 port map( A1 => ML_int_2_3_port, A2 => n17, ZN => 
                           ML_int_3_3_port);
   U15 : AND2_X1 port map( A1 => ML_int_2_0_port, A2 => n17, ZN => 
                           ML_int_3_0_port);
   U16 : AND2_X1 port map( A1 => ML_int_2_1_port, A2 => n17, ZN => 
                           ML_int_3_1_port);
   U17 : INV_X1 port map( A => n21, ZN => n20);
   U18 : INV_X1 port map( A => n19, ZN => n18);
   U19 : INV_X1 port map( A => SH(0), ZN => n13);
   U20 : INV_X1 port map( A => SH(1), ZN => n15);
   U21 : INV_X1 port map( A => SH(2), ZN => n17);
   U22 : NAND2_X1 port map( A1 => ML_int_3_0_port, A2 => n19, ZN => n10);
   U23 : NAND2_X1 port map( A1 => ML_int_3_1_port, A2 => n19, ZN => n9);
   U24 : NAND2_X1 port map( A1 => ML_int_3_2_port, A2 => n19, ZN => n8);
   U25 : NAND2_X1 port map( A1 => ML_int_3_3_port, A2 => n19, ZN => n7);
   U26 : NAND2_X1 port map( A1 => ML_int_3_4_port, A2 => n19, ZN => n6);
   U27 : NAND2_X1 port map( A1 => ML_int_3_5_port, A2 => n19, ZN => n5);
   U28 : NAND2_X1 port map( A1 => ML_int_3_6_port, A2 => n19, ZN => n4);
   U29 : NAND2_X1 port map( A1 => ML_int_3_7_port, A2 => n19, ZN => n3);
   U30 : INV_X1 port map( A => n9, ZN => ML_int_4_1_port);
   U31 : INV_X1 port map( A => n8, ZN => ML_int_4_2_port);
   U32 : INV_X1 port map( A => n7, ZN => ML_int_4_3_port);
   U33 : INV_X1 port map( A => n6, ZN => ML_int_4_4_port);
   U34 : INV_X1 port map( A => n5, ZN => ML_int_4_5_port);
   U35 : INV_X1 port map( A => n4, ZN => ML_int_4_6_port);
   U36 : INV_X1 port map( A => n3, ZN => ML_int_4_7_port);
   U37 : AND2_X1 port map( A1 => ML_int_1_0_port, A2 => n15, ZN => 
                           ML_int_2_0_port);
   U38 : AND2_X1 port map( A1 => ML_int_1_1_port, A2 => n15, ZN => 
                           ML_int_2_1_port);
   U39 : AND2_X1 port map( A1 => ML_int_4_11_port, A2 => n21, ZN => B(11));
   U40 : AND2_X1 port map( A1 => ML_int_4_12_port, A2 => n21, ZN => B(12));
   U41 : AND2_X1 port map( A1 => ML_int_4_13_port, A2 => n21, ZN => B(13));
   U42 : AND2_X1 port map( A1 => ML_int_4_14_port, A2 => n21, ZN => B(14));
   U43 : AND2_X1 port map( A1 => ML_int_4_15_port, A2 => n21, ZN => B(15));
   U44 : NOR2_X1 port map( A1 => n20, A2 => n6, ZN => B(4));
   U45 : NOR2_X1 port map( A1 => n20, A2 => n4, ZN => B(6));
   U46 : AND2_X1 port map( A1 => ML_int_4_8_port, A2 => n21, ZN => B(8));
   U47 : AND2_X1 port map( A1 => ML_int_4_9_port, A2 => n21, ZN => B(9));
   U48 : NOR2_X1 port map( A1 => n20, A2 => n10, ZN => B(0));
   U49 : AND2_X1 port map( A1 => ML_int_4_10_port, A2 => n21, ZN => B(10));
   U50 : INV_X1 port map( A => SH(4), ZN => n21);
   U51 : AND2_X1 port map( A1 => A(0), A2 => n13, ZN => ML_int_1_0_port);
   U52 : INV_X1 port map( A => SH(3), ZN => n19);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderSumGenerator_DATA_SIZE32_SPARSITY4_0 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic_vector 
         (7 downto 0);  sum : out std_logic_vector (31 downto 0));

end AdderSumGenerator_DATA_SIZE32_SPARSITY4_0;

architecture SYN_adder_sum_generator_arch of 
   AdderSumGenerator_DATA_SIZE32_SPARSITY4_0 is

   component AdderCarrySelect_DATA_SIZE4_77
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_78
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_79
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_80
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_81
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_82
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_83
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_0
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;

begin
   
   ACSi_0 : AdderCarrySelect_DATA_SIZE4_0 port map( a(3) => a(3), a(2) => a(2),
                           a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), sel => cin(0), 
                           sum(3) => sum(3), sum(2) => sum(2), sum(1) => sum(1)
                           , sum(0) => sum(0));
   ACSi_1 : AdderCarrySelect_DATA_SIZE4_83 port map( a(3) => a(7), a(2) => a(6)
                           , a(1) => a(5), a(0) => a(4), b(3) => b(7), b(2) => 
                           b(6), b(1) => b(5), b(0) => b(4), sel => cin(1), 
                           sum(3) => sum(7), sum(2) => sum(6), sum(1) => sum(5)
                           , sum(0) => sum(4));
   ACSi_2 : AdderCarrySelect_DATA_SIZE4_82 port map( a(3) => a(11), a(2) => 
                           a(10), a(1) => a(9), a(0) => a(8), b(3) => b(11), 
                           b(2) => b(10), b(1) => b(9), b(0) => b(8), sel => 
                           cin(2), sum(3) => sum(11), sum(2) => sum(10), sum(1)
                           => sum(9), sum(0) => sum(8));
   ACSi_3 : AdderCarrySelect_DATA_SIZE4_81 port map( a(3) => a(15), a(2) => 
                           a(14), a(1) => a(13), a(0) => a(12), b(3) => b(15), 
                           b(2) => b(14), b(1) => b(13), b(0) => b(12), sel => 
                           cin(3), sum(3) => sum(15), sum(2) => sum(14), sum(1)
                           => sum(13), sum(0) => sum(12));
   ACSi_4 : AdderCarrySelect_DATA_SIZE4_80 port map( a(3) => a(19), a(2) => 
                           a(18), a(1) => a(17), a(0) => a(16), b(3) => b(19), 
                           b(2) => b(18), b(1) => b(17), b(0) => b(16), sel => 
                           cin(4), sum(3) => sum(19), sum(2) => sum(18), sum(1)
                           => sum(17), sum(0) => sum(16));
   ACSi_5 : AdderCarrySelect_DATA_SIZE4_79 port map( a(3) => a(23), a(2) => 
                           a(22), a(1) => a(21), a(0) => a(20), b(3) => b(23), 
                           b(2) => b(22), b(1) => b(21), b(0) => b(20), sel => 
                           cin(5), sum(3) => sum(23), sum(2) => sum(22), sum(1)
                           => sum(21), sum(0) => sum(20));
   ACSi_6 : AdderCarrySelect_DATA_SIZE4_78 port map( a(3) => a(27), a(2) => 
                           a(26), a(1) => a(25), a(0) => a(24), b(3) => b(27), 
                           b(2) => b(26), b(1) => b(25), b(0) => b(24), sel => 
                           cin(6), sum(3) => sum(27), sum(2) => sum(26), sum(1)
                           => sum(25), sum(0) => sum(24));
   ACSi_7 : AdderCarrySelect_DATA_SIZE4_77 port map( a(3) => a(31), a(2) => 
                           a(30), a(1) => a(29), a(0) => a(28), b(3) => b(31), 
                           b(2) => b(30), b(1) => b(29), b(0) => b(28), sel => 
                           cin(7), sum(3) => sum(31), sum(2) => sum(30), sum(1)
                           => sum(29), sum(0) => sum(28));

end SYN_adder_sum_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4CarryGenerator_DATA_SIZE32_SPARSITY4_0 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  cout :
         out std_logic_vector (7 downto 0));

end P4CarryGenerator_DATA_SIZE32_SPARSITY4_0;

architecture SYN_p4_carry_generator_arch of 
   P4CarryGenerator_DATA_SIZE32_SPARSITY4_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n267, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n69, n73, n74
      , n75, n76, n77, n78, n79, n82, n102, n103, net138479, net138523, 
      net138522, net138519, net138537, net138629, net138840, net149048, 
      net150785, net150986, net150985, net150984, net150981, net150978, 
      net150977, net150964, net150962, net150961, net150953, net150952, 
      net150951, net150938, net150936, net150935, net150934, net150929, 
      net150923, net150922, net150920, net150919, net150916, net150902, 
      net150897, net150882, net151486, net151669, net151668, net151667, 
      net151653, net151647, net151646, net151645, net151639, net151615, 
      net152639, net152653, net152678, net152799, net152783, net152766, 
      net152763, net152760, net152759, net152747, net152743, net152737, 
      net152735, net153401, net153399, net153520, net153540, net153539, 
      net153553, net153787, net153762, net153760, net154049, net154277, 
      net154289, net153400, net138535, n104, n105, n106, n107, n108, n109, n110
      , n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n264, n265 : std_logic;

begin
   
   cout_5_inst : NAND3_X1 port map( A1 => n233, A2 => net150882, A3 => n234, ZN
                           => cout(5));
   net151579 : NAND3_X1 port map( A1 => a(16), A2 => b(16), A3 => n79, ZN => 
                           n78);
   net152714 : NAND3_X1 port map( A1 => net152735, A2 => n187, A3 => net152737,
                           ZN => net138537);
   syn97 : NAND3_X1 port map( A1 => n180, A2 => n181, A3 => n104, ZN => n179);
   syn172 : NAND3_X1 port map( A1 => n164, A2 => net153400, A3 => n105, ZN => 
                           n157);
   U1 : INV_X1 port map( A => a(12), ZN => n171);
   U2 : NAND2_X1 port map( A1 => net150923, A2 => n242, ZN => net150922);
   U3 : NAND2_X1 port map( A1 => n110, A2 => n111, ZN => net150923);
   U4 : NAND2_X1 port map( A1 => n238, A2 => n239, ZN => n242);
   U5 : INV_X1 port map( A => b(27), ZN => n238);
   U6 : INV_X1 port map( A => n112, ZN => n115);
   U7 : OAI211_X1 port map( C1 => n110, C2 => n111, A => n113, B => net150916, 
                           ZN => n112);
   U8 : NAND2_X1 port map( A1 => b(25), A2 => a(25), ZN => n113);
   U9 : INV_X1 port map( A => a(4), ZN => n205);
   U10 : INV_X1 port map( A => a(18), ZN => n227);
   U11 : INV_X1 port map( A => a(22), ZN => n253);
   U12 : NAND2_X1 port map( A1 => a(21), A2 => b(21), ZN => net150964);
   U13 : NAND2_X1 port map( A1 => n218, A2 => n219, ZN => n212);
   U14 : INV_X1 port map( A => b(21), ZN => n218);
   U15 : INV_X1 port map( A => a(21), ZN => n219);
   U16 : INV_X1 port map( A => n140, ZN => net151667);
   U17 : NAND2_X1 port map( A1 => net151653, A2 => n224, ZN => n225);
   U18 : NAND2_X1 port map( A1 => net150964, A2 => n253, ZN => net150935);
   U19 : NAND2_X1 port map( A1 => net150964, A2 => n254, ZN => net150934);
   U20 : NOR2_X1 port map( A1 => net150922, A2 => n122, ZN => n123);
   U21 : NAND2_X1 port map( A1 => n115, A2 => net150919, ZN => n114);
   U22 : INV_X1 port map( A => b(24), ZN => net150919);
   U23 : NOR2_X1 port map( A1 => a(5), A2 => b(5), ZN => net152747);
   U24 : INV_X1 port map( A => a(5), ZN => n206);
   U25 : INV_X1 port map( A => a(9), ZN => n153);
   U26 : NAND2_X1 port map( A1 => a(8), A2 => b(8), ZN => n156);
   U27 : INV_X1 port map( A => a(8), ZN => n154);
   U28 : AND3_X1 port map( A1 => n166, A2 => n171, A3 => n104, ZN => n182);
   U29 : NAND2_X1 port map( A1 => n254, A2 => n253, ZN => net150929);
   U30 : INV_X1 port map( A => n114, ZN => net150938);
   U31 : NAND2_X1 port map( A1 => n124, A2 => n129, ZN => n118);
   U32 : AOI21_X1 port map( B1 => n124, B2 => a(24), A => n125, ZN => n119);
   U33 : INV_X1 port map( A => net150882, ZN => n129);
   U34 : NAND2_X1 port map( A1 => net150936, A2 => n115, ZN => net150951);
   U35 : NOR2_X1 port map( A1 => b(25), A2 => a(25), ZN => net150936);
   U36 : AND2_X1 port map( A1 => n176, A2 => net153762, ZN => net153760);
   U37 : NAND2_X1 port map( A1 => a(9), A2 => b(9), ZN => net153762);
   U38 : NAND2_X1 port map( A1 => b(10), A2 => a(10), ZN => n176);
   U39 : NAND2_X1 port map( A1 => b(19), A2 => a(19), ZN => n220);
   U40 : NAND2_X1 port map( A1 => n216, A2 => n217, ZN => n230);
   U41 : NAND2_X1 port map( A1 => n215, A2 => n214, ZN => n231);
   U42 : NAND2_X1 port map( A1 => n227, A2 => n226, ZN => n229);
   U43 : NAND2_X1 port map( A1 => a(23), A2 => net150929, ZN => n243);
   U44 : NAND2_X1 port map( A1 => b(23), A2 => net150929, ZN => n240);
   U45 : INV_X1 port map( A => a(7), ZN => n102);
   U46 : INV_X1 port map( A => a(6), ZN => n148);
   U47 : OAI22_X1 port map( A1 => a(7), A2 => b(7), B1 => a(6), B2 => b(6), ZN 
                           => n146);
   U48 : INV_X1 port map( A => net151639, ZN => n141);
   U49 : NAND2_X1 port map( A1 => net151669, A2 => n141, ZN => n136);
   U50 : INV_X1 port map( A => n243, ZN => n255);
   U51 : NAND2_X1 port map( A1 => a(23), A2 => b(23), ZN => net150882);
   U52 : NAND2_X1 port map( A1 => net150934, A2 => net150935, ZN => net150984);
   U53 : NAND2_X1 port map( A1 => net150934, A2 => net150935, ZN => net150985);
   U54 : INV_X1 port map( A => n240, ZN => n256);
   U55 : NAND2_X1 port map( A1 => net151653, A2 => n224, ZN => n223);
   U56 : INV_X1 port map( A => cin, ZN => n108);
   U57 : INV_X1 port map( A => a(27), ZN => n239);
   U58 : INV_X1 port map( A => a(26), ZN => n111);
   U59 : INV_X1 port map( A => b(26), ZN => n110);
   U60 : NAND2_X1 port map( A1 => a(27), A2 => b(27), ZN => net150916);
   U61 : NAND2_X1 port map( A1 => b(23), A2 => net150929, ZN => n122);
   U62 : NAND2_X1 port map( A1 => net150934, A2 => net150935, ZN => n132);
   U63 : NOR2_X1 port map( A1 => net150922, A2 => n120, ZN => n121);
   U64 : NAND2_X1 port map( A1 => a(23), A2 => net150929, ZN => n120);
   U65 : NAND2_X1 port map( A1 => net150934, A2 => net150935, ZN => n133);
   U66 : NAND2_X1 port map( A1 => net150934, A2 => net150935, ZN => net150986);
   U67 : NAND2_X1 port map( A1 => net150934, A2 => net150935, ZN => n258);
   U68 : NOR2_X1 port map( A1 => a(4), A2 => b(4), ZN => n191);
   U69 : INV_X1 port map( A => b(4), ZN => n201);
   U70 : INV_X1 port map( A => net150929, ZN => net150952);
   U71 : AOI21_X1 port map( B1 => net150934, B2 => net150935, A => net150897, 
                           ZN => n246);
   U72 : INV_X1 port map( A => net150916, ZN => n125);
   U73 : INV_X1 port map( A => net150922, ZN => n124);
   U74 : INV_X1 port map( A => b(2), ZN => n195);
   U75 : INV_X1 port map( A => b(5), ZN => n147);
   U76 : INV_X1 port map( A => b(9), ZN => n152);
   U77 : INV_X1 port map( A => a(13), ZN => net138522);
   U78 : INV_X1 port map( A => b(13), ZN => net138523);
   U79 : INV_X1 port map( A => b(12), ZN => n180);
   U80 : NAND2_X1 port map( A1 => n175, A2 => n177, ZN => n173);
   U81 : NOR2_X1 port map( A1 => n178, A2 => n171, ZN => n177);
   U82 : INV_X1 port map( A => n174, ZN => n178);
   U83 : INV_X1 port map( A => b(18), ZN => n226);
   U84 : INV_X1 port map( A => a(16), ZN => n215);
   U85 : INV_X1 port map( A => b(16), ZN => n214);
   U86 : INV_X1 port map( A => a(19), ZN => n216);
   U87 : INV_X1 port map( A => b(19), ZN => n217);
   U88 : NAND2_X1 port map( A1 => n141, A2 => n138, ZN => n140);
   U89 : INV_X1 port map( A => a(20), ZN => n138);
   U90 : NAND2_X1 port map( A1 => n139, A2 => a(20), ZN => net151645);
   U91 : NAND2_X1 port map( A1 => net151669, A2 => n141, ZN => n139);
   U92 : NAND2_X1 port map( A1 => net151639, A2 => a(20), ZN => net151653);
   U93 : INV_X1 port map( A => b(20), ZN => n224);
   U94 : INV_X1 port map( A => b(22), ZN => n254);
   U95 : NOR2_X1 port map( A1 => net150952, A2 => net150922, ZN => n244);
   U96 : NAND2_X1 port map( A1 => net150934, A2 => net150935, ZN => n259);
   U97 : NOR2_X1 port map( A1 => n236, A2 => n237, ZN => n235);
   U98 : NOR2_X1 port map( A1 => n240, A2 => n241, ZN => n236);
   U99 : OAI21_X1 port map( B1 => n243, B2 => n246, A => net150882, ZN => n237)
                           ;
   U100 : AOI21_X1 port map( B1 => net150934, B2 => net150935, A => net150897, 
                           ZN => n241);
   U101 : INV_X1 port map( A => a(24), ZN => net150902);
   U102 : NAND2_X1 port map( A1 => n106, A2 => a(23), ZN => n252);
   U103 : NAND2_X1 port map( A1 => net150938, A2 => net150882, ZN => n247);
   U104 : INV_X1 port map( A => b(3), ZN => n198);
   U105 : INV_X1 port map( A => b(6), ZN => net152763);
   U106 : NAND2_X1 port map( A1 => n167, A2 => n168, ZN => n174);
   U107 : INV_X1 port map( A => b(10), ZN => n168);
   U108 : INV_X1 port map( A => a(10), ZN => n167);
   U109 : NAND2_X1 port map( A1 => n169, A2 => n170, ZN => n175);
   U110 : INV_X1 port map( A => b(11), ZN => n169);
   U111 : INV_X1 port map( A => a(11), ZN => n170);
   U112 : NAND2_X1 port map( A1 => n156, A2 => n154, ZN => n158);
   U113 : NAND2_X1 port map( A1 => n152, A2 => n153, ZN => n159);
   U114 : OAI211_X1 port map( C1 => n117, C2 => net150953, A => net150951, B =>
                           net150962, ZN => net150961);
   U115 : NAND2_X1 port map( A1 => n251, A2 => n252, ZN => net150953);
   U116 : OAI21_X1 port map( B1 => n235, B2 => net150902, A => net150938, ZN =>
                           net150962);
   U117 : NAND2_X1 port map( A1 => n106, A2 => b(23), ZN => n251);
   U118 : INV_X1 port map( A => a(3), ZN => n204);
   U119 : INV_X1 port map( A => b(7), ZN => n103);
   U120 : NAND2_X1 port map( A1 => a(11), A2 => b(11), ZN => n166);
   U121 : NAND2_X1 port map( A1 => n174, A2 => n175, ZN => n165);
   U122 : INV_X1 port map( A => net150961, ZN => net138479);
   U123 : INV_X1 port map( A => n146, ZN => net152737);
   U124 : AND2_X1 port map( A1 => n136, A2 => n137, ZN => cout(4));
   U125 : NAND2_X1 port map( A1 => net150977, A2 => n255, ZN => n233);
   U126 : NAND2_X1 port map( A1 => net150978, A2 => n256, ZN => n234);
   U127 : OAI21_X1 port map( B1 => net154277, B2 => n165, A => n166, ZN => 
                           cout(2));
   U128 : AND2_X1 port map( A1 => n261, A2 => n260, ZN => n104);
   U129 : NAND2_X1 port map( A1 => n146, A2 => net138535, ZN => n105);
   U130 : AND2_X1 port map( A1 => n244, A2 => n245, ZN => n106);
   U131 : NAND2_X1 port map( A1 => a(0), A2 => b(0), ZN => n109);
   U132 : NOR2_X1 port map( A1 => b(0), A2 => a(0), ZN => n107);
   U133 : OAI21_X1 port map( B1 => n107, B2 => n108, A => n109, ZN => net153553
                           );
   U134 : NOR2_X1 port map( A1 => net153553, A2 => b(1), ZN => net152743);
   U135 : OAI22_X1 port map( A1 => n126, A2 => n117, B1 => a(24), B2 => n114, 
                           ZN => n116);
   U136 : NOR2_X1 port map( A1 => n116, A2 => net150920, ZN => cout(6));
   U137 : NAND2_X1 port map( A1 => n127, A2 => n128, ZN => n126);
   U138 : NAND2_X1 port map( A1 => n130, A2 => n121, ZN => n128);
   U139 : NAND2_X1 port map( A1 => net151486, A2 => n132, ZN => n130);
   U140 : NAND2_X1 port map( A1 => n131, A2 => n123, ZN => n127);
   U141 : NAND2_X1 port map( A1 => n133, A2 => net152653, ZN => n131);
   U142 : OAI211_X1 port map( C1 => n115, C2 => net150922, A => n118, B => n119
                           , ZN => n117);
   U143 : AOI21_X1 port map( B1 => n143, B2 => n136, A => n140, ZN => n142);
   U144 : NOR2_X1 port map( A1 => net154289, A2 => n142, ZN => net153399);
   U145 : NOR2_X1 port map( A1 => net151646, A2 => n142, ZN => net151615);
   U146 : NAND2_X1 port map( A1 => n134, A2 => n144, ZN => n143);
   U147 : NAND2_X1 port map( A1 => n145, A2 => n136, ZN => net151668);
   U148 : NAND2_X1 port map( A1 => net153539, A2 => n141, ZN => n137);
   U149 : NAND2_X1 port map( A1 => net138840, A2 => a(15), ZN => n134);
   U150 : NAND2_X1 port map( A1 => n134, A2 => n82, ZN => n145);
   U151 : OAI21_X1 port map( B1 => net149048, B2 => a(15), A => b(15), ZN => 
                           n144);
   U152 : AND2_X1 port map( A1 => net152678, A2 => n144, ZN => net153539);
   U153 : CLKBUF_X1 port map( A => net138840, Z => n135);
   U154 : NAND2_X1 port map( A1 => net138840, A2 => a(15), ZN => net152678);
   U155 : OAI21_X1 port map( B1 => net149048, B2 => a(15), A => b(15), ZN => 
                           n82);
   U156 : OAI21_X1 port map( B1 => a(15), B2 => n135, A => b(15), ZN => 
                           net138629);
   U157 : OAI221_X1 port map( B1 => n161, B2 => n158, C1 => n163, C2 => n155, A
                           => n159, ZN => n160);
   U158 : AND2_X1 port map( A1 => n160, A2 => net153760, ZN => net154277);
   U159 : AND2_X1 port map( A1 => n160, A2 => net153760, ZN => net153787);
   U160 : NAND2_X1 port map( A1 => n156, A2 => n157, ZN => n155);
   U161 : NAND2_X1 port map( A1 => net153400, A2 => n105, ZN => n162);
   U162 : NAND2_X1 port map( A1 => net153540, A2 => net152799, ZN => n164);
   U163 : NOR2_X1 port map( A1 => n162, A2 => net154049, ZN => n163);
   U164 : NOR2_X1 port map( A1 => net154049, A2 => n162, ZN => n161);
   U165 : NAND2_X1 port map( A1 => n149, A2 => n150, ZN => net153400);
   U166 : AND2_X1 port map( A1 => n148, A2 => net138535, ZN => n150);
   U167 : NAND2_X1 port map( A1 => n148, A2 => net153520, ZN => net152735);
   U168 : NAND2_X1 port map( A1 => n151, A2 => net152783, ZN => n149);
   U169 : AOI21_X1 port map( B1 => net152760, B2 => n147, A => net152747, ZN =>
                           n151);
   U170 : AOI21_X1 port map( B1 => net152760, B2 => n147, A => net152747, ZN =>
                           net152759);
   U171 : OR2_X1 port map( A1 => n102, A2 => n103, ZN => net138535);
   U172 : AND2_X1 port map( A1 => net152763, A2 => net138535, ZN => net152799);
   U173 : AOI21_X1 port map( B1 => n267, B2 => net151647, A => n223, ZN => 
                           net154289);
   U174 : NAND2_X1 port map( A1 => net153401, A2 => b(8), ZN => net154049);
   U175 : NAND2_X1 port map( A1 => n220, A2 => n221, ZN => net151639);
   U176 : NAND3_X1 port map( A1 => a(11), A2 => b(11), A3 => a(12), ZN => n181)
                           ;
   U177 : NAND3_X1 port map( A1 => net138523, A2 => net138522, A3 => n104, ZN 
                           => n185);
   U178 : OAI211_X1 port map( C1 => n179, C2 => n172, A => n184, B => n185, ZN 
                           => n183);
   U179 : INV_X1 port map( A => n183, ZN => net138519);
   U180 : OAI21_X1 port map( B1 => net153787, B2 => n165, A => n182, ZN => n184
                           );
   U181 : NOR2_X1 port map( A1 => net154277, A2 => n173, ZN => n172);
   U182 : NOR2_X1 port map( A1 => a(3), A2 => b(3), ZN => n190);
   U183 : INV_X1 port map( A => a(1), ZN => n202);
   U184 : NAND2_X1 port map( A1 => n202, A2 => net152766, ZN => n207);
   U185 : OAI21_X1 port map( B1 => a(19), B2 => b(19), A => n228, ZN => n221);
   U186 : NOR2_X1 port map( A1 => a(1), A2 => b(1), ZN => n188);
   U187 : NAND2_X1 port map( A1 => n194, A2 => n203, ZN => n208);
   U188 : CLKBUF_X1 port map( A => n200, Z => n186);
   U189 : NAND2_X1 port map( A1 => net152759, A2 => net152783, ZN => net153540)
                           ;
   U190 : CLKBUF_X1 port map( A => net153540, Z => net153520);
   U191 : NAND2_X1 port map( A1 => n196, A2 => n209, ZN => n200);
   U192 : INV_X1 port map( A => n186, ZN => cout(0));
   U193 : NAND2_X1 port map( A1 => net152760, A2 => n206, ZN => net152783);
   U194 : NAND2_X1 port map( A1 => n200, A2 => n205, ZN => n210);
   U195 : AOI21_X1 port map( B1 => n200, B2 => n201, A => n191, ZN => n199);
   U196 : NAND2_X1 port map( A1 => n197, A2 => n204, ZN => n209);
   U197 : AOI21_X1 port map( B1 => n197, B2 => n198, A => n190, ZN => n196);
   U198 : NAND2_X1 port map( A1 => n199, A2 => n210, ZN => net152760);
   U199 : NAND2_X1 port map( A1 => n192, A2 => n207, ZN => n194);
   U200 : NAND2_X1 port map( A1 => net152763, A2 => net153520, ZN => n187);
   U201 : NOR2_X1 port map( A1 => n188, A2 => net152743, ZN => n192);
   U202 : NAND2_X1 port map( A1 => net153540, A2 => net152799, ZN => net153401)
                           ;
   U203 : NAND2_X1 port map( A1 => n193, A2 => n208, ZN => n197);
   U204 : AOI21_X1 port map( B1 => n194, B2 => n195, A => n189, ZN => n193);
   U205 : INV_X1 port map( A => a(2), ZN => n203);
   U206 : NOR2_X1 port map( A1 => a(2), A2 => b(2), ZN => n189);
   U207 : INV_X1 port map( A => net153553, ZN => net152766);
   U208 : NAND2_X1 port map( A1 => net153399, A2 => n212, ZN => net152653);
   U209 : CLKBUF_X1 port map( A => net152653, Z => net152639);
   U210 : NAND2_X1 port map( A1 => net151615, A2 => n212, ZN => net151486);
   U211 : OAI211_X1 port map( C1 => n222, C2 => n225, A => n232, B => n212, ZN 
                           => n211);
   U212 : OAI211_X1 port map( C1 => n222, C2 => n225, A => n232, B => n212, ZN 
                           => n213);
   U213 : NAND4_X1 port map( A1 => n230, A2 => n229, A3 => n231, A4 => n79, ZN 
                           => net151669);
   U214 : INV_X1 port map( A => n69, ZN => n228);
   U215 : NAND2_X1 port map( A1 => n211, A2 => net150984, ZN => net150977);
   U216 : NAND2_X1 port map( A1 => n211, A2 => net150985, ZN => net150978);
   U217 : NAND2_X1 port map( A1 => n213, A2 => net150986, ZN => net150981);
   U218 : NOR2_X1 port map( A1 => net153539, A2 => net151645, ZN => n222);
   U219 : NAND2_X1 port map( A1 => net151667, A2 => net151668, ZN => n232);
   U220 : AOI21_X1 port map( B1 => n267, B2 => net151647, A => n223, ZN => 
                           net151646);
   U221 : INV_X1 port map( A => net151645, ZN => net151647);
   U222 : NAND2_X1 port map( A1 => n249, A2 => n250, ZN => n248);
   U223 : NAND2_X1 port map( A1 => net150981, A2 => n255, ZN => n250);
   U224 : NAND2_X1 port map( A1 => n257, A2 => n256, ZN => n249);
   U225 : INV_X1 port map( A => net152639, ZN => net150897);
   U226 : NAND2_X1 port map( A1 => n259, A2 => net152639, ZN => n245);
   U227 : NAND2_X1 port map( A1 => net151486, A2 => n258, ZN => n257);
   U228 : OAI21_X1 port map( B1 => n248, B2 => n247, A => net150951, ZN => 
                           net150920);
   U229 : CLKBUF_X1 port map( A => net152678, Z => net150785);
   U230 : OR2_X1 port map( A1 => n264, A2 => n265, ZN => n260);
   U231 : OR2_X1 port map( A1 => net138522, A2 => net138523, ZN => n261);
   U232 : AND2_X1 port map( A1 => net138519, A2 => n262, ZN => net149048);
   U233 : INV_X1 port map( A => a(17), ZN => n76);
   U234 : NAND2_X1 port map( A1 => n77, A2 => n76, ZN => n79);
   U235 : OAI21_X1 port map( B1 => n36, B2 => n37, A => n38, ZN => cout(7));
   U236 : INV_X1 port map( A => a(31), ZN => n37);
   U237 : INV_X1 port map( A => b(14), ZN => n265);
   U238 : OAI21_X1 port map( B1 => a(18), B2 => n73, A => n74, ZN => n69);
   U239 : INV_X1 port map( A => n75, ZN => n74);
   U240 : AOI21_X1 port map( B1 => n73, B2 => a(18), A => b(18), ZN => n75);
   U241 : OAI21_X1 port map( B1 => n76, B2 => n77, A => n78, ZN => n73);
   U242 : OAI21_X1 port map( B1 => n42, B2 => n43, A => n44, ZN => n40);
   U243 : INV_X1 port map( A => b(29), ZN => n43);
   U244 : OAI21_X1 port map( B1 => n39, B2 => a(31), A => b(31), ZN => n38);
   U245 : INV_X1 port map( A => n36, ZN => n39);
   U246 : INV_X1 port map( A => b(17), ZN => n77);
   U247 : INV_X1 port map( A => a(29), ZN => n42);
   U248 : AND2_X1 port map( A1 => n40, A2 => a(30), ZN => n41);
   U249 : OAI22_X1 port map( A1 => a(30), A2 => n40, B1 => b(30), B2 => n41, ZN
                           => n36);
   U250 : INV_X1 port map( A => a(14), ZN => n264);
   U251 : AND2_X1 port map( A1 => net138519, A2 => n262, ZN => net138840);
   U252 : OR2_X1 port map( A1 => b(14), A2 => a(14), ZN => n262);
   U253 : NAND2_X1 port map( A1 => net138629, A2 => net150785, ZN => cout(3));
   U254 : NAND2_X1 port map( A1 => net152678, A2 => n82, ZN => n267);
   U255 : OAI21_X1 port map( B1 => n102, B2 => n103, A => net138537, ZN => 
                           cout(1));
   U256 : OAI222_X1 port map( A1 => a(28), A2 => net138479, B1 => b(28), B2 => 
                           n45, C1 => b(29), C2 => a(29), ZN => n44);
   U257 : AND2_X1 port map( A1 => net138479, A2 => a(28), ZN => n45);

end SYN_p4_carry_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Div_DATA_SIZE32_DIV_STAGE34_SQRT_STAGE18_DW01_inc_0 is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end Div_DATA_SIZE32_DIV_STAGE34_SQRT_STAGE18_DW01_inc_0;

architecture SYN_rpl of Div_DATA_SIZE32_DIV_STAGE34_SQRT_STAGE18_DW01_inc_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port : std_logic;

begin
   
   U1_1_30 : HA_X1 port map( A => A(30), B => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_1_29 : HA_X1 port map( A => A(29), B => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_1_28 : HA_X1 port map( A => A(28), B => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_1_27 : HA_X1 port map( A => A(27), B => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_1_26 : HA_X1 port map( A => A(26), B => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_1_25 : HA_X1 port map( A => A(25), B => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_1_24 : HA_X1 port map( A => A(24), B => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_1_23 : HA_X1 port map( A => A(23), B => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_1_22 : HA_X1 port map( A => A(22), B => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_1_21 : HA_X1 port map( A => A(21), B => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_1_20 : HA_X1 port map( A => A(20), B => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_1_19 : HA_X1 port map( A => A(19), B => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_1_18 : HA_X1 port map( A => A(18), B => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_1_17 : HA_X1 port map( A => A(17), B => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_1_16 : HA_X1 port map( A => A(16), B => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_1_15 : HA_X1 port map( A => A(15), B => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : XOR2_X1 port map( A => carry_31_port, B => A(31), Z => SUM(31));
   U2 : INV_X1 port map( A => A(0), ZN => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Sipo_DATA_SIZE32 is

   port( rst, en, clk, din : in std_logic;  dout : out std_logic_vector (31 
         downto 0));

end Sipo_DATA_SIZE32;

architecture SYN_sipo_arch of Sipo_DATA_SIZE32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
      n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n65, n66, n67
      , n68, n69, n70, net108809, net108810, net108811, net108812, net108813, 
      net108814, net108815, net108816, net108817, net108818, net108819, 
      net108820, net108821, net108822, net108823, net108824, net108825, 
      net108826, net108827, net108828, net108829, net108830, net108831, 
      net108832, net108833, net108834, net108835, net108836, net108837, 
      net108838, net108839, net108840, n38, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, net164139, net164140, net164141, net164142, net164143, 
      net164144, net164145, net164146, net164147, net164148, net164149, 
      net164150, net164151, net164152, net164153, net164154, net164155, 
      net164156, net164157, net164158, net164159, net164160, net164161, 
      net164162, net164163, net164164, net164165, net164166, net164167, 
      net164168 : std_logic;

begin
   
   dout_reg_1_inst : DFFR_X1 port map( D => n161, CK => clk, RN => n84, Q => 
                           dout(1), QN => net108839);
   data_reg_2_inst : DFF_X1 port map( D => n160, CK => clk, Q => net164168, QN 
                           => n69);
   dout_reg_2_inst : DFFR_X1 port map( D => n159, CK => clk, RN => n84, Q => 
                           dout(2), QN => net108838);
   data_reg_3_inst : DFF_X1 port map( D => n158, CK => clk, Q => net164167, QN 
                           => n68);
   dout_reg_3_inst : DFFR_X1 port map( D => n157, CK => clk, RN => n84, Q => 
                           dout(3), QN => net108837);
   data_reg_4_inst : DFF_X1 port map( D => n156, CK => clk, Q => net164166, QN 
                           => n67);
   dout_reg_4_inst : DFFR_X1 port map( D => n155, CK => clk, RN => n84, Q => 
                           dout(4), QN => net108836);
   data_reg_5_inst : DFF_X1 port map( D => n154, CK => clk, Q => net164165, QN 
                           => n66);
   dout_reg_5_inst : DFFR_X1 port map( D => n153, CK => clk, RN => n84, Q => 
                           dout(5), QN => net108835);
   data_reg_6_inst : DFF_X1 port map( D => n152, CK => clk, Q => net164164, QN 
                           => n65);
   dout_reg_6_inst : DFFR_X1 port map( D => n151, CK => clk, RN => n84, Q => 
                           dout(6), QN => net108834);
   data_reg_7_inst : DFF_X1 port map( D => n150, CK => clk, Q => net164163, QN 
                           => n74);
   dout_reg_7_inst : DFFR_X1 port map( D => n149, CK => clk, RN => n84, Q => 
                           dout(7), QN => net108833);
   data_reg_8_inst : DFF_X1 port map( D => n148, CK => clk, Q => net164162, QN 
                           => n72);
   dout_reg_8_inst : DFFR_X1 port map( D => n147, CK => clk, RN => n84, Q => 
                           dout(8), QN => net108832);
   data_reg_9_inst : DFF_X1 port map( D => n146, CK => clk, Q => net164161, QN 
                           => n73);
   dout_reg_9_inst : DFFR_X1 port map( D => n145, CK => clk, RN => n84, Q => 
                           dout(9), QN => net108831);
   data_reg_10_inst : DFF_X1 port map( D => n144, CK => clk, Q => net164160, QN
                           => n61);
   dout_reg_10_inst : DFFR_X1 port map( D => n143, CK => clk, RN => n84, Q => 
                           dout(10), QN => net108830);
   data_reg_11_inst : DFF_X1 port map( D => n142, CK => clk, Q => net164159, QN
                           => n60);
   dout_reg_11_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n84, Q => 
                           dout(11), QN => net108829);
   data_reg_12_inst : DFF_X1 port map( D => n140, CK => clk, Q => net164158, QN
                           => n59);
   dout_reg_12_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n84, Q => 
                           dout(12), QN => net108828);
   data_reg_13_inst : DFF_X1 port map( D => n138, CK => clk, Q => net164157, QN
                           => n58);
   dout_reg_13_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n84, Q => 
                           dout(13), QN => net108827);
   data_reg_14_inst : DFF_X1 port map( D => n136, CK => clk, Q => net164156, QN
                           => n57);
   dout_reg_14_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n84, Q => 
                           dout(14), QN => net108826);
   data_reg_15_inst : DFF_X1 port map( D => n134, CK => clk, Q => net164155, QN
                           => n56);
   dout_reg_15_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n84, Q => 
                           dout(15), QN => net108825);
   data_reg_16_inst : DFF_X1 port map( D => n132, CK => clk, Q => net164154, QN
                           => n55);
   dout_reg_16_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n84, Q => 
                           dout(16), QN => net108824);
   data_reg_17_inst : DFF_X1 port map( D => n130, CK => clk, Q => net164153, QN
                           => n54);
   dout_reg_17_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n83, Q => 
                           dout(17), QN => net108823);
   data_reg_18_inst : DFF_X1 port map( D => n128, CK => clk, Q => net164152, QN
                           => n53);
   dout_reg_18_inst : DFFR_X1 port map( D => n127, CK => clk, RN => n83, Q => 
                           dout(18), QN => net108822);
   data_reg_19_inst : DFF_X1 port map( D => n126, CK => clk, Q => net164151, QN
                           => n52);
   dout_reg_19_inst : DFFR_X1 port map( D => n125, CK => clk, RN => n83, Q => 
                           dout(19), QN => net108821);
   data_reg_20_inst : DFF_X1 port map( D => n124, CK => clk, Q => net164150, QN
                           => n51);
   dout_reg_20_inst : DFFR_X1 port map( D => n123, CK => clk, RN => n83, Q => 
                           dout(20), QN => net108820);
   data_reg_21_inst : DFF_X1 port map( D => n122, CK => clk, Q => net164149, QN
                           => n50);
   dout_reg_21_inst : DFFR_X1 port map( D => n121, CK => clk, RN => n83, Q => 
                           dout(21), QN => net108819);
   data_reg_22_inst : DFF_X1 port map( D => n120, CK => clk, Q => net164148, QN
                           => n49);
   dout_reg_22_inst : DFFR_X1 port map( D => n119, CK => clk, RN => n83, Q => 
                           dout(22), QN => net108818);
   data_reg_23_inst : DFF_X1 port map( D => n118, CK => clk, Q => net164147, QN
                           => n48);
   dout_reg_23_inst : DFFR_X1 port map( D => n117, CK => clk, RN => n83, Q => 
                           dout(23), QN => net108817);
   data_reg_24_inst : DFF_X1 port map( D => n116, CK => clk, Q => net164146, QN
                           => n47);
   dout_reg_24_inst : DFFR_X1 port map( D => n115, CK => clk, RN => n83, Q => 
                           dout(24), QN => net108816);
   data_reg_25_inst : DFF_X1 port map( D => n114, CK => clk, Q => net164145, QN
                           => n46);
   dout_reg_25_inst : DFFR_X1 port map( D => n113, CK => clk, RN => n83, Q => 
                           dout(25), QN => net108815);
   data_reg_26_inst : DFF_X1 port map( D => n112, CK => clk, Q => net164144, QN
                           => n45);
   dout_reg_26_inst : DFFR_X1 port map( D => n111, CK => clk, RN => n83, Q => 
                           dout(26), QN => net108814);
   data_reg_27_inst : DFF_X1 port map( D => n110, CK => clk, Q => net164143, QN
                           => n44);
   dout_reg_27_inst : DFFR_X1 port map( D => n109, CK => clk, RN => n83, Q => 
                           dout(27), QN => net108813);
   data_reg_28_inst : DFF_X1 port map( D => n108, CK => clk, Q => net164142, QN
                           => n43);
   dout_reg_28_inst : DFFR_X1 port map( D => n107, CK => clk, RN => n83, Q => 
                           dout(28), QN => net108812);
   data_reg_29_inst : DFF_X1 port map( D => n106, CK => clk, Q => net164141, QN
                           => n42);
   dout_reg_29_inst : DFFR_X1 port map( D => n105, CK => clk, RN => n83, Q => 
                           dout(29), QN => net108811);
   data_reg_30_inst : DFF_X1 port map( D => n104, CK => clk, Q => net164140, QN
                           => n41);
   dout_reg_30_inst : DFFR_X1 port map( D => n103, CK => clk, RN => n83, Q => 
                           dout(30), QN => net108810);
   data_reg_31_inst : DFF_X1 port map( D => n102, CK => clk, Q => net164139, QN
                           => n40);
   dout_reg_31_inst : DFFR_X1 port map( D => n101, CK => clk, RN => n83, Q => 
                           dout(31), QN => net108809);
   dout_reg_0_inst : DFFR_X1 port map( D => n163, CK => clk, RN => n84, Q => 
                           dout(0), QN => net108840);
   data_reg_1_inst : DFF_X1 port map( D => n162, CK => clk, Q => n71, QN => n70
                           );
   U3 : OR2_X1 port map( A1 => n82, A2 => n70, ZN => n75);
   U4 : NAND2_X1 port map( A1 => n95, A2 => n75, ZN => n162);
   U5 : INV_X1 port map( A => n76, ZN => n78);
   U6 : BUF_X1 port map( A => n38, Z => n81);
   U7 : BUF_X1 port map( A => n38, Z => n80);
   U8 : BUF_X1 port map( A => n38, Z => n82);
   U9 : NAND2_X1 port map( A1 => n83, A2 => n86, ZN => n38);
   U10 : BUF_X1 port map( A => n94, Z => n93);
   U11 : AND2_X1 port map( A1 => n83, A2 => en, ZN => n76);
   U12 : BUF_X1 port map( A => n94, Z => n86);
   U13 : BUF_X1 port map( A => n94, Z => n87);
   U14 : BUF_X1 port map( A => n94, Z => n88);
   U15 : BUF_X1 port map( A => n88, Z => n89);
   U16 : BUF_X1 port map( A => n88, Z => n90);
   U17 : BUF_X1 port map( A => n88, Z => n91);
   U18 : BUF_X1 port map( A => n88, Z => n92);
   U19 : BUF_X1 port map( A => rst, Z => n83);
   U20 : INV_X1 port map( A => n85, ZN => n94);
   U21 : BUF_X1 port map( A => rst, Z => n84);
   U22 : BUF_X1 port map( A => en, Z => n85);
   U23 : OAI22_X1 port map( A1 => n82, A2 => n73, B1 => n79, B2 => n72, ZN => 
                           n146);
   U24 : OAI22_X1 port map( A1 => n82, A2 => n72, B1 => n79, B2 => n74, ZN => 
                           n148);
   U25 : OAI22_X1 port map( A1 => n40, A2 => n90, B1 => net108809, B2 => n85, 
                           ZN => n101);
   U26 : OAI22_X1 port map( A1 => n41, A2 => n86, B1 => net108810, B2 => n85, 
                           ZN => n103);
   U27 : OAI22_X1 port map( A1 => n42, A2 => n86, B1 => net108811, B2 => n85, 
                           ZN => n105);
   U28 : OAI22_X1 port map( A1 => n43, A2 => n86, B1 => net108812, B2 => n85, 
                           ZN => n107);
   U29 : OAI22_X1 port map( A1 => n44, A2 => n87, B1 => net108813, B2 => n85, 
                           ZN => n109);
   U30 : OAI22_X1 port map( A1 => n45, A2 => n87, B1 => net108814, B2 => en, ZN
                           => n111);
   U31 : OAI22_X1 port map( A1 => n46, A2 => n87, B1 => net108815, B2 => n85, 
                           ZN => n113);
   U32 : OAI22_X1 port map( A1 => n47, A2 => n87, B1 => net108816, B2 => n85, 
                           ZN => n115);
   U33 : OAI22_X1 port map( A1 => n61, A2 => n80, B1 => n79, B2 => n73, ZN => 
                           n144);
   U34 : OAI22_X1 port map( A1 => n69, A2 => n80, B1 => n70, B2 => n78, ZN => 
                           n160);
   U35 : OAI22_X1 port map( A1 => n40, A2 => n82, B1 => n41, B2 => n78, ZN => 
                           n102);
   U36 : OAI22_X1 port map( A1 => n41, A2 => n82, B1 => n42, B2 => n78, ZN => 
                           n104);
   U37 : OAI22_X1 port map( A1 => n44, A2 => n81, B1 => n45, B2 => n79, ZN => 
                           n110);
   U38 : OAI22_X1 port map( A1 => n46, A2 => n81, B1 => n47, B2 => n78, ZN => 
                           n114);
   U39 : OAI22_X1 port map( A1 => n47, A2 => n81, B1 => n48, B2 => n79, ZN => 
                           n116);
   U40 : OAI22_X1 port map( A1 => n48, A2 => n81, B1 => n49, B2 => n78, ZN => 
                           n118);
   U41 : OAI22_X1 port map( A1 => n49, A2 => n81, B1 => n50, B2 => n79, ZN => 
                           n120);
   U42 : OAI22_X1 port map( A1 => n50, A2 => n81, B1 => n51, B2 => n79, ZN => 
                           n122);
   U43 : OAI22_X1 port map( A1 => n51, A2 => n81, B1 => n52, B2 => n79, ZN => 
                           n124);
   U44 : OAI22_X1 port map( A1 => n52, A2 => n81, B1 => n53, B2 => n79, ZN => 
                           n126);
   U45 : OAI22_X1 port map( A1 => n53, A2 => n81, B1 => n54, B2 => n79, ZN => 
                           n128);
   U46 : OAI22_X1 port map( A1 => n54, A2 => n80, B1 => n55, B2 => n79, ZN => 
                           n130);
   U47 : OAI22_X1 port map( A1 => n55, A2 => n80, B1 => n56, B2 => n78, ZN => 
                           n132);
   U48 : OAI22_X1 port map( A1 => n56, A2 => n80, B1 => n57, B2 => n78, ZN => 
                           n134);
   U49 : OAI22_X1 port map( A1 => n57, A2 => n80, B1 => n58, B2 => n78, ZN => 
                           n136);
   U50 : OAI22_X1 port map( A1 => n58, A2 => n80, B1 => n59, B2 => n78, ZN => 
                           n138);
   U51 : OAI22_X1 port map( A1 => n59, A2 => n80, B1 => n60, B2 => n78, ZN => 
                           n140);
   U52 : OAI22_X1 port map( A1 => n60, A2 => n80, B1 => n61, B2 => n78, ZN => 
                           n142);
   U53 : OAI22_X1 port map( A1 => n82, A2 => n74, B1 => n65, B2 => n78, ZN => 
                           n150);
   U54 : OAI22_X1 port map( A1 => n65, A2 => n80, B1 => n66, B2 => n78, ZN => 
                           n152);
   U55 : OAI22_X1 port map( A1 => n66, A2 => n81, B1 => n67, B2 => n79, ZN => 
                           n154);
   U56 : OAI22_X1 port map( A1 => n67, A2 => n80, B1 => n68, B2 => n78, ZN => 
                           n156);
   U57 : OAI22_X1 port map( A1 => n68, A2 => n80, B1 => n69, B2 => n78, ZN => 
                           n158);
   U58 : OAI22_X1 port map( A1 => n59, A2 => n91, B1 => net108828, B2 => en, ZN
                           => n139);
   U59 : OAI22_X1 port map( A1 => n60, A2 => n91, B1 => net108829, B2 => en, ZN
                           => n141);
   U60 : OAI22_X1 port map( A1 => n61, A2 => n91, B1 => net108830, B2 => en, ZN
                           => n143);
   U61 : OAI22_X1 port map( A1 => n93, A2 => n73, B1 => net108831, B2 => n85, 
                           ZN => n145);
   U62 : OAI22_X1 port map( A1 => n93, A2 => n72, B1 => net108832, B2 => n85, 
                           ZN => n147);
   U63 : OAI22_X1 port map( A1 => n93, A2 => n74, B1 => net108833, B2 => n85, 
                           ZN => n149);
   U64 : OAI22_X1 port map( A1 => n65, A2 => n92, B1 => net108834, B2 => n85, 
                           ZN => n151);
   U65 : OAI22_X1 port map( A1 => n66, A2 => n92, B1 => net108835, B2 => en, ZN
                           => n153);
   U66 : OAI22_X1 port map( A1 => n67, A2 => n91, B1 => net108836, B2 => n85, 
                           ZN => n155);
   U67 : OAI22_X1 port map( A1 => n68, A2 => n92, B1 => net108837, B2 => en, ZN
                           => n157);
   U68 : OAI22_X1 port map( A1 => n69, A2 => n93, B1 => net108838, B2 => en, ZN
                           => n159);
   U69 : OAI22_X1 port map( A1 => n42, A2 => n81, B1 => n43, B2 => n79, ZN => 
                           n106);
   U70 : OAI22_X1 port map( A1 => n43, A2 => n82, B1 => n44, B2 => n79, ZN => 
                           n108);
   U71 : OAI22_X1 port map( A1 => n45, A2 => n81, B1 => n46, B2 => n79, ZN => 
                           n112);
   U72 : OAI22_X1 port map( A1 => n48, A2 => n88, B1 => net108817, B2 => n85, 
                           ZN => n117);
   U73 : OAI22_X1 port map( A1 => n49, A2 => n88, B1 => net108818, B2 => n85, 
                           ZN => n119);
   U74 : OAI22_X1 port map( A1 => n50, A2 => n88, B1 => net108819, B2 => en, ZN
                           => n121);
   U75 : OAI22_X1 port map( A1 => n51, A2 => n88, B1 => net108820, B2 => en, ZN
                           => n123);
   U76 : OAI22_X1 port map( A1 => n52, A2 => n89, B1 => net108821, B2 => en, ZN
                           => n125);
   U77 : OAI22_X1 port map( A1 => n53, A2 => n89, B1 => net108822, B2 => en, ZN
                           => n127);
   U78 : OAI22_X1 port map( A1 => n54, A2 => n89, B1 => net108823, B2 => en, ZN
                           => n129);
   U79 : OAI22_X1 port map( A1 => n55, A2 => n89, B1 => net108824, B2 => en, ZN
                           => n131);
   U80 : OAI22_X1 port map( A1 => n56, A2 => n90, B1 => net108825, B2 => n85, 
                           ZN => n133);
   U81 : OAI22_X1 port map( A1 => n57, A2 => n90, B1 => net108826, B2 => en, ZN
                           => n135);
   U82 : OAI22_X1 port map( A1 => n58, A2 => n90, B1 => net108827, B2 => n85, 
                           ZN => n137);
   U83 : OAI22_X1 port map( A1 => n70, A2 => n92, B1 => net108839, B2 => n85, 
                           ZN => n161);
   U84 : OR2_X1 port map( A1 => en, A2 => net108840, ZN => n77);
   U85 : NAND2_X1 port map( A1 => n95, A2 => n77, ZN => n163);
   U86 : NAND2_X1 port map( A1 => din, A2 => n76, ZN => n95);
   U87 : INV_X1 port map( A => n76, ZN => n79);

end SYN_sipo_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE64 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (63 downto 0);
         dout : out std_logic_vector (63 downto 0));

end Reg_DATA_SIZE64;

architecture SYN_reg_arch of Reg_DATA_SIZE64 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal dout_59_port, dout_58_port, dout_57_port, dout_56_port, dout_55_port,
      dout_54_port, dout_53_port, dout_52_port, dout_51_port, dout_50_port, 
      dout_49_port, dout_48_port, dout_47_port, dout_46_port, dout_45_port, 
      dout_44_port, dout_43_port, dout_42_port, dout_41_port, dout_40_port, 
      dout_39_port, dout_38_port, dout_37_port, dout_36_port, dout_35_port, 
      dout_34_port, dout_33_port, dout_32_port, dout_31_port, dout_30_port, 
      dout_29_port, dout_28_port, dout_27_port, dout_26_port, dout_25_port, 
      dout_24_port, dout_23_port, dout_22_port, dout_21_port, dout_20_port, 
      dout_19_port, dout_18_port, dout_17_port, dout_16_port, dout_15_port, 
      dout_14_port, dout_13_port, dout_12_port, dout_11_port, dout_10_port, 
      dout_9_port, dout_8_port, dout_7_port, dout_6_port, dout_5_port, 
      dout_4_port, dout_3_port, dout_2_port, dout_1_port, dout_0_port, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, 
      n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, 
      n190, n191, n192, net108745, net108746, net108747, net108748, net108749, 
      net108750, net108751, net108752, net108753, net108754, net108755, 
      net108756, net108757, net108758, net108759, net108760, net108761, 
      net108762, net108763, net108764, net108765, net108766, net108767, 
      net108768, net108769, net108770, net108771, net108772, net108773, 
      net108774, net108775, net108776, net108777, net108778, net108779, 
      net108780, net108781, net108782, net108783, net108784, net108785, 
      net108786, net108787, net108788, net108789, net108790, net108791, 
      net108792, net108793, net108794, net108795, net108796, net108797, 
      net108798, net108799, net108800, net108801, net108802, net108803, 
      net108804, net108805, net108806, net108807, net108808, n17, n18, n19, n20
      , n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, 
      n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49
      , n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, 
      n64, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n65, n66, n67, n68, 
      n69, n70, n71, n72, dout_60_port, dout_61_port, dout_62_port, 
      dout_63_port : std_logic;

begin
   dout <= ( dout_63_port, dout_62_port, dout_61_port, dout_60_port, 
      dout_59_port, dout_58_port, dout_57_port, dout_56_port, dout_55_port, 
      dout_54_port, dout_53_port, dout_52_port, dout_51_port, dout_50_port, 
      dout_49_port, dout_48_port, dout_47_port, dout_46_port, dout_45_port, 
      dout_44_port, dout_43_port, dout_42_port, dout_41_port, dout_40_port, 
      dout_39_port, dout_38_port, dout_37_port, dout_36_port, dout_35_port, 
      dout_34_port, dout_33_port, dout_32_port, dout_31_port, dout_30_port, 
      dout_29_port, dout_28_port, dout_27_port, dout_26_port, dout_25_port, 
      dout_24_port, dout_23_port, dout_22_port, dout_21_port, dout_20_port, 
      dout_19_port, dout_18_port, dout_17_port, dout_16_port, dout_15_port, 
      dout_14_port, dout_13_port, dout_12_port, dout_11_port, dout_10_port, 
      dout_9_port, dout_8_port, dout_7_port, dout_6_port, dout_5_port, 
      dout_4_port, dout_3_port, dout_2_port, dout_1_port, dout_0_port );
   
   dout_reg_63_inst : DFFR_X1 port map( D => n192, CK => clk, RN => n11, Q => 
                           dout_63_port, QN => net108808);
   dout_reg_62_inst : DFFR_X1 port map( D => n191, CK => clk, RN => n12, Q => 
                           dout_62_port, QN => net108807);
   dout_reg_61_inst : DFFR_X1 port map( D => n190, CK => clk, RN => n12, Q => 
                           dout_61_port, QN => net108806);
   dout_reg_60_inst : DFFR_X1 port map( D => n189, CK => clk, RN => n12, Q => 
                           dout_60_port, QN => net108805);
   dout_reg_59_inst : DFFR_X1 port map( D => n188, CK => clk, RN => n7, Q => 
                           dout_59_port, QN => net108804);
   dout_reg_58_inst : DFFR_X1 port map( D => n187, CK => clk, RN => n7, Q => 
                           dout_58_port, QN => net108803);
   dout_reg_57_inst : DFFR_X1 port map( D => n186, CK => clk, RN => n7, Q => 
                           dout_57_port, QN => net108802);
   dout_reg_56_inst : DFFR_X1 port map( D => n185, CK => clk, RN => n7, Q => 
                           dout_56_port, QN => net108801);
   dout_reg_55_inst : DFFR_X1 port map( D => n184, CK => clk, RN => n7, Q => 
                           dout_55_port, QN => net108800);
   dout_reg_54_inst : DFFR_X1 port map( D => n183, CK => clk, RN => n7, Q => 
                           dout_54_port, QN => net108799);
   dout_reg_53_inst : DFFR_X1 port map( D => n182, CK => clk, RN => n7, Q => 
                           dout_53_port, QN => net108798);
   dout_reg_52_inst : DFFR_X1 port map( D => n181, CK => clk, RN => n7, Q => 
                           dout_52_port, QN => net108797);
   dout_reg_51_inst : DFFR_X1 port map( D => n180, CK => clk, RN => n7, Q => 
                           dout_51_port, QN => net108796);
   dout_reg_50_inst : DFFR_X1 port map( D => n179, CK => clk, RN => n7, Q => 
                           dout_50_port, QN => net108795);
   dout_reg_49_inst : DFFR_X1 port map( D => n178, CK => clk, RN => n7, Q => 
                           dout_49_port, QN => net108794);
   dout_reg_48_inst : DFFR_X1 port map( D => n177, CK => clk, RN => n7, Q => 
                           dout_48_port, QN => net108793);
   dout_reg_47_inst : DFFR_X1 port map( D => n176, CK => clk, RN => n8, Q => 
                           dout_47_port, QN => net108792);
   dout_reg_46_inst : DFFR_X1 port map( D => n175, CK => clk, RN => n8, Q => 
                           dout_46_port, QN => net108791);
   dout_reg_45_inst : DFFR_X1 port map( D => n174, CK => clk, RN => n8, Q => 
                           dout_45_port, QN => net108790);
   dout_reg_44_inst : DFFR_X1 port map( D => n173, CK => clk, RN => n8, Q => 
                           dout_44_port, QN => net108789);
   dout_reg_43_inst : DFFR_X1 port map( D => n172, CK => clk, RN => n8, Q => 
                           dout_43_port, QN => net108788);
   dout_reg_42_inst : DFFR_X1 port map( D => n171, CK => clk, RN => n8, Q => 
                           dout_42_port, QN => net108787);
   dout_reg_41_inst : DFFR_X1 port map( D => n170, CK => clk, RN => n8, Q => 
                           dout_41_port, QN => net108786);
   dout_reg_40_inst : DFFR_X1 port map( D => n169, CK => clk, RN => n12, Q => 
                           dout_40_port, QN => net108785);
   dout_reg_39_inst : DFFR_X1 port map( D => n168, CK => clk, RN => n8, Q => 
                           dout_39_port, QN => net108784);
   dout_reg_38_inst : DFFR_X1 port map( D => n167, CK => clk, RN => n8, Q => 
                           dout_38_port, QN => net108783);
   dout_reg_37_inst : DFFR_X1 port map( D => n166, CK => clk, RN => n8, Q => 
                           dout_37_port, QN => net108782);
   dout_reg_36_inst : DFFR_X1 port map( D => n165, CK => clk, RN => n8, Q => 
                           dout_36_port, QN => net108781);
   dout_reg_35_inst : DFFR_X1 port map( D => n164, CK => clk, RN => n8, Q => 
                           dout_35_port, QN => net108780);
   dout_reg_34_inst : DFFR_X1 port map( D => n163, CK => clk, RN => n9, Q => 
                           dout_34_port, QN => net108779);
   dout_reg_33_inst : DFFR_X1 port map( D => n162, CK => clk, RN => n9, Q => 
                           dout_33_port, QN => net108778);
   dout_reg_32_inst : DFFR_X1 port map( D => n161, CK => clk, RN => n9, Q => 
                           dout_32_port, QN => net108777);
   dout_reg_31_inst : DFFR_X1 port map( D => n160, CK => clk, RN => n9, Q => 
                           dout_31_port, QN => net108776);
   dout_reg_30_inst : DFFR_X1 port map( D => n159, CK => clk, RN => n9, Q => 
                           dout_30_port, QN => net108775);
   dout_reg_29_inst : DFFR_X1 port map( D => n158, CK => clk, RN => n9, Q => 
                           dout_29_port, QN => net108774);
   dout_reg_28_inst : DFFR_X1 port map( D => n157, CK => clk, RN => n9, Q => 
                           dout_28_port, QN => net108773);
   dout_reg_27_inst : DFFR_X1 port map( D => n156, CK => clk, RN => n9, Q => 
                           dout_27_port, QN => net108772);
   dout_reg_26_inst : DFFR_X1 port map( D => n155, CK => clk, RN => n9, Q => 
                           dout_26_port, QN => net108771);
   dout_reg_25_inst : DFFR_X1 port map( D => n154, CK => clk, RN => n9, Q => 
                           dout_25_port, QN => net108770);
   dout_reg_24_inst : DFFR_X1 port map( D => n153, CK => clk, RN => n9, Q => 
                           dout_24_port, QN => net108769);
   dout_reg_23_inst : DFFR_X1 port map( D => n152, CK => clk, RN => n9, Q => 
                           dout_23_port, QN => net108768);
   dout_reg_22_inst : DFFR_X1 port map( D => n151, CK => clk, RN => n10, Q => 
                           dout_22_port, QN => net108767);
   dout_reg_21_inst : DFFR_X1 port map( D => n150, CK => clk, RN => n10, Q => 
                           dout_21_port, QN => net108766);
   dout_reg_20_inst : DFFR_X1 port map( D => n149, CK => clk, RN => n10, Q => 
                           dout_20_port, QN => net108765);
   dout_reg_19_inst : DFFR_X1 port map( D => n148, CK => clk, RN => n10, Q => 
                           dout_19_port, QN => net108764);
   dout_reg_18_inst : DFFR_X1 port map( D => n147, CK => clk, RN => n10, Q => 
                           dout_18_port, QN => net108763);
   dout_reg_17_inst : DFFR_X1 port map( D => n146, CK => clk, RN => n10, Q => 
                           dout_17_port, QN => net108762);
   dout_reg_16_inst : DFFR_X1 port map( D => n145, CK => clk, RN => n10, Q => 
                           dout_16_port, QN => net108761);
   dout_reg_15_inst : DFFR_X1 port map( D => n144, CK => clk, RN => n10, Q => 
                           dout_15_port, QN => net108760);
   dout_reg_14_inst : DFFR_X1 port map( D => n143, CK => clk, RN => n10, Q => 
                           dout_14_port, QN => net108759);
   dout_reg_13_inst : DFFR_X1 port map( D => n142, CK => clk, RN => n10, Q => 
                           dout_13_port, QN => net108758);
   dout_reg_12_inst : DFFR_X1 port map( D => n141, CK => clk, RN => n10, Q => 
                           dout_12_port, QN => net108757);
   dout_reg_11_inst : DFFR_X1 port map( D => n140, CK => clk, RN => n10, Q => 
                           dout_11_port, QN => net108756);
   dout_reg_10_inst : DFFR_X1 port map( D => n139, CK => clk, RN => n11, Q => 
                           dout_10_port, QN => net108755);
   dout_reg_9_inst : DFFR_X1 port map( D => n138, CK => clk, RN => n11, Q => 
                           dout_9_port, QN => net108754);
   dout_reg_8_inst : DFFR_X1 port map( D => n137, CK => clk, RN => n11, Q => 
                           dout_8_port, QN => net108753);
   dout_reg_7_inst : DFFR_X1 port map( D => n136, CK => clk, RN => n11, Q => 
                           dout_7_port, QN => net108752);
   dout_reg_6_inst : DFFR_X1 port map( D => n135, CK => clk, RN => n11, Q => 
                           dout_6_port, QN => net108751);
   dout_reg_5_inst : DFFR_X1 port map( D => n134, CK => clk, RN => n11, Q => 
                           dout_5_port, QN => net108750);
   dout_reg_4_inst : DFFR_X1 port map( D => n133, CK => clk, RN => n11, Q => 
                           dout_4_port, QN => net108749);
   dout_reg_3_inst : DFFR_X1 port map( D => n132, CK => clk, RN => n11, Q => 
                           dout_3_port, QN => net108748);
   dout_reg_2_inst : DFFR_X1 port map( D => n131, CK => clk, RN => n11, Q => 
                           dout_2_port, QN => net108747);
   dout_reg_1_inst : DFFR_X1 port map( D => n130, CK => clk, RN => n11, Q => 
                           dout_1_port, QN => net108746);
   dout_reg_0_inst : DFFR_X1 port map( D => n129, CK => clk, RN => n11, Q => 
                           dout_0_port, QN => net108745);
   U2 : BUF_X1 port map( A => n14, Z => n67);
   U3 : BUF_X1 port map( A => n13, Z => n66);
   U4 : BUF_X1 port map( A => n13, Z => n65);
   U5 : BUF_X1 port map( A => n13, Z => n16);
   U6 : BUF_X1 port map( A => n15, Z => n71);
   U7 : BUF_X1 port map( A => n14, Z => n69);
   U8 : BUF_X1 port map( A => n14, Z => n68);
   U9 : BUF_X1 port map( A => n15, Z => n70);
   U10 : BUF_X1 port map( A => n15, Z => n72);
   U11 : OAI21_X1 port map( B1 => net108777, B2 => n69, A => n32, ZN => n161);
   U12 : NAND2_X1 port map( A1 => din(32), A2 => n66, ZN => n32);
   U13 : OAI21_X1 port map( B1 => net108778, B2 => n68, A => n31, ZN => n162);
   U14 : NAND2_X1 port map( A1 => din(33), A2 => n66, ZN => n31);
   U15 : OAI21_X1 port map( B1 => net108779, B2 => n68, A => n30, ZN => n163);
   U16 : NAND2_X1 port map( A1 => din(34), A2 => n66, ZN => n30);
   U17 : OAI21_X1 port map( B1 => net108780, B2 => n68, A => n29, ZN => n164);
   U18 : NAND2_X1 port map( A1 => din(35), A2 => n65, ZN => n29);
   U19 : OAI21_X1 port map( B1 => net108789, B2 => n68, A => n20, ZN => n173);
   U20 : NAND2_X1 port map( A1 => din(44), A2 => n16, ZN => n20);
   U21 : OAI21_X1 port map( B1 => net108790, B2 => n69, A => n19, ZN => n174);
   U22 : NAND2_X1 port map( A1 => din(45), A2 => n16, ZN => n19);
   U23 : OAI21_X1 port map( B1 => net108791, B2 => n68, A => n18, ZN => n175);
   U24 : NAND2_X1 port map( A1 => din(46), A2 => n16, ZN => n18);
   U25 : OAI21_X1 port map( B1 => net108792, B2 => n70, A => n17, ZN => n176);
   U26 : NAND2_X1 port map( A1 => din(47), A2 => n16, ZN => n17);
   U27 : OAI21_X1 port map( B1 => net108785, B2 => n69, A => n24, ZN => n169);
   U28 : NAND2_X1 port map( A1 => din(40), A2 => n16, ZN => n24);
   U29 : OAI21_X1 port map( B1 => net108786, B2 => n68, A => n23, ZN => n170);
   U30 : NAND2_X1 port map( A1 => din(41), A2 => n16, ZN => n23);
   U31 : OAI21_X1 port map( B1 => net108787, B2 => n68, A => n22, ZN => n171);
   U32 : NAND2_X1 port map( A1 => din(42), A2 => n16, ZN => n22);
   U33 : OAI21_X1 port map( B1 => net108788, B2 => n68, A => n21, ZN => n172);
   U34 : NAND2_X1 port map( A1 => din(43), A2 => n16, ZN => n21);
   U35 : OAI21_X1 port map( B1 => net108781, B2 => n68, A => n28, ZN => n165);
   U36 : NAND2_X1 port map( A1 => din(36), A2 => n16, ZN => n28);
   U37 : OAI21_X1 port map( B1 => net108782, B2 => n69, A => n27, ZN => n166);
   U38 : NAND2_X1 port map( A1 => din(37), A2 => n65, ZN => n27);
   U39 : OAI21_X1 port map( B1 => net108783, B2 => n68, A => n26, ZN => n167);
   U40 : NAND2_X1 port map( A1 => din(38), A2 => n65, ZN => n26);
   U41 : OAI21_X1 port map( B1 => net108784, B2 => n68, A => n25, ZN => n168);
   U42 : NAND2_X1 port map( A1 => din(39), A2 => n16, ZN => n25);
   U43 : OAI21_X1 port map( B1 => net108769, B2 => n69, A => n40, ZN => n153);
   U44 : NAND2_X1 port map( A1 => din(24), A2 => n67, ZN => n40);
   U45 : OAI21_X1 port map( B1 => net108770, B2 => n69, A => n39, ZN => n154);
   U46 : NAND2_X1 port map( A1 => din(25), A2 => n67, ZN => n39);
   U47 : OAI21_X1 port map( B1 => net108771, B2 => n69, A => n38, ZN => n155);
   U48 : NAND2_X1 port map( A1 => din(26), A2 => n66, ZN => n38);
   U49 : OAI21_X1 port map( B1 => net108772, B2 => n69, A => n37, ZN => n156);
   U50 : NAND2_X1 port map( A1 => din(27), A2 => n67, ZN => n37);
   U51 : OAI21_X1 port map( B1 => net108773, B2 => n69, A => n36, ZN => n157);
   U52 : NAND2_X1 port map( A1 => din(28), A2 => n67, ZN => n36);
   U53 : OAI21_X1 port map( B1 => net108774, B2 => n69, A => n35, ZN => n158);
   U54 : NAND2_X1 port map( A1 => din(29), A2 => n67, ZN => n35);
   U55 : OAI21_X1 port map( B1 => net108775, B2 => n69, A => n34, ZN => n159);
   U56 : NAND2_X1 port map( A1 => din(30), A2 => n66, ZN => n34);
   U57 : OAI21_X1 port map( B1 => net108776, B2 => n68, A => n33, ZN => n160);
   U58 : NAND2_X1 port map( A1 => din(31), A2 => n67, ZN => n33);
   U59 : OAI21_X1 port map( B1 => net108752, B2 => n71, A => n57, ZN => n136);
   U60 : NAND2_X1 port map( A1 => din(7), A2 => n65, ZN => n57);
   U61 : OAI21_X1 port map( B1 => net108756, B2 => n71, A => n53, ZN => n140);
   U62 : NAND2_X1 port map( A1 => din(11), A2 => n65, ZN => n53);
   U63 : OAI21_X1 port map( B1 => net108757, B2 => n70, A => n52, ZN => n141);
   U64 : NAND2_X1 port map( A1 => din(12), A2 => n66, ZN => n52);
   U65 : OAI21_X1 port map( B1 => net108758, B2 => n70, A => n51, ZN => n142);
   U66 : NAND2_X1 port map( A1 => din(13), A2 => n65, ZN => n51);
   U67 : OAI21_X1 port map( B1 => net108759, B2 => n70, A => n50, ZN => n143);
   U68 : NAND2_X1 port map( A1 => din(14), A2 => n66, ZN => n50);
   U69 : OAI21_X1 port map( B1 => net108760, B2 => n70, A => n49, ZN => n144);
   U70 : NAND2_X1 port map( A1 => din(15), A2 => n66, ZN => n49);
   U71 : OAI21_X1 port map( B1 => net108761, B2 => n70, A => n48, ZN => n145);
   U72 : NAND2_X1 port map( A1 => din(16), A2 => n66, ZN => n48);
   U73 : OAI21_X1 port map( B1 => net108762, B2 => n70, A => n47, ZN => n146);
   U74 : NAND2_X1 port map( A1 => din(17), A2 => n67, ZN => n47);
   U75 : OAI21_X1 port map( B1 => net108763, B2 => n70, A => n46, ZN => n147);
   U76 : NAND2_X1 port map( A1 => din(18), A2 => n67, ZN => n46);
   U77 : OAI21_X1 port map( B1 => net108764, B2 => n69, A => n45, ZN => n148);
   U78 : NAND2_X1 port map( A1 => din(19), A2 => n67, ZN => n45);
   U79 : OAI21_X1 port map( B1 => net108765, B2 => n70, A => n44, ZN => n149);
   U80 : NAND2_X1 port map( A1 => din(20), A2 => n67, ZN => n44);
   U81 : OAI21_X1 port map( B1 => net108766, B2 => n70, A => n43, ZN => n150);
   U82 : NAND2_X1 port map( A1 => din(21), A2 => n66, ZN => n43);
   U83 : OAI21_X1 port map( B1 => net108767, B2 => n70, A => n42, ZN => n151);
   U84 : NAND2_X1 port map( A1 => din(22), A2 => n67, ZN => n42);
   U85 : OAI21_X1 port map( B1 => net108768, B2 => n70, A => n41, ZN => n152);
   U86 : NAND2_X1 port map( A1 => din(23), A2 => n67, ZN => n41);
   U87 : OAI21_X1 port map( B1 => net108745, B2 => n71, A => n64, ZN => n129);
   U88 : NAND2_X1 port map( A1 => din(0), A2 => n16, ZN => n64);
   U89 : OAI21_X1 port map( B1 => net108750, B2 => n71, A => n59, ZN => n134);
   U90 : NAND2_X1 port map( A1 => din(5), A2 => n65, ZN => n59);
   U91 : OAI21_X1 port map( B1 => net108746, B2 => n71, A => n63, ZN => n130);
   U92 : NAND2_X1 port map( A1 => din(1), A2 => n16, ZN => n63);
   U93 : OAI21_X1 port map( B1 => net108747, B2 => n71, A => n62, ZN => n131);
   U94 : NAND2_X1 port map( A1 => din(2), A2 => n65, ZN => n62);
   U95 : OAI21_X1 port map( B1 => net108748, B2 => n71, A => n61, ZN => n132);
   U96 : NAND2_X1 port map( A1 => din(3), A2 => n65, ZN => n61);
   U97 : OAI21_X1 port map( B1 => net108749, B2 => n71, A => n60, ZN => n133);
   U98 : NAND2_X1 port map( A1 => din(4), A2 => n65, ZN => n60);
   U99 : OAI21_X1 port map( B1 => net108751, B2 => n71, A => n58, ZN => n135);
   U100 : NAND2_X1 port map( A1 => din(6), A2 => n65, ZN => n58);
   U101 : OAI21_X1 port map( B1 => net108753, B2 => n71, A => n56, ZN => n137);
   U102 : NAND2_X1 port map( A1 => din(8), A2 => n65, ZN => n56);
   U103 : OAI21_X1 port map( B1 => net108754, B2 => n71, A => n55, ZN => n138);
   U104 : NAND2_X1 port map( A1 => din(9), A2 => n66, ZN => n55);
   U105 : OAI21_X1 port map( B1 => net108755, B2 => n71, A => n54, ZN => n139);
   U106 : NAND2_X1 port map( A1 => din(10), A2 => n66, ZN => n54);
   U107 : CLKBUF_X1 port map( A => rst, Z => n7);
   U108 : CLKBUF_X1 port map( A => rst, Z => n8);
   U109 : CLKBUF_X1 port map( A => rst, Z => n9);
   U110 : CLKBUF_X1 port map( A => rst, Z => n10);
   U111 : CLKBUF_X1 port map( A => rst, Z => n11);
   U112 : CLKBUF_X1 port map( A => rst, Z => n12);
   U113 : CLKBUF_X1 port map( A => en, Z => n13);
   U114 : CLKBUF_X1 port map( A => en, Z => n14);
   U115 : CLKBUF_X1 port map( A => en, Z => n15);
   U116 : MUX2_X1 port map( A => dout_48_port, B => din(48), S => n72, Z => 
                           n177);
   U117 : MUX2_X1 port map( A => dout_49_port, B => din(49), S => n72, Z => 
                           n178);
   U118 : MUX2_X1 port map( A => dout_50_port, B => din(50), S => n72, Z => 
                           n179);
   U119 : MUX2_X1 port map( A => dout_51_port, B => din(51), S => n72, Z => 
                           n180);
   U120 : MUX2_X1 port map( A => dout_52_port, B => din(52), S => n72, Z => 
                           n181);
   U121 : MUX2_X1 port map( A => dout_53_port, B => din(53), S => n72, Z => 
                           n182);
   U122 : MUX2_X1 port map( A => dout_54_port, B => din(54), S => n72, Z => 
                           n183);
   U123 : MUX2_X1 port map( A => dout_55_port, B => din(55), S => n72, Z => 
                           n184);
   U124 : MUX2_X1 port map( A => dout_56_port, B => din(56), S => n72, Z => 
                           n185);
   U125 : MUX2_X1 port map( A => dout_57_port, B => din(57), S => n72, Z => 
                           n186);
   U126 : MUX2_X1 port map( A => dout_58_port, B => din(58), S => n72, Z => 
                           n187);
   U127 : MUX2_X1 port map( A => dout_59_port, B => din(59), S => n72, Z => 
                           n188);
   U128 : MUX2_X1 port map( A => dout_60_port, B => din(60), S => n72, Z => 
                           n189);
   U129 : MUX2_X1 port map( A => dout_61_port, B => din(61), S => n72, Z => 
                           n190);
   U130 : MUX2_X1 port map( A => dout_62_port, B => din(62), S => n72, Z => 
                           n191);
   U131 : MUX2_X1 port map( A => dout_63_port, B => din(63), S => n72, Z => 
                           n192);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AddSub_DATA_SIZE64 is

   port( as : in std_logic;  a, b : in std_logic_vector (63 downto 0);  re : 
         out std_logic_vector (63 downto 0);  cout : out std_logic);

end AddSub_DATA_SIZE64;

architecture SYN_add_sub_arch of AddSub_DATA_SIZE64 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component Adder_DATA_SIZE64
      port( cin : in std_logic;  a, b : in std_logic_vector (63 downto 0);  s :
            out std_logic_vector (63 downto 0);  cout : out std_logic);
   end component;
   
   signal b_new_63_port, b_new_62_port, b_new_61_port, b_new_60_port, 
      b_new_59_port, b_new_58_port, b_new_57_port, b_new_56_port, b_new_55_port
      , b_new_54_port, b_new_53_port, b_new_52_port, b_new_51_port, 
      b_new_50_port, b_new_49_port, b_new_48_port, b_new_47_port, b_new_46_port
      , b_new_45_port, b_new_44_port, b_new_43_port, b_new_42_port, 
      b_new_41_port, b_new_40_port, b_new_39_port, b_new_38_port, b_new_37_port
      , b_new_36_port, b_new_35_port, b_new_34_port, b_new_33_port, 
      b_new_32_port, b_new_31_port, b_new_30_port, b_new_29_port, b_new_28_port
      , b_new_27_port, b_new_26_port, b_new_25_port, b_new_24_port, 
      b_new_23_port, b_new_22_port, b_new_21_port, b_new_20_port, b_new_19_port
      , b_new_18_port, b_new_17_port, b_new_16_port, b_new_15_port, 
      b_new_14_port, b_new_13_port, b_new_12_port, b_new_11_port, b_new_10_port
      , b_new_9_port, b_new_8_port, b_new_7_port, b_new_6_port, b_new_5_port, 
      b_new_4_port, b_new_3_port, b_new_2_port, b_new_1_port, b_new_0_port, n1,
      n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17 : 
      std_logic;

begin
   
   U5 : XOR2_X1 port map( A => b(63), B => n9, Z => b_new_63_port);
   U6 : XOR2_X1 port map( A => b(62), B => n8, Z => b_new_62_port);
   U7 : XOR2_X1 port map( A => b(61), B => n8, Z => b_new_61_port);
   U8 : XOR2_X1 port map( A => b(60), B => n9, Z => b_new_60_port);
   U10 : XOR2_X1 port map( A => b(59), B => n8, Z => b_new_59_port);
   U11 : XOR2_X1 port map( A => b(58), B => n9, Z => b_new_58_port);
   U12 : XOR2_X1 port map( A => b(57), B => n9, Z => b_new_57_port);
   U13 : XOR2_X1 port map( A => b(56), B => n8, Z => b_new_56_port);
   U14 : XOR2_X1 port map( A => b(55), B => n9, Z => b_new_55_port);
   U15 : XOR2_X1 port map( A => b(54), B => n8, Z => b_new_54_port);
   U16 : XOR2_X1 port map( A => b(53), B => n9, Z => b_new_53_port);
   U17 : XOR2_X1 port map( A => b(52), B => n8, Z => b_new_52_port);
   U18 : XOR2_X1 port map( A => b(51), B => n9, Z => b_new_51_port);
   U19 : XOR2_X1 port map( A => b(50), B => n8, Z => b_new_50_port);
   U21 : XOR2_X1 port map( A => b(49), B => n9, Z => b_new_49_port);
   U22 : XOR2_X1 port map( A => b(48), B => n9, Z => b_new_48_port);
   U23 : XOR2_X1 port map( A => b(47), B => n8, Z => b_new_47_port);
   U24 : XOR2_X1 port map( A => b(46), B => n9, Z => b_new_46_port);
   U25 : XOR2_X1 port map( A => b(45), B => n8, Z => b_new_45_port);
   U26 : XOR2_X1 port map( A => b(44), B => n9, Z => b_new_44_port);
   U27 : XOR2_X1 port map( A => b(43), B => n8, Z => b_new_43_port);
   U28 : XOR2_X1 port map( A => b(42), B => n8, Z => b_new_42_port);
   U29 : XOR2_X1 port map( A => b(41), B => n8, Z => b_new_41_port);
   U30 : XOR2_X1 port map( A => b(40), B => n9, Z => b_new_40_port);
   U32 : XOR2_X1 port map( A => b(39), B => n8, Z => b_new_39_port);
   U33 : XOR2_X1 port map( A => b(38), B => n9, Z => b_new_38_port);
   U34 : XOR2_X1 port map( A => b(37), B => n9, Z => b_new_37_port);
   U35 : XOR2_X1 port map( A => b(36), B => n8, Z => b_new_36_port);
   U36 : XOR2_X1 port map( A => b(35), B => n9, Z => b_new_35_port);
   U37 : XOR2_X1 port map( A => b(34), B => n9, Z => b_new_34_port);
   U38 : XOR2_X1 port map( A => b(33), B => n9, Z => b_new_33_port);
   U39 : XOR2_X1 port map( A => b(32), B => n9, Z => b_new_32_port);
   U40 : XOR2_X1 port map( A => b(31), B => n9, Z => b_new_31_port);
   U41 : XOR2_X1 port map( A => b(30), B => n8, Z => b_new_30_port);
   U43 : XOR2_X1 port map( A => b(29), B => n9, Z => b_new_29_port);
   U44 : XOR2_X1 port map( A => b(28), B => n8, Z => b_new_28_port);
   U45 : XOR2_X1 port map( A => b(27), B => n8, Z => b_new_27_port);
   U46 : XOR2_X1 port map( A => b(26), B => n8, Z => b_new_26_port);
   U47 : XOR2_X1 port map( A => b(25), B => n9, Z => b_new_25_port);
   U48 : XOR2_X1 port map( A => b(24), B => n8, Z => b_new_24_port);
   U49 : XOR2_X1 port map( A => b(23), B => n8, Z => b_new_23_port);
   U50 : XOR2_X1 port map( A => b(22), B => n8, Z => b_new_22_port);
   U51 : XOR2_X1 port map( A => b(21), B => n9, Z => b_new_21_port);
   U52 : XOR2_X1 port map( A => b(20), B => n8, Z => b_new_20_port);
   U54 : XOR2_X1 port map( A => b(19), B => n9, Z => b_new_19_port);
   U55 : XOR2_X1 port map( A => b(18), B => n8, Z => b_new_18_port);
   U56 : XOR2_X1 port map( A => b(17), B => n9, Z => b_new_17_port);
   U57 : XOR2_X1 port map( A => b(16), B => n9, Z => b_new_16_port);
   U58 : XOR2_X1 port map( A => b(15), B => n8, Z => b_new_15_port);
   U59 : XOR2_X1 port map( A => b(14), B => n8, Z => b_new_14_port);
   U60 : XOR2_X1 port map( A => b(13), B => n8, Z => b_new_13_port);
   U61 : XOR2_X1 port map( A => b(12), B => n9, Z => b_new_12_port);
   ADDER0 : Adder_DATA_SIZE64 port map( cin => n5, a(63) => a(63), a(62) => 
                           a(62), a(61) => a(61), a(60) => a(60), a(59) => 
                           a(59), a(58) => a(58), a(57) => a(57), a(56) => 
                           a(56), a(55) => a(55), a(54) => a(54), a(53) => 
                           a(53), a(52) => a(52), a(51) => a(51), a(50) => 
                           a(50), a(49) => a(49), a(48) => a(48), a(47) => 
                           a(47), a(46) => a(46), a(45) => a(45), a(44) => 
                           a(44), a(43) => a(43), a(42) => a(42), a(41) => 
                           a(41), a(40) => a(40), a(39) => a(39), a(38) => 
                           a(38), a(37) => a(37), a(36) => a(36), a(35) => 
                           a(35), a(34) => a(34), a(33) => a(33), a(32) => 
                           a(32), a(31) => a(31), a(30) => a(30), a(29) => 
                           a(29), a(28) => a(28), a(27) => a(27), a(26) => 
                           a(26), a(25) => a(25), a(24) => a(24), a(23) => 
                           a(23), a(22) => a(22), a(21) => a(21), a(20) => 
                           a(20), a(19) => a(19), a(18) => a(18), a(17) => 
                           a(17), a(16) => a(16), a(15) => a(15), a(14) => 
                           a(14), a(13) => a(13), a(12) => a(12), a(11) => 
                           a(11), a(10) => a(10), a(9) => a(9), a(8) => a(8), 
                           a(7) => a(7), a(6) => a(6), a(5) => a(5), a(4) => 
                           a(4), a(3) => a(3), a(2) => a(2), a(1) => a(1), a(0)
                           => a(0), b(63) => b_new_63_port, b(62) => 
                           b_new_62_port, b(61) => b_new_61_port, b(60) => 
                           b_new_60_port, b(59) => b_new_59_port, b(58) => 
                           b_new_58_port, b(57) => b_new_57_port, b(56) => 
                           b_new_56_port, b(55) => b_new_55_port, b(54) => 
                           b_new_54_port, b(53) => b_new_53_port, b(52) => 
                           b_new_52_port, b(51) => b_new_51_port, b(50) => 
                           b_new_50_port, b(49) => b_new_49_port, b(48) => 
                           b_new_48_port, b(47) => b_new_47_port, b(46) => 
                           b_new_46_port, b(45) => b_new_45_port, b(44) => 
                           b_new_44_port, b(43) => b_new_43_port, b(42) => 
                           b_new_42_port, b(41) => b_new_41_port, b(40) => 
                           b_new_40_port, b(39) => b_new_39_port, b(38) => 
                           b_new_38_port, b(37) => b_new_37_port, b(36) => 
                           b_new_36_port, b(35) => b_new_35_port, b(34) => 
                           b_new_34_port, b(33) => b_new_33_port, b(32) => 
                           b_new_32_port, b(31) => b_new_31_port, b(30) => 
                           b_new_30_port, b(29) => b_new_29_port, b(28) => 
                           b_new_28_port, b(27) => b_new_27_port, b(26) => 
                           b_new_26_port, b(25) => b_new_25_port, b(24) => 
                           b_new_24_port, b(23) => b_new_23_port, b(22) => 
                           b_new_22_port, b(21) => b_new_21_port, b(20) => 
                           b_new_20_port, b(19) => b_new_19_port, b(18) => 
                           b_new_18_port, b(17) => b_new_17_port, b(16) => 
                           b_new_16_port, b(15) => b_new_15_port, b(14) => 
                           b_new_14_port, b(13) => b_new_13_port, b(12) => 
                           b_new_12_port, b(11) => b_new_11_port, b(10) => 
                           b_new_10_port, b(9) => b_new_9_port, b(8) => 
                           b_new_8_port, b(7) => b_new_7_port, b(6) => 
                           b_new_6_port, b(5) => b_new_5_port, b(4) => 
                           b_new_4_port, b(3) => b_new_3_port, b(2) => 
                           b_new_2_port, b(1) => b_new_1_port, b(0) => 
                           b_new_0_port, s(63) => re(63), s(62) => re(62), 
                           s(61) => re(61), s(60) => re(60), s(59) => re(59), 
                           s(58) => re(58), s(57) => re(57), s(56) => re(56), 
                           s(55) => re(55), s(54) => re(54), s(53) => re(53), 
                           s(52) => re(52), s(51) => re(51), s(50) => re(50), 
                           s(49) => re(49), s(48) => re(48), s(47) => re(47), 
                           s(46) => re(46), s(45) => re(45), s(44) => re(44), 
                           s(43) => re(43), s(42) => re(42), s(41) => re(41), 
                           s(40) => re(40), s(39) => re(39), s(38) => re(38), 
                           s(37) => re(37), s(36) => re(36), s(35) => re(35), 
                           s(34) => re(34), s(33) => re(33), s(32) => re(32), 
                           s(31) => re(31), s(30) => re(30), s(29) => re(29), 
                           s(28) => re(28), s(27) => re(27), s(26) => re(26), 
                           s(25) => re(25), s(24) => re(24), s(23) => re(23), 
                           s(22) => re(22), s(21) => re(21), s(20) => re(20), 
                           s(19) => re(19), s(18) => re(18), s(17) => re(17), 
                           s(16) => re(16), s(15) => re(15), s(14) => re(14), 
                           s(13) => re(13), s(12) => re(12), s(11) => re(11), 
                           s(10) => re(10), s(9) => re(9), s(8) => re(8), s(7) 
                           => re(7), s(6) => re(6), s(5) => re(5), s(4) => 
                           re(4), s(3) => re(3), s(2) => re(2), s(1) => re(1), 
                           s(0) => re(0), cout => cout);
   U1 : INV_X1 port map( A => b(2), ZN => n1);
   U2 : BUF_X1 port map( A => n15, Z => n7);
   U3 : BUF_X1 port map( A => as, Z => n6);
   U4 : XNOR2_X1 port map( A => n7, B => n1, ZN => b_new_2_port);
   U9 : BUF_X1 port map( A => as, Z => n14);
   U20 : BUF_X1 port map( A => n6, Z => n5);
   U31 : BUF_X1 port map( A => as, Z => n15);
   U42 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => b_new_1_port);
   U53 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => b_new_0_port);
   U62 : NAND2_X1 port map( A1 => n6, A2 => n17, ZN => n3);
   U63 : NAND2_X1 port map( A1 => n2, A2 => b(1), ZN => n4);
   U64 : INV_X1 port map( A => n15, ZN => n2);
   U65 : BUF_X4 port map( A => n14, Z => n8);
   U66 : BUF_X4 port map( A => n15, Z => n9);
   U67 : NAND2_X1 port map( A1 => n6, A2 => n11, ZN => n12);
   U68 : NAND2_X1 port map( A1 => n10, A2 => b(0), ZN => n13);
   U69 : INV_X1 port map( A => n14, ZN => n10);
   U70 : INV_X1 port map( A => b(0), ZN => n11);
   U71 : XOR2_X1 port map( A => n7, B => b(4), Z => b_new_4_port);
   U72 : XOR2_X1 port map( A => n8, B => b(10), Z => b_new_10_port);
   U73 : XOR2_X1 port map( A => n8, B => b(6), Z => b_new_6_port);
   U74 : XOR2_X1 port map( A => n8, B => b(8), Z => b_new_8_port);
   U75 : XOR2_X1 port map( A => n9, B => b(9), Z => b_new_9_port);
   U76 : XOR2_X1 port map( A => n9, B => b(11), Z => b_new_11_port);
   U77 : XOR2_X1 port map( A => n9, B => b(7), Z => b_new_7_port);
   U78 : XOR2_X1 port map( A => n7, B => b(3), Z => b_new_3_port);
   U79 : INV_X1 port map( A => b(5), ZN => n16);
   U80 : XNOR2_X1 port map( A => n9, B => n16, ZN => b_new_5_port);
   U81 : INV_X1 port map( A => b(1), ZN => n17);

end SYN_add_sub_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE64 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (63 downto 0);  
         dout : out std_logic_vector (63 downto 0));

end Mux_DATA_SIZE64;

architecture SYN_mux_arch of Mux_DATA_SIZE64 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : MUX2_X1 port map( A => din0(0), B => din1(0), S => n3, Z => dout(0));
   U2 : CLKBUF_X1 port map( A => n4, Z => n5);
   U3 : CLKBUF_X1 port map( A => sel, Z => n4);
   U4 : BUF_X1 port map( A => n3, Z => n2);
   U5 : BUF_X1 port map( A => n3, Z => n1);
   U6 : CLKBUF_X1 port map( A => sel, Z => n3);
   U7 : CLKBUF_X1 port map( A => n4, Z => n6);
   U8 : CLKBUF_X1 port map( A => n4, Z => n7);
   U9 : MUX2_X1 port map( A => din0(1), B => din1(1), S => n1, Z => dout(1));
   U10 : MUX2_X1 port map( A => din0(2), B => din1(2), S => n2, Z => dout(2));
   U11 : MUX2_X1 port map( A => din0(3), B => din1(3), S => n1, Z => dout(3));
   U12 : MUX2_X1 port map( A => din0(4), B => din1(4), S => n2, Z => dout(4));
   U13 : MUX2_X1 port map( A => din0(5), B => din1(5), S => n1, Z => dout(5));
   U14 : MUX2_X1 port map( A => din0(6), B => din1(6), S => n2, Z => dout(6));
   U15 : MUX2_X1 port map( A => din0(7), B => din1(7), S => n1, Z => dout(7));
   U16 : MUX2_X1 port map( A => din0(8), B => din1(8), S => n2, Z => dout(8));
   U17 : MUX2_X1 port map( A => din0(9), B => din1(9), S => n1, Z => dout(9));
   U18 : MUX2_X1 port map( A => din0(10), B => din1(10), S => n2, Z => dout(10)
                           );
   U19 : MUX2_X1 port map( A => din0(11), B => din1(11), S => n1, Z => dout(11)
                           );
   U20 : MUX2_X1 port map( A => din0(12), B => din1(12), S => n4, Z => dout(12)
                           );
   U21 : MUX2_X1 port map( A => din0(13), B => din1(13), S => n4, Z => dout(13)
                           );
   U22 : MUX2_X1 port map( A => din0(14), B => din1(14), S => n4, Z => dout(14)
                           );
   U23 : MUX2_X1 port map( A => din0(15), B => din1(15), S => n4, Z => dout(15)
                           );
   U24 : MUX2_X1 port map( A => din0(16), B => din1(16), S => n4, Z => dout(16)
                           );
   U25 : MUX2_X1 port map( A => din0(17), B => din1(17), S => n4, Z => dout(17)
                           );
   U26 : MUX2_X1 port map( A => din0(18), B => din1(18), S => n4, Z => dout(18)
                           );
   U27 : MUX2_X1 port map( A => din0(19), B => din1(19), S => n4, Z => dout(19)
                           );
   U28 : MUX2_X1 port map( A => din0(20), B => din1(20), S => n4, Z => dout(20)
                           );
   U29 : MUX2_X1 port map( A => din0(21), B => din1(21), S => n4, Z => dout(21)
                           );
   U30 : MUX2_X1 port map( A => din0(22), B => din1(22), S => n4, Z => dout(22)
                           );
   U31 : MUX2_X1 port map( A => din0(23), B => din1(23), S => n4, Z => dout(23)
                           );
   U32 : MUX2_X1 port map( A => din0(24), B => din1(24), S => n5, Z => dout(24)
                           );
   U33 : MUX2_X1 port map( A => din0(25), B => din1(25), S => n5, Z => dout(25)
                           );
   U34 : MUX2_X1 port map( A => din0(26), B => din1(26), S => n5, Z => dout(26)
                           );
   U35 : MUX2_X1 port map( A => din0(27), B => din1(27), S => n5, Z => dout(27)
                           );
   U36 : MUX2_X1 port map( A => din0(28), B => din1(28), S => n5, Z => dout(28)
                           );
   U37 : MUX2_X1 port map( A => din0(29), B => din1(29), S => n5, Z => dout(29)
                           );
   U38 : MUX2_X1 port map( A => din0(30), B => din1(30), S => n5, Z => dout(30)
                           );
   U39 : MUX2_X1 port map( A => din0(31), B => din1(31), S => n5, Z => dout(31)
                           );
   U40 : MUX2_X1 port map( A => din0(32), B => din1(32), S => n5, Z => dout(32)
                           );
   U41 : MUX2_X1 port map( A => din0(33), B => din1(33), S => n5, Z => dout(33)
                           );
   U42 : MUX2_X1 port map( A => din0(34), B => din1(34), S => n5, Z => dout(34)
                           );
   U43 : MUX2_X1 port map( A => din0(35), B => din1(35), S => n5, Z => dout(35)
                           );
   U44 : MUX2_X1 port map( A => din0(36), B => din1(36), S => n6, Z => dout(36)
                           );
   U45 : MUX2_X1 port map( A => din0(37), B => din1(37), S => n6, Z => dout(37)
                           );
   U46 : MUX2_X1 port map( A => din0(38), B => din1(38), S => n6, Z => dout(38)
                           );
   U47 : MUX2_X1 port map( A => din0(39), B => din1(39), S => n6, Z => dout(39)
                           );
   U48 : MUX2_X1 port map( A => din0(40), B => din1(40), S => n6, Z => dout(40)
                           );
   U49 : MUX2_X1 port map( A => din0(41), B => din1(41), S => n6, Z => dout(41)
                           );
   U50 : MUX2_X1 port map( A => din0(42), B => din1(42), S => n6, Z => dout(42)
                           );
   U51 : MUX2_X1 port map( A => din0(43), B => din1(43), S => n6, Z => dout(43)
                           );
   U52 : MUX2_X1 port map( A => din0(44), B => din1(44), S => n6, Z => dout(44)
                           );
   U53 : MUX2_X1 port map( A => din0(45), B => din1(45), S => n6, Z => dout(45)
                           );
   U54 : MUX2_X1 port map( A => din0(46), B => din1(46), S => n6, Z => dout(46)
                           );
   U55 : MUX2_X1 port map( A => din0(47), B => din1(47), S => n6, Z => dout(47)
                           );
   U56 : MUX2_X1 port map( A => din0(48), B => din1(48), S => n7, Z => dout(48)
                           );
   U57 : MUX2_X1 port map( A => din0(49), B => din1(49), S => n7, Z => dout(49)
                           );
   U58 : MUX2_X1 port map( A => din0(50), B => din1(50), S => n7, Z => dout(50)
                           );
   U59 : MUX2_X1 port map( A => din0(51), B => din1(51), S => n7, Z => dout(51)
                           );
   U60 : MUX2_X1 port map( A => din0(52), B => din1(52), S => n7, Z => dout(52)
                           );
   U61 : MUX2_X1 port map( A => din0(53), B => din1(53), S => n7, Z => dout(53)
                           );
   U62 : MUX2_X1 port map( A => din0(54), B => din1(54), S => n7, Z => dout(54)
                           );
   U63 : MUX2_X1 port map( A => din0(55), B => din1(55), S => n7, Z => dout(55)
                           );
   U64 : MUX2_X1 port map( A => din0(56), B => din1(56), S => n7, Z => dout(56)
                           );
   U65 : MUX2_X1 port map( A => din0(57), B => din1(57), S => n7, Z => dout(57)
                           );
   U66 : MUX2_X1 port map( A => din0(58), B => din1(58), S => n7, Z => dout(58)
                           );
   U67 : MUX2_X1 port map( A => din0(59), B => din1(59), S => n7, Z => dout(59)
                           );
   U68 : MUX2_X1 port map( A => din0(60), B => din1(60), S => n7, Z => dout(60)
                           );
   U69 : MUX2_X1 port map( A => din0(61), B => din1(61), S => n7, Z => dout(61)
                           );
   U70 : MUX2_X1 port map( A => din0(62), B => din1(62), S => n7, Z => dout(62)
                           );
   U71 : MUX2_X1 port map( A => din0(63), B => din1(63), S => sel, Z => 
                           dout(63));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AddSub_DATA_SIZE32_0 is

   port( as : in std_logic;  a, b : in std_logic_vector (31 downto 0);  re : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end AddSub_DATA_SIZE32_0;

architecture SYN_add_sub_arch of AddSub_DATA_SIZE32_0 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component Adder_DATA_SIZE32_4
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal b_new_31_port, b_new_30_port, b_new_29_port, b_new_28_port, 
      b_new_27_port, b_new_26_port, b_new_25_port, b_new_24_port, b_new_23_port
      , b_new_22_port, b_new_21_port, b_new_20_port, b_new_19_port, 
      b_new_18_port, b_new_17_port, b_new_16_port, b_new_15_port, b_new_14_port
      , b_new_13_port, b_new_12_port, b_new_11_port, b_new_10_port, 
      b_new_9_port, b_new_8_port, b_new_7_port, b_new_6_port, b_new_5_port, 
      b_new_4_port, b_new_3_port, b_new_2_port, b_new_1_port, b_new_0_port, n1,
      n2, n3, n4, n5 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b(9), B => n3, Z => b_new_9_port);
   U2 : XOR2_X1 port map( A => b(8), B => n2, Z => b_new_8_port);
   U3 : XOR2_X1 port map( A => b(7), B => n5, Z => b_new_7_port);
   U4 : XOR2_X1 port map( A => b(6), B => n5, Z => b_new_6_port);
   U5 : XOR2_X1 port map( A => b(5), B => n5, Z => b_new_5_port);
   U6 : XOR2_X1 port map( A => b(4), B => n2, Z => b_new_4_port);
   U7 : XOR2_X1 port map( A => b(3), B => n3, Z => b_new_3_port);
   U8 : XOR2_X1 port map( A => b(31), B => n2, Z => b_new_31_port);
   U9 : XOR2_X1 port map( A => b(30), B => n2, Z => b_new_30_port);
   U10 : XOR2_X1 port map( A => b(2), B => n5, Z => b_new_2_port);
   U11 : XOR2_X1 port map( A => b(29), B => n5, Z => b_new_29_port);
   U12 : XOR2_X1 port map( A => b(28), B => n5, Z => b_new_28_port);
   U13 : XOR2_X1 port map( A => b(27), B => n2, Z => b_new_27_port);
   U14 : XOR2_X1 port map( A => b(26), B => n3, Z => b_new_26_port);
   U15 : XOR2_X1 port map( A => b(25), B => n3, Z => b_new_25_port);
   U16 : XOR2_X1 port map( A => b(24), B => n2, Z => b_new_24_port);
   U17 : XOR2_X1 port map( A => b(23), B => n3, Z => b_new_23_port);
   U18 : XOR2_X1 port map( A => b(22), B => n2, Z => b_new_22_port);
   U19 : XOR2_X1 port map( A => b(21), B => n5, Z => b_new_21_port);
   U20 : XOR2_X1 port map( A => b(20), B => n3, Z => b_new_20_port);
   U21 : XOR2_X1 port map( A => b(1), B => n2, Z => b_new_1_port);
   U22 : XOR2_X1 port map( A => b(19), B => n3, Z => b_new_19_port);
   U23 : XOR2_X1 port map( A => b(18), B => n5, Z => b_new_18_port);
   U24 : XOR2_X1 port map( A => b(17), B => n5, Z => b_new_17_port);
   U25 : XOR2_X1 port map( A => b(16), B => n2, Z => b_new_16_port);
   U26 : XOR2_X1 port map( A => b(15), B => n5, Z => b_new_15_port);
   U27 : XOR2_X1 port map( A => b(14), B => n3, Z => b_new_14_port);
   U28 : XOR2_X1 port map( A => b(13), B => n2, Z => b_new_13_port);
   U29 : XOR2_X1 port map( A => b(12), B => n3, Z => b_new_12_port);
   U30 : XOR2_X1 port map( A => b(11), B => n5, Z => b_new_11_port);
   U31 : XOR2_X1 port map( A => b(10), B => n5, Z => b_new_10_port);
   ADDER0 : Adder_DATA_SIZE32_4 port map( cin => n3, a(31) => a(31), a(30) => 
                           a(30), a(29) => a(29), a(28) => a(28), a(27) => 
                           a(27), a(26) => a(26), a(25) => a(25), a(24) => 
                           a(24), a(23) => a(23), a(22) => a(22), a(21) => 
                           a(21), a(20) => a(20), a(19) => a(19), a(18) => 
                           a(18), a(17) => a(17), a(16) => a(16), a(15) => 
                           a(15), a(14) => a(14), a(13) => a(13), a(12) => 
                           a(12), a(11) => a(11), a(10) => a(10), a(9) => a(9),
                           a(8) => a(8), a(7) => a(7), a(6) => a(6), a(5) => 
                           a(5), a(4) => a(4), a(3) => a(3), a(2) => a(2), a(1)
                           => a(1), a(0) => a(0), b(31) => b_new_31_port, b(30)
                           => b_new_30_port, b(29) => b_new_29_port, b(28) => 
                           b_new_28_port, b(27) => b_new_27_port, b(26) => 
                           b_new_26_port, b(25) => b_new_25_port, b(24) => 
                           b_new_24_port, b(23) => b_new_23_port, b(22) => 
                           b_new_22_port, b(21) => b_new_21_port, b(20) => 
                           b_new_20_port, b(19) => b_new_19_port, b(18) => 
                           b_new_18_port, b(17) => b_new_17_port, b(16) => 
                           b_new_16_port, b(15) => b_new_15_port, b(14) => 
                           b_new_14_port, b(13) => b_new_13_port, b(12) => 
                           b_new_12_port, b(11) => b_new_11_port, b(10) => 
                           b_new_10_port, b(9) => b_new_9_port, b(8) => 
                           b_new_8_port, b(7) => b_new_7_port, b(6) => 
                           b_new_6_port, b(5) => b_new_5_port, b(4) => 
                           b_new_4_port, b(3) => b_new_3_port, b(2) => 
                           b_new_2_port, b(1) => b_new_1_port, b(0) => 
                           b_new_0_port, s(31) => re(31), s(30) => re(30), 
                           s(29) => re(29), s(28) => re(28), s(27) => re(27), 
                           s(26) => re(26), s(25) => re(25), s(24) => re(24), 
                           s(23) => re(23), s(22) => re(22), s(21) => re(21), 
                           s(20) => re(20), s(19) => re(19), s(18) => re(18), 
                           s(17) => re(17), s(16) => re(16), s(15) => re(15), 
                           s(14) => re(14), s(13) => re(13), s(12) => re(12), 
                           s(11) => re(11), s(10) => re(10), s(9) => re(9), 
                           s(8) => re(8), s(7) => re(7), s(6) => re(6), s(5) =>
                           re(5), s(4) => re(4), s(3) => re(3), s(2) => re(2), 
                           s(1) => re(1), s(0) => re(0), cout => cout);
   U32 : BUF_X2 port map( A => as, Z => n3);
   U33 : INV_X1 port map( A => b(0), ZN => n4);
   U34 : CLKBUF_X1 port map( A => as, Z => n1);
   U35 : CLKBUF_X1 port map( A => n1, Z => n5);
   U36 : CLKBUF_X3 port map( A => n1, Z => n2);
   U37 : XNOR2_X1 port map( A => n4, B => as, ZN => b_new_0_port);

end SYN_add_sub_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity BoothMul_DATA_SIZE16_STAGE10 is

   port( rst, clk, en, lock, sign : in std_logic;  a, b : in std_logic_vector 
         (15 downto 0);  o : out std_logic_vector (31 downto 0));

end BoothMul_DATA_SIZE16_STAGE10;

architecture SYN_booth_mul_arch of BoothMul_DATA_SIZE16_STAGE10 is

   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BoothMul_DATA_SIZE16_STAGE10_DW01_inc_0
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component Adder_DATA_SIZE32_5
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;
   
   component Reg_DATA_SIZE32_1
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 
            0);  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component AddSub_DATA_SIZE32_1
      port( as : in std_logic;  a, b : in std_logic_vector (31 downto 0);  re :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;
   
   component Mux_DATA_SIZE32_1
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0)
            ;  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component BoothEncoder
      port( din : in std_logic_vector (2 downto 0);  sel : out std_logic_vector
            (2 downto 0));
   end component;
   
   component Adder_DATA_SIZE16
      port( cin : in std_logic;  a, b : in std_logic_vector (15 downto 0);  s :
            out std_logic_vector (15 downto 0);  cout : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic0_port, e_a_31_port, e_a_30_port, e_a_29_port, e_a_28_port, 
      e_a_27_port, e_a_26_port, e_a_25_port, e_a_24_port, e_a_23_port, 
      e_a_22_port, e_a_21_port, e_a_20_port, e_a_19_port, e_a_18_port, 
      e_a_17_port, e_a_16_port, e_a_15_port, e_a_14_port, e_a_13_port, 
      e_a_12_port, e_a_11_port, e_a_10_port, e_a_9_port, e_a_8_port, e_a_7_port
      , e_a_6_port, e_a_5_port, e_a_4_port, e_a_3_port, e_a_2_port, e_a_1_port,
      e_a_0_port, e_b_16_port, e_b_15_port, e_b_14_port, e_b_13_port, 
      e_b_12_port, e_b_11_port, e_b_10_port, e_b_9_port, e_b_8_port, e_b_7_port
      , e_b_6_port, e_b_5_port, e_b_4_port, e_b_3_port, e_b_2_port, e_b_1_port,
      e_b_0_port, adj_final_mod_31_port, adj_final_mod_30_port, 
      adj_final_mod_29_port, adj_final_mod_28_port, adj_final_mod_27_port, 
      adj_final_mod_26_port, adj_final_mod_25_port, adj_final_mod_24_port, 
      adj_final_mod_23_port, adj_final_mod_22_port, adj_final_mod_21_port, 
      adj_final_mod_20_port, adj_final_mod_19_port, adj_final_mod_18_port, 
      adj_final_mod_17_port, adj_final_mod_16_port, adj_final_mod_15_port, 
      adj_final_mod_14_port, adj_final_mod_13_port, adj_final_mod_12_port, 
      adj_final_mod_11_port, adj_final_mod_10_port, adj_final_mod_9_port, 
      adj_final_mod_8_port, adj_final_mod_7_port, adj_final_mod_6_port, 
      adj_final_mod_5_port, adj_final_mod_4_port, adj_final_mod_3_port, 
      adj_final_mod_2_port, adj_final_mod_1_port, adj_final_mod_0_port, N9, N10
      , N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, 
      N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39
      , N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, 
      N54, N55, N56, N57, adj_sum_15_port, adj_sum_14_port, adj_sum_13_port, 
      adj_sum_12_port, adj_sum_11_port, adj_sum_10_port, adj_sum_9_port, 
      adj_sum_8_port, adj_sum_7_port, adj_sum_6_port, adj_sum_5_port, 
      adj_sum_4_port, adj_sum_3_port, adj_sum_2_port, adj_sum_1_port, 
      adj_sum_0_port, adj_cout, sel_2_port, sel_1_port, sel_0_port, 
      mux_out_31_port, mux_out_30_port, mux_out_29_port, mux_out_28_port, 
      mux_out_27_port, mux_out_26_port, mux_out_25_port, mux_out_24_port, 
      mux_out_23_port, mux_out_22_port, mux_out_21_port, mux_out_20_port, 
      mux_out_19_port, mux_out_18_port, mux_out_17_port, mux_out_16_port, 
      mux_out_15_port, mux_out_14_port, mux_out_13_port, mux_out_12_port, 
      mux_out_11_port, mux_out_10_port, mux_out_9_port, mux_out_8_port, 
      mux_out_7_port, mux_out_6_port, mux_out_5_port, mux_out_4_port, 
      mux_out_3_port, mux_out_2_port, mux_out_1_port, mux_out_0_port, 
      zero_out_31_port, zero_out_30_port, zero_out_29_port, zero_out_28_port, 
      zero_out_27_port, zero_out_26_port, zero_out_25_port, zero_out_24_port, 
      zero_out_23_port, zero_out_22_port, zero_out_21_port, zero_out_20_port, 
      zero_out_19_port, zero_out_18_port, zero_out_17_port, zero_out_16_port, 
      zero_out_15_port, zero_out_14_port, zero_out_13_port, zero_out_12_port, 
      zero_out_11_port, zero_out_10_port, zero_out_9_port, zero_out_8_port, 
      zero_out_7_port, zero_out_6_port, zero_out_5_port, zero_out_4_port, 
      zero_out_3_port, zero_out_2_port, zero_out_1_port, zero_out_0_port, 
      add_out_reg_31_port, add_out_reg_30_port, add_out_reg_29_port, 
      add_out_reg_28_port, add_out_reg_27_port, add_out_reg_26_port, 
      add_out_reg_25_port, add_out_reg_24_port, add_out_reg_23_port, 
      add_out_reg_22_port, add_out_reg_21_port, add_out_reg_20_port, 
      add_out_reg_19_port, add_out_reg_18_port, add_out_reg_17_port, 
      add_out_reg_16_port, add_out_reg_15_port, add_out_reg_14_port, 
      add_out_reg_13_port, add_out_reg_12_port, add_out_reg_11_port, 
      add_out_reg_10_port, add_out_reg_9_port, add_out_reg_8_port, 
      add_out_reg_7_port, add_out_reg_6_port, add_out_reg_5_port, 
      add_out_reg_4_port, add_out_reg_3_port, add_out_reg_2_port, 
      add_out_reg_1_port, add_out_reg_0_port, add_out_31_port, add_out_30_port,
      add_out_29_port, add_out_28_port, add_out_27_port, add_out_26_port, 
      add_out_25_port, add_out_24_port, add_out_23_port, add_out_22_port, 
      add_out_21_port, add_out_20_port, add_out_19_port, add_out_18_port, 
      add_out_17_port, add_out_16_port, add_out_15_port, add_out_14_port, 
      add_out_13_port, add_out_12_port, add_out_11_port, add_out_10_port, 
      add_out_9_port, add_out_8_port, add_out_7_port, add_out_6_port, 
      add_out_5_port, add_out_4_port, add_out_3_port, add_out_2_port, 
      add_out_1_port, add_out_0_port, reg_rst, en_o, n_state_31_port, 
      n_state_30_port, n_state_29_port, n_state_28_port, n_state_27_port, 
      n_state_26_port, n_state_25_port, n_state_24_port, n_state_23_port, 
      n_state_22_port, n_state_21_port, n_state_20_port, n_state_19_port, 
      n_state_18_port, n_state_17_port, n_state_16_port, n_state_15_port, 
      n_state_14_port, n_state_13_port, n_state_12_port, n_state_11_port, 
      n_state_10_port, n_state_9_port, n_state_8_port, n_state_7_port, 
      n_state_6_port, n_state_5_port, n_state_4_port, n_state_3_port, 
      n_state_2_port, n_state_1_port, n_state_0_port, c_state_31_port, 
      c_state_30_port, c_state_29_port, c_state_28_port, c_state_27_port, 
      c_state_26_port, c_state_25_port, c_state_24_port, c_state_23_port, 
      c_state_22_port, c_state_21_port, c_state_20_port, c_state_19_port, 
      c_state_18_port, c_state_17_port, c_state_16_port, c_state_15_port, 
      c_state_14_port, c_state_13_port, c_state_12_port, c_state_11_port, 
      c_state_10_port, c_state_9_port, c_state_8_port, c_state_7_port, 
      c_state_6_port, c_state_5_port, c_state_4_port, c_state_3_port, 
      c_state_2_port, c_state_1_port, c_state_0_port, N70, N71, N72, N73, N74, 
      N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89
      , N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, net4347, 
      net4348, n12_port, n13_port, n22_port, n23_port, n24_port, n31_port, n58,
      n65, n66, n67, n68, n69, n70_port, n71_port, n72_port, n79_port, n80_port
      , n81_port, n82_port, n83_port, n84_port, n85_port, n86_port, n87_port, 
      n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, 
      n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, 
      n53_port, n54_port, n55_port, n56_port, n57_port, n59, n60, net108691, 
      net108692, net108693, net108694, net108695, net108696, net108697, 
      net108698, net108699, net108700, net108701, net108702, net108703, 
      net108704, net108705, net108706, net108707, net108708, net108709, 
      net108710, net108711, net108712, net108713, net108714, net108715, 
      net108716, net108717, net108718, net108719, net108720, net108721, 
      net108722, net108723, net108724, net108725, net108726, net108727, 
      net108728, net108729, net108730, net108731, net108732, net108733, 
      net108734, net108735, net108736, net108737, net108738, net108739, 
      net108740, net108741, net108742, net108743, net108744, n77_port, n78_port
      , n88_port, n89_port, n90_port, n91_port, n92_port, n93_port, n95_port, 
      n96_port, n97_port, n98_port, n99_port, n100_port, n101_port, n102, n103,
      n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, 
      n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, 
      n140, n141, n142, n143, n144, n145, n146, n148, n149, n150, n151, n152, 
      n153, n154, n155, n156, n64, n73_port, n74_port, n75_port, n76_port, 
      n94_port, n147, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, 
      net164133, net164134, net164135, net164136, net164137, net164138 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   c_state_reg_0_inst : DFFR_X1 port map( D => n_state_0_port, CK => clk, RN =>
                           n174, Q => c_state_0_port, QN => n211);
   c_state_reg_10_inst : DFFR_X1 port map( D => n_state_10_port, CK => clk, RN 
                           => n176, Q => c_state_10_port, QN => n12_port);
   c_state_reg_1_inst : DFFR_X1 port map( D => n_state_1_port, CK => clk, RN =>
                           n174, Q => c_state_1_port, QN => n13_port);
   c_state_reg_2_inst : DFFR_X1 port map( D => n_state_2_port, CK => clk, RN =>
                           n174, Q => c_state_2_port, QN => n55_port);
   c_state_reg_3_inst : DFFR_X1 port map( D => n_state_3_port, CK => clk, RN =>
                           n174, Q => c_state_3_port, QN => n54_port);
   c_state_reg_4_inst : DFFR_X1 port map( D => n_state_4_port, CK => clk, RN =>
                           n174, Q => c_state_4_port, QN => n57_port);
   c_state_reg_5_inst : DFFR_X1 port map( D => n_state_5_port, CK => clk, RN =>
                           n174, Q => c_state_5_port, QN => n59);
   c_state_reg_6_inst : DFFR_X1 port map( D => n_state_6_port, CK => clk, RN =>
                           n174, Q => c_state_6_port, QN => net108744);
   c_state_reg_7_inst : DFFR_X1 port map( D => n_state_7_port, CK => clk, RN =>
                           n174, Q => c_state_7_port, QN => net108743);
   c_state_reg_8_inst : DFFR_X1 port map( D => n_state_8_port, CK => clk, RN =>
                           n174, Q => c_state_8_port, QN => net108742);
   c_state_reg_9_inst : DFFR_X1 port map( D => n_state_9_port, CK => clk, RN =>
                           n174, Q => c_state_9_port, QN => n56_port);
   c_state_reg_11_inst : DFFR_X1 port map( D => n_state_11_port, CK => clk, RN 
                           => n176, Q => c_state_11_port, QN => n22_port);
   c_state_reg_12_inst : DFFR_X1 port map( D => n_state_12_port, CK => clk, RN 
                           => n176, Q => c_state_12_port, QN => n23_port);
   c_state_reg_13_inst : DFFR_X1 port map( D => n_state_13_port, CK => clk, RN 
                           => n176, Q => c_state_13_port, QN => n24_port);
   c_state_reg_14_inst : DFFR_X1 port map( D => n_state_14_port, CK => clk, RN 
                           => n176, Q => c_state_14_port, QN => net108741);
   c_state_reg_15_inst : DFFR_X1 port map( D => n_state_15_port, CK => clk, RN 
                           => n176, Q => c_state_15_port, QN => net108740);
   c_state_reg_16_inst : DFFR_X1 port map( D => n_state_16_port, CK => clk, RN 
                           => n176, Q => c_state_16_port, QN => net108739);
   c_state_reg_17_inst : DFFR_X1 port map( D => n_state_17_port, CK => clk, RN 
                           => n176, Q => c_state_17_port, QN => net164138);
   c_state_reg_18_inst : DFFR_X1 port map( D => n_state_18_port, CK => clk, RN 
                           => n175, Q => c_state_18_port, QN => net164137);
   c_state_reg_19_inst : DFFR_X1 port map( D => n_state_19_port, CK => clk, RN 
                           => n175, Q => c_state_19_port, QN => net164136);
   c_state_reg_20_inst : DFFR_X1 port map( D => n_state_20_port, CK => clk, RN 
                           => n175, Q => c_state_20_port, QN => n31_port);
   c_state_reg_21_inst : DFFR_X1 port map( D => n_state_21_port, CK => clk, RN 
                           => n175, Q => c_state_21_port, QN => net108738);
   c_state_reg_22_inst : DFFR_X1 port map( D => n_state_22_port, CK => clk, RN 
                           => n175, Q => c_state_22_port, QN => net108737);
   c_state_reg_23_inst : DFFR_X1 port map( D => n_state_23_port, CK => clk, RN 
                           => n175, Q => c_state_23_port, QN => net108736);
   c_state_reg_24_inst : DFFR_X1 port map( D => n_state_24_port, CK => clk, RN 
                           => n175, Q => c_state_24_port, QN => net164135);
   c_state_reg_25_inst : DFFR_X1 port map( D => n_state_25_port, CK => clk, RN 
                           => n175, Q => c_state_25_port, QN => net164134);
   c_state_reg_26_inst : DFFR_X1 port map( D => n_state_26_port, CK => clk, RN 
                           => n175, Q => c_state_26_port, QN => net108735);
   c_state_reg_27_inst : DFFR_X1 port map( D => n_state_27_port, CK => clk, RN 
                           => n175, Q => c_state_27_port, QN => net108734);
   c_state_reg_28_inst : DFFR_X1 port map( D => n_state_28_port, CK => clk, RN 
                           => n175, Q => c_state_28_port, QN => n60);
   c_state_reg_29_inst : DFFR_X1 port map( D => n_state_29_port, CK => clk, RN 
                           => n175, Q => c_state_29_port, QN => net164133);
   c_state_reg_30_inst : DFFR_X1 port map( D => n_state_30_port, CK => clk, RN 
                           => n174, Q => c_state_30_port, QN => net108733);
   c_state_reg_31_inst : DFFR_X1 port map( D => n_state_31_port, CK => clk, RN 
                           => n174, Q => c_state_31_port, QN => n53_port);
   adj_final_mod_reg_31_inst : DFF_X1 port map( D => n210, CK => clk, Q => 
                           adj_final_mod_31_port, QN => n189);
   adj_final_mod_reg_30_inst : DFF_X1 port map( D => n209, CK => clk, Q => 
                           adj_final_mod_30_port, QN => n188);
   adj_final_mod_reg_29_inst : DFF_X1 port map( D => n208, CK => clk, Q => 
                           adj_final_mod_29_port, QN => net108732);
   adj_final_mod_reg_28_inst : DFF_X1 port map( D => n207, CK => clk, Q => 
                           adj_final_mod_28_port, QN => net108731);
   adj_final_mod_reg_27_inst : DFF_X1 port map( D => n206, CK => clk, Q => 
                           adj_final_mod_27_port, QN => net108730);
   adj_final_mod_reg_26_inst : DFF_X1 port map( D => n205, CK => clk, Q => 
                           adj_final_mod_26_port, QN => net108729);
   adj_final_mod_reg_25_inst : DFF_X1 port map( D => n204, CK => clk, Q => 
                           adj_final_mod_25_port, QN => net108728);
   adj_final_mod_reg_24_inst : DFF_X1 port map( D => n203, CK => clk, Q => 
                           adj_final_mod_24_port, QN => net108727);
   adj_final_mod_reg_23_inst : DFF_X1 port map( D => n202, CK => clk, Q => 
                           adj_final_mod_23_port, QN => net108726);
   adj_final_mod_reg_22_inst : DFF_X1 port map( D => n201, CK => clk, Q => 
                           adj_final_mod_22_port, QN => net108725);
   adj_final_mod_reg_21_inst : DFF_X1 port map( D => n200, CK => clk, Q => 
                           adj_final_mod_21_port, QN => net108724);
   adj_final_mod_reg_20_inst : DFF_X1 port map( D => n199, CK => clk, Q => 
                           adj_final_mod_20_port, QN => net108723);
   adj_final_mod_reg_19_inst : DFF_X1 port map( D => n198, CK => clk, Q => 
                           adj_final_mod_19_port, QN => net108722);
   adj_final_mod_reg_18_inst : DFF_X1 port map( D => n197, CK => clk, Q => 
                           adj_final_mod_18_port, QN => net108721);
   adj_final_mod_reg_17_inst : DFF_X1 port map( D => n196, CK => clk, Q => 
                           adj_final_mod_17_port, QN => net108720);
   adj_final_mod_reg_16_inst : DFF_X1 port map( D => n195, CK => clk, Q => 
                           adj_final_mod_16_port, QN => net108719);
   adj_final_mod_reg_15_inst : DFF_X1 port map( D => n194, CK => clk, Q => 
                           adj_final_mod_15_port, QN => net108718);
   e_a_reg_0_inst : DFF_X1 port map( D => N9, CK => clk, Q => e_a_0_port, QN =>
                           net108717);
   e_b_reg_16_inst : DFF_X1 port map( D => N57, CK => clk, Q => e_b_16_port, QN
                           => net108716);
   e_b_reg_15_inst : DFF_X1 port map( D => N56, CK => clk, Q => e_b_15_port, QN
                           => net108715);
   e_b_reg_14_inst : DFF_X1 port map( D => N55, CK => clk, Q => e_b_14_port, QN
                           => net108714);
   e_b_reg_13_inst : DFF_X1 port map( D => N54, CK => clk, Q => e_b_13_port, QN
                           => net108713);
   e_b_reg_12_inst : DFF_X1 port map( D => N53, CK => clk, Q => e_b_12_port, QN
                           => net108712);
   e_b_reg_11_inst : DFF_X1 port map( D => N52, CK => clk, Q => e_b_11_port, QN
                           => net108711);
   e_b_reg_10_inst : DFF_X1 port map( D => N51, CK => clk, Q => e_b_10_port, QN
                           => net108710);
   e_b_reg_9_inst : DFF_X1 port map( D => N50, CK => clk, Q => e_b_9_port, QN 
                           => net108709);
   e_b_reg_8_inst : DFF_X1 port map( D => N49, CK => clk, Q => e_b_8_port, QN 
                           => net108708);
   e_b_reg_7_inst : DFF_X1 port map( D => N48, CK => clk, Q => e_b_7_port, QN 
                           => net108707);
   e_b_reg_6_inst : DFF_X1 port map( D => N47, CK => clk, Q => e_b_6_port, QN 
                           => net108706);
   e_b_reg_5_inst : DFF_X1 port map( D => N46, CK => clk, Q => e_b_5_port, QN 
                           => net108705);
   e_b_reg_4_inst : DFF_X1 port map( D => N45, CK => clk, Q => e_b_4_port, QN 
                           => net108704);
   e_b_reg_3_inst : DFF_X1 port map( D => N44, CK => clk, Q => e_b_3_port, QN 
                           => net108703);
   e_b_reg_2_inst : DFF_X1 port map( D => N43, CK => clk, Q => e_b_2_port, QN 
                           => n58);
   e_b_reg_0_inst : DFF_X1 port map( D => N41, CK => clk, Q => e_b_0_port, QN 
                           => n193);
   e_b_reg_1_inst : DFF_X1 port map( D => N42, CK => clk, Q => e_b_1_port, QN 
                           => n192);
   e_a_reg_2_inst : DFF_X1 port map( D => N11, CK => clk, Q => e_a_2_port, QN 
                           => net108702);
   e_a_reg_4_inst : DFF_X1 port map( D => N13, CK => clk, Q => e_a_4_port, QN 
                           => net108701);
   e_a_reg_6_inst : DFF_X1 port map( D => N15, CK => clk, Q => e_a_6_port, QN 
                           => net108700);
   e_a_reg_8_inst : DFF_X1 port map( D => N17, CK => clk, Q => e_a_8_port, QN 
                           => net108699);
   e_a_reg_10_inst : DFF_X1 port map( D => N19, CK => clk, Q => e_a_10_port, QN
                           => net108698);
   e_a_reg_12_inst : DFF_X1 port map( D => N21, CK => clk, Q => e_a_12_port, QN
                           => net108697);
   e_a_reg_14_inst : DFF_X1 port map( D => N23, CK => clk, Q => e_a_14_port, QN
                           => n65);
   e_a_reg_16_inst : DFF_X1 port map( D => N25, CK => clk, Q => e_a_16_port, QN
                           => n66);
   e_a_reg_18_inst : DFF_X1 port map( D => N27, CK => clk, Q => e_a_18_port, QN
                           => n67);
   e_a_reg_20_inst : DFF_X1 port map( D => N29, CK => clk, Q => e_a_20_port, QN
                           => n68);
   e_a_reg_22_inst : DFF_X1 port map( D => N31, CK => clk, Q => e_a_22_port, QN
                           => n69);
   e_a_reg_24_inst : DFF_X1 port map( D => N33, CK => clk, Q => e_a_24_port, QN
                           => n70_port);
   e_a_reg_26_inst : DFF_X1 port map( D => N35, CK => clk, Q => e_a_26_port, QN
                           => n71_port);
   e_a_reg_28_inst : DFF_X1 port map( D => N37, CK => clk, Q => e_a_28_port, QN
                           => n72_port);
   e_a_reg_30_inst : DFF_X1 port map( D => N39, CK => clk, Q => e_a_30_port, QN
                           => n191);
   e_a_reg_1_inst : DFF_X1 port map( D => N10, CK => clk, Q => e_a_1_port, QN 
                           => net108696);
   e_a_reg_3_inst : DFF_X1 port map( D => N12, CK => clk, Q => e_a_3_port, QN 
                           => net108695);
   e_a_reg_5_inst : DFF_X1 port map( D => N14, CK => clk, Q => e_a_5_port, QN 
                           => net108694);
   e_a_reg_7_inst : DFF_X1 port map( D => N16, CK => clk, Q => e_a_7_port, QN 
                           => net108693);
   e_a_reg_9_inst : DFF_X1 port map( D => N18, CK => clk, Q => e_a_9_port, QN 
                           => net108692);
   e_a_reg_11_inst : DFF_X1 port map( D => N20, CK => clk, Q => e_a_11_port, QN
                           => net108691);
   e_a_reg_13_inst : DFF_X1 port map( D => N22, CK => clk, Q => e_a_13_port, QN
                           => n79_port);
   e_a_reg_15_inst : DFF_X1 port map( D => N24, CK => clk, Q => e_a_15_port, QN
                           => n80_port);
   e_a_reg_17_inst : DFF_X1 port map( D => N26, CK => clk, Q => e_a_17_port, QN
                           => n81_port);
   e_a_reg_19_inst : DFF_X1 port map( D => N28, CK => clk, Q => e_a_19_port, QN
                           => n82_port);
   e_a_reg_21_inst : DFF_X1 port map( D => N30, CK => clk, Q => e_a_21_port, QN
                           => n83_port);
   e_a_reg_23_inst : DFF_X1 port map( D => N32, CK => clk, Q => e_a_23_port, QN
                           => n84_port);
   e_a_reg_25_inst : DFF_X1 port map( D => N34, CK => clk, Q => e_a_25_port, QN
                           => n85_port);
   e_a_reg_27_inst : DFF_X1 port map( D => N36, CK => clk, Q => e_a_27_port, QN
                           => n86_port);
   e_a_reg_29_inst : DFF_X1 port map( D => N38, CK => clk, Q => e_a_29_port, QN
                           => n87_port);
   e_a_reg_31_inst : DFF_X1 port map( D => N40, CK => clk, Q => e_a_31_port, QN
                           => n190);
   adj_final_mod_0_port <= '0';
   adj_final_mod_1_port <= '0';
   adj_final_mod_2_port <= '0';
   adj_final_mod_3_port <= '0';
   adj_final_mod_4_port <= '0';
   adj_final_mod_5_port <= '0';
   adj_final_mod_6_port <= '0';
   adj_final_mod_7_port <= '0';
   adj_final_mod_8_port <= '0';
   adj_final_mod_9_port <= '0';
   adj_final_mod_10_port <= '0';
   adj_final_mod_11_port <= '0';
   adj_final_mod_12_port <= '0';
   adj_final_mod_13_port <= '0';
   adj_final_mod_14_port <= '0';
   U203 : XOR2_X1 port map( A => adj_sum_15_port, B => adj_cout, Z => n96_port)
                           ;
   U205 : NAND3_X1 port map( A1 => net108734, A2 => net108733, A3 => net108735,
                           ZN => n156);
   ADJUST0 : Adder_DATA_SIZE16 port map( cin => X_Logic0_port, a(15) => a(15), 
                           a(14) => a(14), a(13) => a(13), a(12) => a(12), 
                           a(11) => a(11), a(10) => a(10), a(9) => a(9), a(8) 
                           => a(8), a(7) => a(7), a(6) => a(6), a(5) => a(5), 
                           a(4) => a(4), a(3) => a(3), a(2) => a(2), a(1) => 
                           a(1), a(0) => a(0), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           s(15) => adj_sum_15_port, s(14) => adj_sum_14_port, 
                           s(13) => adj_sum_13_port, s(12) => adj_sum_12_port, 
                           s(11) => adj_sum_11_port, s(10) => adj_sum_10_port, 
                           s(9) => adj_sum_9_port, s(8) => adj_sum_8_port, s(7)
                           => adj_sum_7_port, s(6) => adj_sum_6_port, s(5) => 
                           adj_sum_5_port, s(4) => adj_sum_4_port, s(3) => 
                           adj_sum_3_port, s(2) => adj_sum_2_port, s(1) => 
                           adj_sum_1_port, s(0) => adj_sum_0_port, cout => 
                           adj_cout);
   BEC0 : BoothEncoder port map( din(2) => e_b_2_port, din(1) => e_b_1_port, 
                           din(0) => e_b_0_port, sel(2) => sel_2_port, sel(1) 
                           => sel_1_port, sel(0) => sel_0_port);
   MUX0 : Mux_DATA_SIZE32_1 port map( sel => sel_0_port, din0(31) => 
                           e_a_31_port, din0(30) => e_a_30_port, din0(29) => 
                           e_a_29_port, din0(28) => e_a_28_port, din0(27) => 
                           e_a_27_port, din0(26) => e_a_26_port, din0(25) => 
                           e_a_25_port, din0(24) => e_a_24_port, din0(23) => 
                           e_a_23_port, din0(22) => e_a_22_port, din0(21) => 
                           e_a_21_port, din0(20) => e_a_20_port, din0(19) => 
                           e_a_19_port, din0(18) => e_a_18_port, din0(17) => 
                           e_a_17_port, din0(16) => e_a_16_port, din0(15) => 
                           e_a_15_port, din0(14) => e_a_14_port, din0(13) => 
                           e_a_13_port, din0(12) => e_a_12_port, din0(11) => 
                           e_a_11_port, din0(10) => e_a_10_port, din0(9) => 
                           e_a_9_port, din0(8) => e_a_8_port, din0(7) => 
                           e_a_7_port, din0(6) => e_a_6_port, din0(5) => 
                           e_a_5_port, din0(4) => e_a_4_port, din0(3) => 
                           e_a_3_port, din0(2) => e_a_2_port, din0(1) => 
                           e_a_1_port, din0(0) => e_a_0_port, din1(31) => 
                           e_a_30_port, din1(30) => e_a_29_port, din1(29) => 
                           e_a_28_port, din1(28) => e_a_27_port, din1(27) => 
                           e_a_26_port, din1(26) => e_a_25_port, din1(25) => 
                           e_a_24_port, din1(24) => e_a_23_port, din1(23) => 
                           e_a_22_port, din1(22) => e_a_21_port, din1(21) => 
                           e_a_20_port, din1(20) => e_a_19_port, din1(19) => 
                           e_a_18_port, din1(18) => e_a_17_port, din1(17) => 
                           e_a_16_port, din1(16) => e_a_15_port, din1(15) => 
                           e_a_14_port, din1(14) => e_a_13_port, din1(13) => 
                           e_a_12_port, din1(12) => e_a_11_port, din1(11) => 
                           e_a_10_port, din1(10) => e_a_9_port, din1(9) => 
                           e_a_8_port, din1(8) => e_a_7_port, din1(7) => 
                           e_a_6_port, din1(6) => e_a_5_port, din1(5) => 
                           e_a_4_port, din1(4) => e_a_3_port, din1(3) => 
                           e_a_2_port, din1(2) => e_a_1_port, din1(1) => 
                           e_a_0_port, din1(0) => X_Logic0_port, dout(31) => 
                           mux_out_31_port, dout(30) => mux_out_30_port, 
                           dout(29) => mux_out_29_port, dout(28) => 
                           mux_out_28_port, dout(27) => mux_out_27_port, 
                           dout(26) => mux_out_26_port, dout(25) => 
                           mux_out_25_port, dout(24) => mux_out_24_port, 
                           dout(23) => mux_out_23_port, dout(22) => 
                           mux_out_22_port, dout(21) => mux_out_21_port, 
                           dout(20) => mux_out_20_port, dout(19) => 
                           mux_out_19_port, dout(18) => mux_out_18_port, 
                           dout(17) => mux_out_17_port, dout(16) => 
                           mux_out_16_port, dout(15) => mux_out_15_port, 
                           dout(14) => mux_out_14_port, dout(13) => 
                           mux_out_13_port, dout(12) => mux_out_12_port, 
                           dout(11) => mux_out_11_port, dout(10) => 
                           mux_out_10_port, dout(9) => mux_out_9_port, dout(8) 
                           => mux_out_8_port, dout(7) => mux_out_7_port, 
                           dout(6) => mux_out_6_port, dout(5) => mux_out_5_port
                           , dout(4) => mux_out_4_port, dout(3) => 
                           mux_out_3_port, dout(2) => mux_out_2_port, dout(1) 
                           => mux_out_1_port, dout(0) => mux_out_0_port);
   ADDSUBn : AddSub_DATA_SIZE32_1 port map( as => sel_1_port, a(31) => 
                           add_out_reg_31_port, a(30) => add_out_reg_30_port, 
                           a(29) => add_out_reg_29_port, a(28) => 
                           add_out_reg_28_port, a(27) => add_out_reg_27_port, 
                           a(26) => add_out_reg_26_port, a(25) => 
                           add_out_reg_25_port, a(24) => add_out_reg_24_port, 
                           a(23) => add_out_reg_23_port, a(22) => 
                           add_out_reg_22_port, a(21) => add_out_reg_21_port, 
                           a(20) => add_out_reg_20_port, a(19) => 
                           add_out_reg_19_port, a(18) => add_out_reg_18_port, 
                           a(17) => add_out_reg_17_port, a(16) => 
                           add_out_reg_16_port, a(15) => add_out_reg_15_port, 
                           a(14) => add_out_reg_14_port, a(13) => 
                           add_out_reg_13_port, a(12) => add_out_reg_12_port, 
                           a(11) => add_out_reg_11_port, a(10) => 
                           add_out_reg_10_port, a(9) => add_out_reg_9_port, 
                           a(8) => add_out_reg_8_port, a(7) => 
                           add_out_reg_7_port, a(6) => add_out_reg_6_port, a(5)
                           => add_out_reg_5_port, a(4) => add_out_reg_4_port, 
                           a(3) => add_out_reg_3_port, a(2) => 
                           add_out_reg_2_port, a(1) => add_out_reg_1_port, a(0)
                           => add_out_reg_0_port, b(31) => zero_out_31_port, 
                           b(30) => zero_out_30_port, b(29) => zero_out_29_port
                           , b(28) => zero_out_28_port, b(27) => 
                           zero_out_27_port, b(26) => zero_out_26_port, b(25) 
                           => zero_out_25_port, b(24) => zero_out_24_port, 
                           b(23) => zero_out_23_port, b(22) => zero_out_22_port
                           , b(21) => zero_out_21_port, b(20) => 
                           zero_out_20_port, b(19) => zero_out_19_port, b(18) 
                           => zero_out_18_port, b(17) => zero_out_17_port, 
                           b(16) => zero_out_16_port, b(15) => zero_out_15_port
                           , b(14) => zero_out_14_port, b(13) => 
                           zero_out_13_port, b(12) => zero_out_12_port, b(11) 
                           => zero_out_11_port, b(10) => zero_out_10_port, b(9)
                           => zero_out_9_port, b(8) => zero_out_8_port, b(7) =>
                           zero_out_7_port, b(6) => zero_out_6_port, b(5) => 
                           zero_out_5_port, b(4) => zero_out_4_port, b(3) => 
                           zero_out_3_port, b(2) => zero_out_2_port, b(1) => 
                           zero_out_1_port, b(0) => zero_out_0_port, re(31) => 
                           add_out_31_port, re(30) => add_out_30_port, re(29) 
                           => add_out_29_port, re(28) => add_out_28_port, 
                           re(27) => add_out_27_port, re(26) => add_out_26_port
                           , re(25) => add_out_25_port, re(24) => 
                           add_out_24_port, re(23) => add_out_23_port, re(22) 
                           => add_out_22_port, re(21) => add_out_21_port, 
                           re(20) => add_out_20_port, re(19) => add_out_19_port
                           , re(18) => add_out_18_port, re(17) => 
                           add_out_17_port, re(16) => add_out_16_port, re(15) 
                           => add_out_15_port, re(14) => add_out_14_port, 
                           re(13) => add_out_13_port, re(12) => add_out_12_port
                           , re(11) => add_out_11_port, re(10) => 
                           add_out_10_port, re(9) => add_out_9_port, re(8) => 
                           add_out_8_port, re(7) => add_out_7_port, re(6) => 
                           add_out_6_port, re(5) => add_out_5_port, re(4) => 
                           add_out_4_port, re(3) => add_out_3_port, re(2) => 
                           add_out_2_port, re(1) => add_out_1_port, re(0) => 
                           add_out_0_port, cout => net4348);
   REG0 : Reg_DATA_SIZE32_1 port map( rst => reg_rst, en => en_o, clk => clk, 
                           din(31) => add_out_31_port, din(30) => 
                           add_out_30_port, din(29) => add_out_29_port, din(28)
                           => add_out_28_port, din(27) => add_out_27_port, 
                           din(26) => add_out_26_port, din(25) => 
                           add_out_25_port, din(24) => add_out_24_port, din(23)
                           => add_out_23_port, din(22) => add_out_22_port, 
                           din(21) => add_out_21_port, din(20) => 
                           add_out_20_port, din(19) => add_out_19_port, din(18)
                           => add_out_18_port, din(17) => add_out_17_port, 
                           din(16) => add_out_16_port, din(15) => 
                           add_out_15_port, din(14) => add_out_14_port, din(13)
                           => add_out_13_port, din(12) => add_out_12_port, 
                           din(11) => add_out_11_port, din(10) => 
                           add_out_10_port, din(9) => add_out_9_port, din(8) =>
                           add_out_8_port, din(7) => add_out_7_port, din(6) => 
                           add_out_6_port, din(5) => add_out_5_port, din(4) => 
                           add_out_4_port, din(3) => add_out_3_port, din(2) => 
                           add_out_2_port, din(1) => add_out_1_port, din(0) => 
                           add_out_0_port, dout(31) => add_out_reg_31_port, 
                           dout(30) => add_out_reg_30_port, dout(29) => 
                           add_out_reg_29_port, dout(28) => add_out_reg_28_port
                           , dout(27) => add_out_reg_27_port, dout(26) => 
                           add_out_reg_26_port, dout(25) => add_out_reg_25_port
                           , dout(24) => add_out_reg_24_port, dout(23) => 
                           add_out_reg_23_port, dout(22) => add_out_reg_22_port
                           , dout(21) => add_out_reg_21_port, dout(20) => 
                           add_out_reg_20_port, dout(19) => add_out_reg_19_port
                           , dout(18) => add_out_reg_18_port, dout(17) => 
                           add_out_reg_17_port, dout(16) => add_out_reg_16_port
                           , dout(15) => add_out_reg_15_port, dout(14) => 
                           add_out_reg_14_port, dout(13) => add_out_reg_13_port
                           , dout(12) => add_out_reg_12_port, dout(11) => 
                           add_out_reg_11_port, dout(10) => add_out_reg_10_port
                           , dout(9) => add_out_reg_9_port, dout(8) => 
                           add_out_reg_8_port, dout(7) => add_out_reg_7_port, 
                           dout(6) => add_out_reg_6_port, dout(5) => 
                           add_out_reg_5_port, dout(4) => add_out_reg_4_port, 
                           dout(3) => add_out_reg_3_port, dout(2) => 
                           add_out_reg_2_port, dout(1) => add_out_reg_1_port, 
                           dout(0) => add_out_reg_0_port);
   ADJUST1 : Adder_DATA_SIZE32_5 port map( cin => X_Logic0_port, a(31) => 
                           add_out_reg_31_port, a(30) => add_out_reg_30_port, 
                           a(29) => add_out_reg_29_port, a(28) => 
                           add_out_reg_28_port, a(27) => add_out_reg_27_port, 
                           a(26) => add_out_reg_26_port, a(25) => 
                           add_out_reg_25_port, a(24) => add_out_reg_24_port, 
                           a(23) => add_out_reg_23_port, a(22) => 
                           add_out_reg_22_port, a(21) => add_out_reg_21_port, 
                           a(20) => add_out_reg_20_port, a(19) => 
                           add_out_reg_19_port, a(18) => add_out_reg_18_port, 
                           a(17) => add_out_reg_17_port, a(16) => 
                           add_out_reg_16_port, a(15) => add_out_reg_15_port, 
                           a(14) => add_out_reg_14_port, a(13) => 
                           add_out_reg_13_port, a(12) => add_out_reg_12_port, 
                           a(11) => add_out_reg_11_port, a(10) => 
                           add_out_reg_10_port, a(9) => add_out_reg_9_port, 
                           a(8) => add_out_reg_8_port, a(7) => 
                           add_out_reg_7_port, a(6) => add_out_reg_6_port, a(5)
                           => add_out_reg_5_port, a(4) => add_out_reg_4_port, 
                           a(3) => add_out_reg_3_port, a(2) => 
                           add_out_reg_2_port, a(1) => add_out_reg_1_port, a(0)
                           => add_out_reg_0_port, b(31) => 
                           adj_final_mod_31_port, b(30) => 
                           adj_final_mod_30_port, b(29) => 
                           adj_final_mod_29_port, b(28) => 
                           adj_final_mod_28_port, b(27) => 
                           adj_final_mod_27_port, b(26) => 
                           adj_final_mod_26_port, b(25) => 
                           adj_final_mod_25_port, b(24) => 
                           adj_final_mod_24_port, b(23) => 
                           adj_final_mod_23_port, b(22) => 
                           adj_final_mod_22_port, b(21) => 
                           adj_final_mod_21_port, b(20) => 
                           adj_final_mod_20_port, b(19) => 
                           adj_final_mod_19_port, b(18) => 
                           adj_final_mod_18_port, b(17) => 
                           adj_final_mod_17_port, b(16) => 
                           adj_final_mod_16_port, b(15) => 
                           adj_final_mod_15_port, b(14) => 
                           adj_final_mod_14_port, b(13) => 
                           adj_final_mod_13_port, b(12) => 
                           adj_final_mod_12_port, b(11) => 
                           adj_final_mod_11_port, b(10) => 
                           adj_final_mod_10_port, b(9) => adj_final_mod_9_port,
                           b(8) => adj_final_mod_8_port, b(7) => 
                           adj_final_mod_7_port, b(6) => adj_final_mod_6_port, 
                           b(5) => adj_final_mod_5_port, b(4) => 
                           adj_final_mod_4_port, b(3) => adj_final_mod_3_port, 
                           b(2) => adj_final_mod_2_port, b(1) => 
                           adj_final_mod_1_port, b(0) => adj_final_mod_0_port, 
                           s(31) => o(31), s(30) => o(30), s(29) => o(29), 
                           s(28) => o(28), s(27) => o(27), s(26) => o(26), 
                           s(25) => o(25), s(24) => o(24), s(23) => o(23), 
                           s(22) => o(22), s(21) => o(21), s(20) => o(20), 
                           s(19) => o(19), s(18) => o(18), s(17) => o(17), 
                           s(16) => o(16), s(15) => o(15), s(14) => o(14), 
                           s(13) => o(13), s(12) => o(12), s(11) => o(11), 
                           s(10) => o(10), s(9) => o(9), s(8) => o(8), s(7) => 
                           o(7), s(6) => o(6), s(5) => o(5), s(4) => o(4), s(3)
                           => o(3), s(2) => o(2), s(1) => o(1), s(0) => o(0), 
                           cout => net4347);
   add_189 : BoothMul_DATA_SIZE16_STAGE10_DW01_inc_0 port map( A(31) => 
                           c_state_31_port, A(30) => c_state_30_port, A(29) => 
                           c_state_29_port, A(28) => c_state_28_port, A(27) => 
                           c_state_27_port, A(26) => c_state_26_port, A(25) => 
                           c_state_25_port, A(24) => c_state_24_port, A(23) => 
                           c_state_23_port, A(22) => c_state_22_port, A(21) => 
                           c_state_21_port, A(20) => c_state_20_port, A(19) => 
                           c_state_19_port, A(18) => c_state_18_port, A(17) => 
                           c_state_17_port, A(16) => c_state_16_port, A(15) => 
                           c_state_15_port, A(14) => c_state_14_port, A(13) => 
                           c_state_13_port, A(12) => c_state_12_port, A(11) => 
                           c_state_11_port, A(10) => c_state_10_port, A(9) => 
                           c_state_9_port, A(8) => c_state_8_port, A(7) => 
                           c_state_7_port, A(6) => c_state_6_port, A(5) => 
                           c_state_5_port, A(4) => c_state_4_port, A(3) => 
                           c_state_3_port, A(2) => c_state_2_port, A(1) => 
                           c_state_1_port, A(0) => c_state_0_port, SUM(31) => 
                           N101, SUM(30) => N100, SUM(29) => N99, SUM(28) => 
                           N98, SUM(27) => N97, SUM(26) => N96, SUM(25) => N95,
                           SUM(24) => N94, SUM(23) => N93, SUM(22) => N92, 
                           SUM(21) => N91, SUM(20) => N90, SUM(19) => N89, 
                           SUM(18) => N88, SUM(17) => N87, SUM(16) => N86, 
                           SUM(15) => N85, SUM(14) => N84, SUM(13) => N83, 
                           SUM(12) => N82, SUM(11) => N81, SUM(10) => N80, 
                           SUM(9) => N79, SUM(8) => N78, SUM(7) => N77, SUM(6) 
                           => N76, SUM(5) => N75, SUM(4) => N74, SUM(3) => N73,
                           SUM(2) => N72, SUM(1) => N71, SUM(0) => N70);
   U3 : AND2_X1 port map( A1 => mux_out_0_port, A2 => n171, ZN => 
                           zero_out_0_port);
   U4 : BUF_X2 port map( A => sel_2_port, Z => n171);
   U5 : INV_X1 port map( A => n159, ZN => n147);
   U6 : INV_X1 port map( A => n162, ZN => n157);
   U7 : BUF_X1 port map( A => n64, Z => n158);
   U8 : BUF_X1 port map( A => n64, Z => n160);
   U9 : BUF_X1 port map( A => n64, Z => n159);
   U10 : BUF_X1 port map( A => n73_port, Z => n162);
   U11 : BUF_X1 port map( A => n73_port, Z => n161);
   U12 : BUF_X1 port map( A => n73_port, Z => n163);
   U13 : BUF_X1 port map( A => n74_port, Z => n166);
   U14 : BUF_X1 port map( A => n74_port, Z => n165);
   U15 : BUF_X1 port map( A => n74_port, Z => n164);
   U16 : BUF_X1 port map( A => n75_port, Z => n167);
   U17 : BUF_X1 port map( A => n75_port, Z => n168);
   U18 : INV_X1 port map( A => n97_port, ZN => n95_port);
   U19 : BUF_X1 port map( A => n94_port, Z => n73_port);
   U20 : BUF_X1 port map( A => n94_port, Z => n64);
   U21 : BUF_X1 port map( A => n76_port, Z => n74_port);
   U22 : BUF_X1 port map( A => n76_port, Z => n75_port);
   U23 : NOR2_X2 port map( A1 => n158, A2 => sign, ZN => n97_port);
   U24 : BUF_X1 port map( A => n99_port, Z => n94_port);
   U25 : BUF_X1 port map( A => n99_port, Z => n76_port);
   U26 : AND2_X1 port map( A1 => n176, A2 => en_o, ZN => reg_rst);
   U27 : CLKBUF_X1 port map( A => sel_2_port, Z => n172);
   U28 : CLKBUF_X1 port map( A => sel_2_port, Z => n173);
   U29 : AND2_X1 port map( A1 => N100, A2 => n170, ZN => n_state_30_port);
   U30 : AND2_X1 port map( A1 => N98, A2 => n170, ZN => n_state_28_port);
   U31 : AND2_X1 port map( A1 => N97, A2 => n170, ZN => n_state_27_port);
   U32 : AND2_X1 port map( A1 => N96, A2 => n170, ZN => n_state_26_port);
   U33 : AND2_X1 port map( A1 => N93, A2 => n169, ZN => n_state_23_port);
   U34 : AND2_X1 port map( A1 => N92, A2 => n169, ZN => n_state_22_port);
   U35 : AND2_X1 port map( A1 => N99, A2 => n170, ZN => n_state_29_port);
   U36 : AND2_X1 port map( A1 => N95, A2 => n169, ZN => n_state_25_port);
   U37 : AND2_X1 port map( A1 => N94, A2 => n169, ZN => n_state_24_port);
   U38 : BUF_X1 port map( A => n77_port, Z => n169);
   U39 : BUF_X1 port map( A => n77_port, Z => n170);
   U40 : INV_X1 port map( A => n114, ZN => en_o);
   U41 : NAND2_X1 port map( A1 => en, A2 => n114, ZN => n99_port);
   U42 : NOR2_X1 port map( A1 => lock, A2 => n90_port, ZN => n89_port);
   U43 : INV_X1 port map( A => n91_port, ZN => n90_port);
   U44 : AND3_X1 port map( A1 => b(15), A2 => n157, A3 => sign, ZN => N57);
   U45 : AND2_X1 port map( A1 => b(14), A2 => n157, ZN => N56);
   U46 : AND2_X1 port map( A1 => N91, A2 => n169, ZN => n_state_21_port);
   U47 : AND2_X1 port map( A1 => N90, A2 => n169, ZN => n_state_20_port);
   U48 : AND2_X1 port map( A1 => N83, A2 => n169, ZN => n_state_13_port);
   U49 : AND2_X1 port map( A1 => N82, A2 => n169, ZN => n_state_12_port);
   U50 : AND2_X1 port map( A1 => N81, A2 => n169, ZN => n_state_11_port);
   U51 : AND2_X1 port map( A1 => N79, A2 => n170, ZN => n_state_9_port);
   U52 : AND2_X1 port map( A1 => N75, A2 => n170, ZN => n_state_5_port);
   U53 : AND2_X1 port map( A1 => N74, A2 => n170, ZN => n_state_4_port);
   U54 : AND2_X1 port map( A1 => N73, A2 => n170, ZN => n_state_3_port);
   U55 : AND2_X1 port map( A1 => N72, A2 => n170, ZN => n_state_2_port);
   U56 : AND2_X1 port map( A1 => N71, A2 => n169, ZN => n_state_1_port);
   U57 : AND2_X1 port map( A1 => N80, A2 => n169, ZN => n_state_10_port);
   U58 : AND2_X1 port map( A1 => N89, A2 => n169, ZN => n_state_19_port);
   U59 : AND2_X1 port map( A1 => N88, A2 => n169, ZN => n_state_18_port);
   U60 : AND2_X1 port map( A1 => N87, A2 => n169, ZN => n_state_17_port);
   U61 : AND2_X1 port map( A1 => N86, A2 => n169, ZN => n_state_16_port);
   U62 : AND2_X1 port map( A1 => N85, A2 => n169, ZN => n_state_15_port);
   U63 : AND2_X1 port map( A1 => N84, A2 => n169, ZN => n_state_14_port);
   U64 : AND2_X1 port map( A1 => N78, A2 => n170, ZN => n_state_8_port);
   U65 : AND2_X1 port map( A1 => N77, A2 => n170, ZN => n_state_7_port);
   U66 : AND2_X1 port map( A1 => N76, A2 => n170, ZN => n_state_6_port);
   U67 : BUF_X1 port map( A => rst, Z => n175);
   U68 : BUF_X1 port map( A => rst, Z => n174);
   U69 : BUF_X1 port map( A => rst, Z => n176);
   U70 : AND2_X1 port map( A1 => mux_out_5_port, A2 => n173, ZN => 
                           zero_out_5_port);
   U71 : AND2_X1 port map( A1 => mux_out_10_port, A2 => n171, ZN => 
                           zero_out_10_port);
   U72 : AND2_X1 port map( A1 => mux_out_19_port, A2 => n171, ZN => 
                           zero_out_19_port);
   U73 : AND2_X1 port map( A1 => mux_out_18_port, A2 => n171, ZN => 
                           zero_out_18_port);
   U74 : AND2_X1 port map( A1 => mux_out_21_port, A2 => n172, ZN => 
                           zero_out_21_port);
   U75 : AND2_X1 port map( A1 => mux_out_11_port, A2 => n171, ZN => 
                           zero_out_11_port);
   U76 : AND2_X1 port map( A1 => mux_out_7_port, A2 => n173, ZN => 
                           zero_out_7_port);
   U77 : AND2_X1 port map( A1 => mux_out_13_port, A2 => n171, ZN => 
                           zero_out_13_port);
   U78 : AND2_X1 port map( A1 => mux_out_14_port, A2 => n171, ZN => 
                           zero_out_14_port);
   U79 : AND2_X1 port map( A1 => mux_out_16_port, A2 => n171, ZN => 
                           zero_out_16_port);
   U80 : AND2_X1 port map( A1 => mux_out_17_port, A2 => n171, ZN => 
                           zero_out_17_port);
   U81 : AND2_X1 port map( A1 => mux_out_3_port, A2 => n173, ZN => 
                           zero_out_3_port);
   U82 : AND2_X1 port map( A1 => mux_out_1_port, A2 => n171, ZN => 
                           zero_out_1_port);
   U83 : AND2_X1 port map( A1 => mux_out_8_port, A2 => n173, ZN => 
                           zero_out_8_port);
   U84 : AND2_X1 port map( A1 => mux_out_2_port, A2 => n172, ZN => 
                           zero_out_2_port);
   U85 : AND2_X1 port map( A1 => mux_out_12_port, A2 => n171, ZN => 
                           zero_out_12_port);
   U86 : AND2_X1 port map( A1 => mux_out_20_port, A2 => n172, ZN => 
                           zero_out_20_port);
   U87 : AND2_X1 port map( A1 => mux_out_6_port, A2 => n173, ZN => 
                           zero_out_6_port);
   U88 : AND2_X1 port map( A1 => mux_out_15_port, A2 => n171, ZN => 
                           zero_out_15_port);
   U89 : AND2_X1 port map( A1 => n173, A2 => mux_out_9_port, ZN => 
                           zero_out_9_port);
   U90 : OAI22_X1 port map( A1 => n189, A2 => n157, B1 => n95_port, B2 => 
                           n96_port, ZN => n210);
   U91 : OAI22_X1 port map( A1 => n188, A2 => n157, B1 => adj_sum_15_port, B2 
                           => n95_port, ZN => n209);
   U92 : AND2_X1 port map( A1 => mux_out_4_port, A2 => n173, ZN => 
                           zero_out_4_port);
   U93 : INV_X1 port map( A => n105, ZN => n202);
   U94 : AOI22_X1 port map( A1 => adj_sum_8_port, A2 => n97_port, B1 => n159, 
                           B2 => adj_final_mod_23_port, ZN => n105);
   U95 : INV_X1 port map( A => n104, ZN => n203);
   U96 : AOI22_X1 port map( A1 => adj_sum_9_port, A2 => n97_port, B1 => n159, 
                           B2 => adj_final_mod_24_port, ZN => n104);
   U97 : INV_X1 port map( A => n103, ZN => n204);
   U98 : AOI22_X1 port map( A1 => adj_sum_10_port, A2 => n97_port, B1 => n158, 
                           B2 => adj_final_mod_25_port, ZN => n103);
   U99 : INV_X1 port map( A => n102, ZN => n205);
   U100 : AOI22_X1 port map( A1 => adj_sum_11_port, A2 => n97_port, B1 => n159,
                           B2 => adj_final_mod_26_port, ZN => n102);
   U101 : INV_X1 port map( A => n101_port, ZN => n206);
   U102 : AOI22_X1 port map( A1 => adj_sum_12_port, A2 => n97_port, B1 => n158,
                           B2 => adj_final_mod_27_port, ZN => n101_port);
   U103 : INV_X1 port map( A => n100_port, ZN => n207);
   U104 : AOI22_X1 port map( A1 => adj_sum_13_port, A2 => n97_port, B1 => n158,
                           B2 => adj_final_mod_28_port, ZN => n100_port);
   U105 : INV_X1 port map( A => n98_port, ZN => n208);
   U106 : AOI22_X1 port map( A1 => adj_sum_14_port, A2 => n97_port, B1 => n163,
                           B2 => adj_final_mod_29_port, ZN => n98_port);
   U107 : AND2_X1 port map( A1 => N101, A2 => n170, ZN => n_state_31_port);
   U108 : AND2_X1 port map( A1 => mux_out_25_port, A2 => n172, ZN => 
                           zero_out_25_port);
   U109 : AND2_X1 port map( A1 => mux_out_29_port, A2 => n172, ZN => 
                           zero_out_29_port);
   U110 : AND2_X1 port map( A1 => mux_out_27_port, A2 => n172, ZN => 
                           zero_out_27_port);
   U111 : AND2_X1 port map( A1 => mux_out_26_port, A2 => n172, ZN => 
                           zero_out_26_port);
   U112 : AND2_X1 port map( A1 => mux_out_31_port, A2 => n173, ZN => 
                           zero_out_31_port);
   U113 : AND2_X1 port map( A1 => mux_out_30_port, A2 => n172, ZN => 
                           zero_out_30_port);
   U114 : AND2_X1 port map( A1 => mux_out_24_port, A2 => n172, ZN => 
                           zero_out_24_port);
   U115 : AND2_X1 port map( A1 => mux_out_23_port, A2 => n172, ZN => 
                           zero_out_23_port);
   U116 : AND2_X1 port map( A1 => mux_out_22_port, A2 => n172, ZN => 
                           zero_out_22_port);
   U117 : AND2_X1 port map( A1 => mux_out_28_port, A2 => n172, ZN => 
                           zero_out_28_port);
   U118 : NOR4_X1 port map( A1 => c_state_3_port, A2 => n146, A3 => n148, A4 =>
                           n145, ZN => n91_port);
   U119 : NAND2_X1 port map( A1 => n13_port, A2 => n55_port, ZN => n148);
   U120 : AOI211_X1 port map( C1 => n91_port, C2 => n211, A => n143, B => n144,
                           ZN => n93_port);
   U121 : AOI21_X1 port map( B1 => n13_port, B2 => n55_port, A => n54_port, ZN 
                           => n143);
   U122 : OR2_X1 port map( A1 => n145, A2 => n146, ZN => n144);
   U123 : NAND3_X1 port map( A1 => sign, A2 => n157, A3 => a(15), ZN => n129);
   U124 : NAND2_X1 port map( A1 => n153, A2 => n154, ZN => n146);
   U125 : NOR4_X1 port map( A1 => n156, A2 => c_state_6_port, A3 => 
                           c_state_8_port, A4 => c_state_7_port, ZN => n153);
   U126 : NOR4_X1 port map( A1 => n155, A2 => c_state_25_port, A3 => 
                           c_state_29_port, A4 => c_state_24_port, ZN => n154);
   U127 : AOI22_X1 port map( A1 => en, A2 => lock, B1 => n92_port, B2 => 
                           n53_port, ZN => n77_port);
   U128 : OAI21_X1 port map( B1 => n211, B2 => n54_port, A => n93_port, ZN => 
                           n92_port);
   U129 : OAI21_X1 port map( B1 => n87_port, B2 => n157, A => n129, ZN => N40);
   U130 : OAI21_X1 port map( B1 => n86_port, B2 => n157, A => n129, ZN => N38);
   U131 : OAI21_X1 port map( B1 => n85_port, B2 => n157, A => n129, ZN => N36);
   U132 : OAI21_X1 port map( B1 => n84_port, B2 => n157, A => n129, ZN => N34);
   U133 : OAI21_X1 port map( B1 => n83_port, B2 => n157, A => n129, ZN => N32);
   U134 : OAI21_X1 port map( B1 => n82_port, B2 => n157, A => n129, ZN => N30);
   U135 : OAI21_X1 port map( B1 => n81_port, B2 => n157, A => n129, ZN => N28);
   U136 : OAI21_X1 port map( B1 => n80_port, B2 => n157, A => n129, ZN => N26);
   U137 : OAI21_X1 port map( B1 => n79_port, B2 => n147, A => n129, ZN => N24);
   U138 : OAI21_X1 port map( B1 => n72_port, B2 => n157, A => n129, ZN => N39);
   U139 : OAI21_X1 port map( B1 => n71_port, B2 => n157, A => n129, ZN => N37);
   U140 : OAI21_X1 port map( B1 => n70_port, B2 => n147, A => n129, ZN => N35);
   U141 : OAI21_X1 port map( B1 => n69, B2 => n157, A => n129, ZN => N33);
   U142 : OAI21_X1 port map( B1 => n68, B2 => n157, A => n129, ZN => N31);
   U143 : OAI21_X1 port map( B1 => n67, B2 => n147, A => n129, ZN => N29);
   U144 : OAI21_X1 port map( B1 => n66, B2 => n157, A => n129, ZN => N27);
   U145 : OAI21_X1 port map( B1 => n65, B2 => n157, A => n129, ZN => N25);
   U146 : NAND4_X1 port map( A1 => n24_port, A2 => n23_port, A3 => n22_port, A4
                           => n12_port, ZN => n151);
   U147 : NAND4_X1 port map( A1 => n60, A2 => n59, A3 => n57_port, A4 => 
                           n56_port, ZN => n155);
   U148 : NAND2_X1 port map( A1 => n149, A2 => n150, ZN => n145);
   U149 : NOR4_X1 port map( A1 => n152, A2 => c_state_14_port, A3 => 
                           c_state_16_port, A4 => c_state_15_port, ZN => n149);
   U150 : NOR4_X1 port map( A1 => n151, A2 => c_state_19_port, A3 => 
                           c_state_17_port, A4 => c_state_18_port, ZN => n150);
   U151 : NAND4_X1 port map( A1 => net108738, A2 => net108737, A3 => net108736,
                           A4 => n31_port, ZN => n152);
   U152 : NAND2_X1 port map( A1 => n53_port, A2 => n93_port, ZN => n114);
   U153 : NOR2_X1 port map( A1 => n58, A2 => n157, ZN => N41);
   U154 : INV_X1 port map( A => n113, ZN => n194);
   U155 : AOI22_X1 port map( A1 => adj_sum_0_port, A2 => n97_port, B1 => n161, 
                           B2 => adj_final_mod_15_port, ZN => n113);
   U156 : INV_X1 port map( A => n112, ZN => n195);
   U157 : AOI22_X1 port map( A1 => adj_sum_1_port, A2 => n97_port, B1 => n161, 
                           B2 => adj_final_mod_16_port, ZN => n112);
   U158 : INV_X1 port map( A => n111, ZN => n196);
   U159 : AOI22_X1 port map( A1 => adj_sum_2_port, A2 => n97_port, B1 => n160, 
                           B2 => adj_final_mod_17_port, ZN => n111);
   U160 : INV_X1 port map( A => n110, ZN => n197);
   U161 : AOI22_X1 port map( A1 => adj_sum_3_port, A2 => n97_port, B1 => n161, 
                           B2 => adj_final_mod_18_port, ZN => n110);
   U162 : INV_X1 port map( A => n109, ZN => n198);
   U163 : AOI22_X1 port map( A1 => adj_sum_4_port, A2 => n97_port, B1 => n160, 
                           B2 => adj_final_mod_19_port, ZN => n109);
   U164 : INV_X1 port map( A => n108, ZN => n199);
   U165 : AOI22_X1 port map( A1 => adj_sum_5_port, A2 => n97_port, B1 => n160, 
                           B2 => adj_final_mod_20_port, ZN => n108);
   U166 : INV_X1 port map( A => n107, ZN => n200);
   U167 : AOI22_X1 port map( A1 => adj_sum_6_port, A2 => n97_port, B1 => n159, 
                           B2 => adj_final_mod_21_port, ZN => n107);
   U168 : INV_X1 port map( A => n106, ZN => n201);
   U169 : AOI22_X1 port map( A1 => adj_sum_7_port, A2 => n97_port, B1 => n160, 
                           B2 => adj_final_mod_22_port, ZN => n106);
   U170 : AND2_X1 port map( A1 => a(0), A2 => n157, ZN => N9);
   U171 : INV_X1 port map( A => n121, ZN => N49);
   U172 : AOI22_X1 port map( A1 => b(7), A2 => n157, B1 => n163, B2 => 
                           e_b_10_port, ZN => n121);
   U173 : INV_X1 port map( A => n115, ZN => N55);
   U174 : AOI22_X1 port map( A1 => b(13), A2 => n147, B1 => n161, B2 => 
                           e_b_16_port, ZN => n115);
   U175 : INV_X1 port map( A => n117, ZN => N53);
   U176 : AOI22_X1 port map( A1 => b(11), A2 => n147, B1 => n162, B2 => 
                           e_b_14_port, ZN => n117);
   U177 : INV_X1 port map( A => n119, ZN => N51);
   U178 : AOI22_X1 port map( A1 => b(9), A2 => n147, B1 => n162, B2 => 
                           e_b_12_port, ZN => n119);
   U179 : INV_X1 port map( A => n118, ZN => N52);
   U180 : AOI22_X1 port map( A1 => b(10), A2 => n147, B1 => n162, B2 => 
                           e_b_13_port, ZN => n118);
   U181 : AND2_X1 port map( A1 => a(1), A2 => n157, ZN => N10);
   U182 : INV_X1 port map( A => n125, ZN => N45);
   U183 : AOI22_X1 port map( A1 => b(3), A2 => n147, B1 => n164, B2 => 
                           e_b_6_port, ZN => n125);
   U184 : INV_X1 port map( A => n124, ZN => N46);
   U185 : AOI22_X1 port map( A1 => b(4), A2 => n147, B1 => n164, B2 => 
                           e_b_7_port, ZN => n124);
   U186 : INV_X1 port map( A => n122, ZN => N48);
   U187 : AOI22_X1 port map( A1 => b(6), A2 => n147, B1 => n163, B2 => 
                           e_b_9_port, ZN => n122);
   U188 : INV_X1 port map( A => n116, ZN => N54);
   U189 : AOI22_X1 port map( A1 => b(12), A2 => n147, B1 => n162, B2 => 
                           e_b_15_port, ZN => n116);
   U190 : INV_X1 port map( A => n120, ZN => N50);
   U191 : AOI22_X1 port map( A1 => b(8), A2 => n147, B1 => n163, B2 => 
                           e_b_11_port, ZN => n120);
   U192 : INV_X1 port map( A => n123, ZN => N47);
   U193 : AOI22_X1 port map( A1 => b(5), A2 => n147, B1 => n164, B2 => 
                           e_b_8_port, ZN => n123);
   U194 : INV_X1 port map( A => n131, ZN => N22);
   U195 : AOI22_X1 port map( A1 => a(13), A2 => n147, B1 => n165, B2 => 
                           e_a_11_port, ZN => n131);
   U196 : INV_X1 port map( A => n139, ZN => N14);
   U197 : AOI22_X1 port map( A1 => a(5), A2 => n157, B1 => n167, B2 => 
                           e_a_3_port, ZN => n139);
   U198 : INV_X1 port map( A => n141, ZN => N12);
   U199 : AOI22_X1 port map( A1 => a(3), A2 => n147, B1 => n168, B2 => 
                           e_a_1_port, ZN => n141);
   U200 : INV_X1 port map( A => n133, ZN => N20);
   U201 : AOI22_X1 port map( A1 => a(11), A2 => n157, B1 => n166, B2 => 
                           e_a_9_port, ZN => n133);
   U202 : INV_X1 port map( A => n137, ZN => N16);
   U204 : AOI22_X1 port map( A1 => a(7), A2 => n147, B1 => n167, B2 => 
                           e_a_5_port, ZN => n137);
   U206 : INV_X1 port map( A => n136, ZN => N17);
   U207 : AOI22_X1 port map( A1 => a(8), A2 => n147, B1 => n167, B2 => 
                           e_a_6_port, ZN => n136);
   U208 : INV_X1 port map( A => n128, ZN => N42);
   U209 : AOI22_X1 port map( A1 => b(0), A2 => n157, B1 => n165, B2 => 
                           e_b_3_port, ZN => n128);
   U210 : INV_X1 port map( A => n132, ZN => N21);
   U211 : AOI22_X1 port map( A1 => a(12), A2 => n147, B1 => n166, B2 => 
                           e_a_10_port, ZN => n132);
   U212 : INV_X1 port map( A => n138, ZN => N15);
   U213 : AOI22_X1 port map( A1 => a(6), A2 => n147, B1 => n167, B2 => 
                           e_a_4_port, ZN => n138);
   U214 : INV_X1 port map( A => n130, ZN => N23);
   U215 : AOI22_X1 port map( A1 => a(14), A2 => n157, B1 => n165, B2 => 
                           e_a_12_port, ZN => n130);
   U216 : INV_X1 port map( A => n140, ZN => N13);
   U217 : AOI22_X1 port map( A1 => a(4), A2 => n147, B1 => n168, B2 => 
                           e_a_2_port, ZN => n140);
   U218 : INV_X1 port map( A => n142, ZN => N11);
   U219 : AOI22_X1 port map( A1 => a(2), A2 => n147, B1 => n168, B2 => 
                           e_a_0_port, ZN => n142);
   U220 : INV_X1 port map( A => n127, ZN => N43);
   U221 : AOI22_X1 port map( A1 => b(1), A2 => n147, B1 => n165, B2 => 
                           e_b_4_port, ZN => n127);
   U222 : INV_X1 port map( A => n126, ZN => N44);
   U223 : AOI22_X1 port map( A1 => b(2), A2 => n147, B1 => n164, B2 => 
                           e_b_5_port, ZN => n126);
   U224 : INV_X1 port map( A => n135, ZN => N18);
   U240 : AOI22_X1 port map( A1 => a(9), A2 => n147, B1 => n166, B2 => 
                           e_a_7_port, ZN => n135);
   U241 : INV_X1 port map( A => n134, ZN => N19);
   U242 : AOI22_X1 port map( A1 => a(10), A2 => n147, B1 => n166, B2 => 
                           e_a_8_port, ZN => n134);
   U243 : INV_X1 port map( A => n78_port, ZN => n_state_0_port);
   U244 : AOI21_X1 port map( B1 => n169, B2 => N70, A => n88_port, ZN => 
                           n78_port);
   U245 : AND4_X1 port map( A1 => en, A2 => n53_port, A3 => n89_port, A4 => 
                           n211, ZN => n88_port);

end SYN_booth_mul_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Shifter_DATA_SIZE32 is

   port( l_r, l_a, s_r : in std_logic;  a, b : in std_logic_vector (31 downto 
         0);  o : out std_logic_vector (31 downto 0));

end Shifter_DATA_SIZE32;

architecture SYN_shifter_arch of Shifter_DATA_SIZE32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component Shifter_DATA_SIZE32_DW_rbsh_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component Shifter_DATA_SIZE32_DW_lbsh_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component Shifter_DATA_SIZE32_DW_sra_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component Shifter_DATA_SIZE32_DW_rash_0
      port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH
            : in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out
            std_logic_vector (31 downto 0));
   end component;
   
   component Shifter_DATA_SIZE32_DW_sla_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component Shifter_DATA_SIZE32_DW01_ash_0
      port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH
            : in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out
            std_logic_vector (31 downto 0));
   end component;
   
   signal N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, 
      N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37
      , N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, 
      N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66
      , N67, N68, N69, N70, N71, N72, N108, N109, N110, N111, N112, N113, N114,
      N115, N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, 
      N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, 
      N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, 
      N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, 
      N163, N164, N165, N166, N167, N168, N169, N170, N171, N205, N206, N207, 
      N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, 
      N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, 
      N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, 
      N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, 
      N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, 
      N268, n1, n2, n3, n4, n5, n6, n11_port, n12_port, n13_port, n20_port, 
      n21_port, n22_port, n23_port, n24_port, n25_port, n26_port, n27_port, 
      n28_port, n29_port, n30_port, n31_port, n32_port, n33_port, n34_port, 
      n35_port, n36_port, n37_port, n38_port, n39_port, n40_port, n41_port, 
      n42_port, n43_port, n44_port, n45_port, n46_port, n47_port, n48_port, 
      n49_port, n50_port, n51_port, n52_port, n53_port, n54_port, n55_port, 
      n56_port, n57_port, n58_port, n59_port, n60_port, n61_port, n62_port, 
      n63_port, n64_port, n65_port, n66_port, n67_port, n68_port, n69_port, 
      n70_port, n71_port, n72_port, n73, n74, n75, n76, n77, n78, n79, n80, n81
      , n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, 
      n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, 
      n108_port, n109_port : std_logic;

begin
   
   n1 <= '0';
   n2 <= '0';
   n3 <= '0';
   n4 <= '0';
   n5 <= '0';
   n6 <= '0';
   C93 : Shifter_DATA_SIZE32_DW01_ash_0 port map( A(31) => a(31), A(30) => 
                           a(30), A(29) => a(29), A(28) => a(28), A(27) => 
                           a(27), A(26) => a(26), A(25) => a(25), A(24) => 
                           a(24), A(23) => a(23), A(22) => a(22), A(21) => 
                           a(21), A(20) => a(20), A(19) => a(19), A(18) => 
                           a(18), A(17) => a(17), A(16) => a(16), A(15) => 
                           a(15), A(14) => a(14), A(13) => a(13), A(12) => 
                           a(12), A(11) => a(11), A(10) => a(10), A(9) => a(9),
                           A(8) => a(8), A(7) => a(7), A(6) => a(6), A(5) => 
                           a(5), A(4) => a(4), A(3) => a(3), A(2) => a(2), A(1)
                           => a(1), A(0) => a(0), DATA_TC => n1, SH(4) => 
                           n109_port, SH(3) => n108_port, SH(2) => b(2), SH(1) 
                           => b(1), SH(0) => b(0), SH_TC => n1, B(31) => N268, 
                           B(30) => N267, B(29) => N266, B(28) => N265, B(27) 
                           => N264, B(26) => N263, B(25) => N262, B(24) => N261
                           , B(23) => N260, B(22) => N259, B(21) => N258, B(20)
                           => N257, B(19) => N256, B(18) => N255, B(17) => N254
                           , B(16) => N253, B(15) => N252, B(14) => N251, B(13)
                           => N250, B(12) => N249, B(11) => N248, B(10) => N247
                           , B(9) => N246, B(8) => N245, B(7) => N244, B(6) => 
                           N243, B(5) => N242, B(4) => N241, B(3) => N240, B(2)
                           => N239, B(1) => N238, B(0) => N237);
   C91 : Shifter_DATA_SIZE32_DW_sla_0 port map( A(31) => a(31), A(30) => a(30),
                           A(29) => a(29), A(28) => a(28), A(27) => a(27), 
                           A(26) => a(26), A(25) => a(25), A(24) => a(24), 
                           A(23) => a(23), A(22) => a(22), A(21) => a(21), 
                           A(20) => a(20), A(19) => a(19), A(18) => a(18), 
                           A(17) => a(17), A(16) => a(16), A(15) => a(15), 
                           A(14) => a(14), A(13) => a(13), A(12) => a(12), 
                           A(11) => a(11), A(10) => a(10), A(9) => a(9), A(8) 
                           => a(8), A(7) => a(7), A(6) => a(6), A(5) => a(5), 
                           A(4) => a(4), A(3) => a(3), A(2) => a(2), A(1) => 
                           a(1), A(0) => a(0), SH(4) => n109_port, SH(3) => 
                           n108_port, SH(2) => b(2), SH(1) => b(1), SH(0) => 
                           b(0), SH_TC => n2, B(31) => N236, B(30) => N235, 
                           B(29) => N234, B(28) => N233, B(27) => N232, B(26) 
                           => N231, B(25) => N230, B(24) => N229, B(23) => N228
                           , B(22) => N227, B(21) => N226, B(20) => N225, B(19)
                           => N224, B(18) => N223, B(17) => N222, B(16) => N221
                           , B(15) => N220, B(14) => N219, B(13) => N218, B(12)
                           => N217, B(11) => N216, B(10) => N215, B(9) => N214,
                           B(8) => N213, B(7) => N212, B(6) => N211, B(5) => 
                           N210, B(4) => N209, B(3) => N208, B(2) => N207, B(1)
                           => N206, B(0) => N205);
   C54 : Shifter_DATA_SIZE32_DW_rash_0 port map( A(31) => a(31), A(30) => a(30)
                           , A(29) => a(29), A(28) => a(28), A(27) => a(27), 
                           A(26) => a(26), A(25) => a(25), A(24) => a(24), 
                           A(23) => a(23), A(22) => a(22), A(21) => a(21), 
                           A(20) => a(20), A(19) => a(19), A(18) => a(18), 
                           A(17) => a(17), A(16) => a(16), A(15) => a(15), 
                           A(14) => a(14), A(13) => a(13), A(12) => a(12), 
                           A(11) => a(11), A(10) => a(10), A(9) => a(9), A(8) 
                           => a(8), A(7) => a(7), A(6) => a(6), A(5) => a(5), 
                           A(4) => a(4), A(3) => a(3), A(2) => a(2), A(1) => 
                           a(1), A(0) => a(0), DATA_TC => n3, SH(4) => 
                           n109_port, SH(3) => n108_port, SH(2) => b(2), SH(1) 
                           => b(1), SH(0) => b(0), SH_TC => n3, B(31) => N171, 
                           B(30) => N170, B(29) => N169, B(28) => N168, B(27) 
                           => N167, B(26) => N166, B(25) => N165, B(24) => N164
                           , B(23) => N163, B(22) => N162, B(21) => N161, B(20)
                           => N160, B(19) => N159, B(18) => N158, B(17) => N157
                           , B(16) => N156, B(15) => N155, B(14) => N154, B(13)
                           => N153, B(12) => N152, B(11) => N151, B(10) => N150
                           , B(9) => N149, B(8) => N148, B(7) => N147, B(6) => 
                           N146, B(5) => N145, B(4) => N144, B(3) => N143, B(2)
                           => N142, B(1) => N141, B(0) => N140);
   C52 : Shifter_DATA_SIZE32_DW_sra_0 port map( A(31) => a(31), A(30) => a(30),
                           A(29) => a(29), A(28) => a(28), A(27) => a(27), 
                           A(26) => a(26), A(25) => a(25), A(24) => a(24), 
                           A(23) => a(23), A(22) => a(22), A(21) => a(21), 
                           A(20) => a(20), A(19) => a(19), A(18) => a(18), 
                           A(17) => a(17), A(16) => a(16), A(15) => a(15), 
                           A(14) => a(14), A(13) => a(13), A(12) => a(12), 
                           A(11) => a(11), A(10) => a(10), A(9) => a(9), A(8) 
                           => a(8), A(7) => a(7), A(6) => a(6), A(5) => a(5), 
                           A(4) => a(4), A(3) => a(3), A(2) => a(2), A(1) => 
                           a(1), A(0) => a(0), SH(4) => n109_port, SH(3) => 
                           n108_port, SH(2) => b(2), SH(1) => b(1), SH(0) => 
                           b(0), SH_TC => n4, B(31) => N139, B(30) => N138, 
                           B(29) => N137, B(28) => N136, B(27) => N135, B(26) 
                           => N134, B(25) => N133, B(24) => N132, B(23) => N131
                           , B(22) => N130, B(21) => N129, B(20) => N128, B(19)
                           => N127, B(18) => N126, B(17) => N125, B(16) => N124
                           , B(15) => N123, B(14) => N122, B(13) => N121, B(12)
                           => N120, B(11) => N119, B(10) => N118, B(9) => N117,
                           B(8) => N116, B(7) => N115, B(6) => N114, B(5) => 
                           N113, B(4) => N112, B(3) => N111, B(2) => N110, B(1)
                           => N109, B(0) => N108);
   C12 : Shifter_DATA_SIZE32_DW_lbsh_0 port map( A(31) => a(31), A(30) => a(30)
                           , A(29) => a(29), A(28) => a(28), A(27) => a(27), 
                           A(26) => a(26), A(25) => a(25), A(24) => a(24), 
                           A(23) => a(23), A(22) => a(22), A(21) => a(21), 
                           A(20) => a(20), A(19) => a(19), A(18) => a(18), 
                           A(17) => a(17), A(16) => a(16), A(15) => a(15), 
                           A(14) => a(14), A(13) => a(13), A(12) => a(12), 
                           A(11) => a(11), A(10) => a(10), A(9) => a(9), A(8) 
                           => a(8), A(7) => a(7), A(6) => a(6), A(5) => a(5), 
                           A(4) => a(4), A(3) => a(3), A(2) => a(2), A(1) => 
                           a(1), A(0) => a(0), SH(4) => n109_port, SH(3) => 
                           n108_port, SH(2) => b(2), SH(1) => b(1), SH(0) => 
                           b(0), SH_TC => n5, B(31) => N72, B(30) => N71, B(29)
                           => N70, B(28) => N69, B(27) => N68, B(26) => N67, 
                           B(25) => N66, B(24) => N65, B(23) => N64, B(22) => 
                           N63, B(21) => N62, B(20) => N61, B(19) => N60, B(18)
                           => N59, B(17) => N58, B(16) => N57, B(15) => N56, 
                           B(14) => N55, B(13) => N54, B(12) => N53, B(11) => 
                           N52, B(10) => N51, B(9) => N50, B(8) => N49, B(7) =>
                           N48, B(6) => N47, B(5) => N46, B(4) => N45, B(3) => 
                           N44, B(2) => N43, B(1) => N42, B(0) => N41);
   C10 : Shifter_DATA_SIZE32_DW_rbsh_0 port map( A(31) => a(31), A(30) => a(30)
                           , A(29) => a(29), A(28) => a(28), A(27) => a(27), 
                           A(26) => a(26), A(25) => a(25), A(24) => a(24), 
                           A(23) => a(23), A(22) => a(22), A(21) => a(21), 
                           A(20) => a(20), A(19) => a(19), A(18) => a(18), 
                           A(17) => a(17), A(16) => a(16), A(15) => a(15), 
                           A(14) => a(14), A(13) => a(13), A(12) => a(12), 
                           A(11) => a(11), A(10) => a(10), A(9) => a(9), A(8) 
                           => a(8), A(7) => a(7), A(6) => a(6), A(5) => a(5), 
                           A(4) => a(4), A(3) => a(3), A(2) => a(2), A(1) => 
                           a(1), A(0) => a(0), SH(4) => n109_port, SH(3) => 
                           n108_port, SH(2) => b(2), SH(1) => b(1), SH(0) => 
                           b(0), SH_TC => n6, B(31) => N40, B(30) => N39, B(29)
                           => N38, B(28) => N37, B(27) => N36, B(26) => N35, 
                           B(25) => N34, B(24) => N33, B(23) => N32, B(22) => 
                           N31, B(21) => N30, B(20) => N29, B(19) => N28, B(18)
                           => N27, B(17) => N26, B(16) => N25, B(15) => N24, 
                           B(14) => N23, B(13) => N22, B(12) => N21, B(11) => 
                           N20, B(10) => N19, B(9) => N18, B(8) => N17, B(7) =>
                           N16, B(6) => N15, B(5) => N14, B(4) => N13, B(3) => 
                           N12, B(2) => N11, B(1) => N10, B(0) => N9);
   U1 : CLKBUF_X1 port map( A => b(3), Z => n108_port);
   U2 : NAND2_X1 port map( A1 => n43_port, A2 => n44_port, ZN => o(29));
   U3 : AOI222_X1 port map( A1 => N38, A2 => n97, B1 => N137, B2 => n94, C1 => 
                           N70, C2 => n91, ZN => n43_port);
   U4 : AOI222_X1 port map( A1 => N234, A2 => n106, B1 => N266, B2 => n103, C1 
                           => N169, C2 => n100, ZN => n44_port);
   U11 : NAND2_X1 port map( A1 => n47_port, A2 => n48_port, ZN => o(27));
   U12 : AOI222_X1 port map( A1 => N36, A2 => n97, B1 => N135, B2 => n94, C1 =>
                           N68, C2 => n91, ZN => n47_port);
   U13 : AOI222_X1 port map( A1 => N232, A2 => n106, B1 => N264, B2 => n103, C1
                           => N167, C2 => n100, ZN => n48_port);
   U14 : NAND2_X1 port map( A1 => n49_port, A2 => n50_port, ZN => o(26));
   U15 : AOI222_X1 port map( A1 => N35, A2 => n97, B1 => N134, B2 => n94, C1 =>
                           N67, C2 => n91, ZN => n49_port);
   U16 : AOI222_X1 port map( A1 => N231, A2 => n106, B1 => N263, B2 => n103, C1
                           => N166, C2 => n100, ZN => n50_port);
   U17 : NAND2_X1 port map( A1 => n51_port, A2 => n52_port, ZN => o(25));
   U18 : AOI222_X1 port map( A1 => N34, A2 => n97, B1 => N133, B2 => n94, C1 =>
                           N66, C2 => n91, ZN => n51_port);
   U19 : AOI222_X1 port map( A1 => N230, A2 => n106, B1 => N262, B2 => n103, C1
                           => N165, C2 => n100, ZN => n52_port);
   U20 : NAND2_X1 port map( A1 => n59_port, A2 => n60_port, ZN => o(21));
   U21 : AOI222_X1 port map( A1 => N30, A2 => n97, B1 => N129, B2 => n94, C1 =>
                           N62, C2 => n91, ZN => n59_port);
   U22 : AOI222_X1 port map( A1 => N226, A2 => n106, B1 => N258, B2 => n103, C1
                           => N161, C2 => n100, ZN => n60_port);
   U23 : NAND2_X1 port map( A1 => n57_port, A2 => n58_port, ZN => o(22));
   U24 : AOI222_X1 port map( A1 => N31, A2 => n97, B1 => N130, B2 => n94, C1 =>
                           N63, C2 => n91, ZN => n57_port);
   U25 : AOI222_X1 port map( A1 => N227, A2 => n106, B1 => N259, B2 => n103, C1
                           => N162, C2 => n100, ZN => n58_port);
   U26 : NAND2_X1 port map( A1 => n55_port, A2 => n56_port, ZN => o(23));
   U27 : AOI222_X1 port map( A1 => N32, A2 => n97, B1 => N131, B2 => n94, C1 =>
                           N64, C2 => n91, ZN => n55_port);
   U28 : AOI222_X1 port map( A1 => N228, A2 => n106, B1 => N260, B2 => n103, C1
                           => N163, C2 => n100, ZN => n56_port);
   U29 : NAND2_X1 port map( A1 => n77, A2 => n78, ZN => o(13));
   U30 : AOI222_X1 port map( A1 => N22, A2 => n96, B1 => N121, B2 => n93, C1 =>
                           N54, C2 => n90, ZN => n77);
   U31 : AOI222_X1 port map( A1 => N218, A2 => n105, B1 => N250, B2 => n102, C1
                           => N153, C2 => n99, ZN => n78);
   U32 : NAND2_X1 port map( A1 => n75, A2 => n76, ZN => o(14));
   U33 : AOI222_X1 port map( A1 => N23, A2 => n96, B1 => N122, B2 => n93, C1 =>
                           N55, C2 => n90, ZN => n75);
   U34 : AOI222_X1 port map( A1 => N219, A2 => n105, B1 => N251, B2 => n102, C1
                           => N154, C2 => n99, ZN => n76);
   U35 : NAND2_X1 port map( A1 => n73, A2 => n74, ZN => o(15));
   U36 : AOI222_X1 port map( A1 => N24, A2 => n96, B1 => N123, B2 => n93, C1 =>
                           N56, C2 => n90, ZN => n73);
   U37 : AOI222_X1 port map( A1 => N220, A2 => n105, B1 => N252, B2 => n102, C1
                           => N155, C2 => n99, ZN => n74);
   U38 : NAND2_X1 port map( A1 => n69_port, A2 => n70_port, ZN => o(17));
   U39 : AOI222_X1 port map( A1 => N222, A2 => n105, B1 => N254, B2 => n102, C1
                           => N157, C2 => n99, ZN => n70_port);
   U40 : AOI222_X1 port map( A1 => N26, A2 => n96, B1 => N125, B2 => n93, C1 =>
                           N58, C2 => n90, ZN => n69_port);
   U41 : NAND2_X1 port map( A1 => n67_port, A2 => n68_port, ZN => o(18));
   U42 : AOI222_X1 port map( A1 => N223, A2 => n105, B1 => N255, B2 => n102, C1
                           => N158, C2 => n99, ZN => n68_port);
   U43 : AOI222_X1 port map( A1 => N27, A2 => n96, B1 => N126, B2 => n93, C1 =>
                           N59, C2 => n90, ZN => n67_port);
   U44 : NAND2_X1 port map( A1 => n65_port, A2 => n66_port, ZN => o(19));
   U45 : AOI222_X1 port map( A1 => N224, A2 => n105, B1 => N256, B2 => n102, C1
                           => N159, C2 => n99, ZN => n66_port);
   U46 : AOI222_X1 port map( A1 => N28, A2 => n96, B1 => N127, B2 => n93, C1 =>
                           N60, C2 => n90, ZN => n65_port);
   U47 : NAND2_X1 port map( A1 => n35_port, A2 => n36_port, ZN => o(3));
   U48 : AOI222_X1 port map( A1 => N12, A2 => n98, B1 => N111, B2 => n95, C1 =>
                           N44, C2 => n92, ZN => n35_port);
   U49 : AOI222_X1 port map( A1 => N208, A2 => n107, B1 => N240, B2 => n104, C1
                           => N143, C2 => n101, ZN => n36_port);
   U50 : NAND2_X1 port map( A1 => n33_port, A2 => n34_port, ZN => o(4));
   U51 : AOI222_X1 port map( A1 => N209, A2 => n107, B1 => N241, B2 => n104, C1
                           => N144, C2 => n101, ZN => n34_port);
   U52 : AOI222_X1 port map( A1 => N13, A2 => n98, B1 => N112, B2 => n95, C1 =>
                           N45, C2 => n92, ZN => n33_port);
   U53 : NAND2_X1 port map( A1 => n31_port, A2 => n32_port, ZN => o(5));
   U54 : AOI222_X1 port map( A1 => N14, A2 => n98, B1 => N113, B2 => n95, C1 =>
                           N46, C2 => n92, ZN => n31_port);
   U55 : AOI222_X1 port map( A1 => N210, A2 => n107, B1 => N242, B2 => n104, C1
                           => N145, C2 => n101, ZN => n32_port);
   U56 : NAND2_X1 port map( A1 => n29_port, A2 => n30_port, ZN => o(6));
   U57 : AOI222_X1 port map( A1 => N211, A2 => n107, B1 => N243, B2 => n104, C1
                           => N146, C2 => n101, ZN => n30_port);
   U58 : AOI222_X1 port map( A1 => N15, A2 => n98, B1 => N114, B2 => n95, C1 =>
                           N47, C2 => n92, ZN => n29_port);
   U59 : NAND2_X1 port map( A1 => n27_port, A2 => n28_port, ZN => o(7));
   U60 : AOI222_X1 port map( A1 => N16, A2 => n98, B1 => N115, B2 => n95, C1 =>
                           N48, C2 => n92, ZN => n27_port);
   U61 : AOI222_X1 port map( A1 => N212, A2 => n107, B1 => N244, B2 => n104, C1
                           => N147, C2 => n101, ZN => n28_port);
   U62 : NAND2_X1 port map( A1 => n25_port, A2 => n26_port, ZN => o(8));
   U63 : AOI222_X1 port map( A1 => N213, A2 => n107, B1 => N245, B2 => n104, C1
                           => N148, C2 => n101, ZN => n26_port);
   U64 : AOI222_X1 port map( A1 => N17, A2 => n98, B1 => N116, B2 => n95, C1 =>
                           N49, C2 => n92, ZN => n25_port);
   U65 : NAND2_X1 port map( A1 => n11_port, A2 => n12_port, ZN => o(9));
   U66 : AOI222_X1 port map( A1 => N214, A2 => n107, B1 => N246, B2 => n104, C1
                           => N149, C2 => n101, ZN => n12_port);
   U67 : AOI222_X1 port map( A1 => N18, A2 => n98, B1 => N117, B2 => n95, C1 =>
                           N50, C2 => n92, ZN => n11_port);
   U68 : NAND2_X1 port map( A1 => n85, A2 => n86, ZN => o(0));
   U69 : AOI222_X1 port map( A1 => N205, A2 => n105, B1 => N237, B2 => n102, C1
                           => N140, C2 => n99, ZN => n86);
   U70 : AOI222_X1 port map( A1 => N9, A2 => n96, B1 => N108, B2 => n93, C1 => 
                           N41, C2 => n90, ZN => n85);
   U71 : NAND2_X1 port map( A1 => n63_port, A2 => n64_port, ZN => o(1));
   U72 : AOI222_X1 port map( A1 => N206, A2 => n105, B1 => N238, B2 => n102, C1
                           => N141, C2 => n99, ZN => n64_port);
   U73 : AOI222_X1 port map( A1 => N10, A2 => n96, B1 => N109, B2 => n93, C1 =>
                           N42, C2 => n90, ZN => n63_port);
   U74 : NAND2_X1 port map( A1 => n41_port, A2 => n42_port, ZN => o(2));
   U75 : AOI222_X1 port map( A1 => N207, A2 => n106, B1 => N239, B2 => n103, C1
                           => N142, C2 => n100, ZN => n42_port);
   U76 : AOI222_X1 port map( A1 => N11, A2 => n97, B1 => N110, B2 => n94, C1 =>
                           N43, C2 => n91, ZN => n41_port);
   U77 : NAND2_X1 port map( A1 => n83, A2 => n84, ZN => o(10));
   U78 : AOI222_X1 port map( A1 => N215, A2 => n105, B1 => N247, B2 => n102, C1
                           => N150, C2 => n99, ZN => n84);
   U79 : AOI222_X1 port map( A1 => N19, A2 => n96, B1 => N118, B2 => n93, C1 =>
                           N51, C2 => n90, ZN => n83);
   U80 : NAND2_X1 port map( A1 => n81, A2 => n82, ZN => o(11));
   U81 : AOI222_X1 port map( A1 => N20, A2 => n96, B1 => N119, B2 => n93, C1 =>
                           N52, C2 => n90, ZN => n81);
   U82 : AOI222_X1 port map( A1 => N216, A2 => n105, B1 => N248, B2 => n102, C1
                           => N151, C2 => n99, ZN => n82);
   U83 : BUF_X1 port map( A => n22_port, Z => n96);
   U84 : BUF_X1 port map( A => n22_port, Z => n97);
   U85 : BUF_X1 port map( A => n22_port, Z => n98);
   U86 : NAND2_X1 port map( A1 => n37_port, A2 => n38_port, ZN => o(31));
   U87 : AOI222_X1 port map( A1 => N40, A2 => n98, B1 => N139, B2 => n95, C1 =>
                           N72, C2 => n92, ZN => n37_port);
   U88 : AOI222_X1 port map( A1 => N236, A2 => n107, B1 => N268, B2 => n104, C1
                           => N171, C2 => n101, ZN => n38_port);
   U89 : NAND2_X1 port map( A1 => n45_port, A2 => n46_port, ZN => o(28));
   U90 : AOI222_X1 port map( A1 => N37, A2 => n97, B1 => N136, B2 => n94, C1 =>
                           N69, C2 => n91, ZN => n45_port);
   U91 : AOI222_X1 port map( A1 => N233, A2 => n106, B1 => N265, B2 => n103, C1
                           => N168, C2 => n100, ZN => n46_port);
   U92 : NAND2_X1 port map( A1 => n39_port, A2 => n40_port, ZN => o(30));
   U93 : AOI222_X1 port map( A1 => N39, A2 => n97, B1 => N138, B2 => n94, C1 =>
                           N71, C2 => n91, ZN => n39_port);
   U94 : AOI222_X1 port map( A1 => N235, A2 => n106, B1 => N267, B2 => n103, C1
                           => N170, C2 => n100, ZN => n40_port);
   U95 : NAND2_X1 port map( A1 => n53_port, A2 => n54_port, ZN => o(24));
   U96 : AOI222_X1 port map( A1 => N33, A2 => n97, B1 => N132, B2 => n94, C1 =>
                           N65, C2 => n91, ZN => n53_port);
   U97 : AOI222_X1 port map( A1 => N229, A2 => n106, B1 => N261, B2 => n103, C1
                           => N164, C2 => n100, ZN => n54_port);
   U98 : NAND2_X1 port map( A1 => n61_port, A2 => n62_port, ZN => o(20));
   U99 : AOI222_X1 port map( A1 => N225, A2 => n106, B1 => N257, B2 => n103, C1
                           => N160, C2 => n100, ZN => n62_port);
   U100 : AOI222_X1 port map( A1 => N29, A2 => n97, B1 => N128, B2 => n94, C1 
                           => N61, C2 => n91, ZN => n61_port);
   U101 : NAND2_X1 port map( A1 => n79, A2 => n80, ZN => o(12));
   U102 : AOI222_X1 port map( A1 => N21, A2 => n96, B1 => N120, B2 => n93, C1 
                           => N53, C2 => n90, ZN => n79);
   U103 : AOI222_X1 port map( A1 => N217, A2 => n105, B1 => N249, B2 => n102, 
                           C1 => N152, C2 => n99, ZN => n80);
   U104 : NAND2_X1 port map( A1 => n71_port, A2 => n72_port, ZN => o(16));
   U105 : AOI222_X1 port map( A1 => N221, A2 => n105, B1 => N253, B2 => n102, 
                           C1 => N156, C2 => n99, ZN => n72_port);
   U106 : AOI222_X1 port map( A1 => N25, A2 => n96, B1 => N124, B2 => n93, C1 
                           => N57, C2 => n90, ZN => n71_port);
   U107 : BUF_X1 port map( A => n13_port, Z => n105);
   U108 : BUF_X1 port map( A => n13_port, Z => n106);
   U109 : BUF_X1 port map( A => n20_port, Z => n102);
   U110 : BUF_X1 port map( A => n20_port, Z => n103);
   U111 : BUF_X1 port map( A => n23_port, Z => n93);
   U112 : BUF_X1 port map( A => n23_port, Z => n94);
   U113 : NOR2_X1 port map( A1 => n89, A2 => n87, ZN => n22_port);
   U114 : BUF_X1 port map( A => n21_port, Z => n99);
   U115 : BUF_X1 port map( A => n21_port, Z => n100);
   U116 : BUF_X1 port map( A => n24_port, Z => n90);
   U117 : BUF_X1 port map( A => n24_port, Z => n91);
   U118 : BUF_X1 port map( A => n20_port, Z => n104);
   U119 : BUF_X1 port map( A => n21_port, Z => n101);
   U120 : BUF_X1 port map( A => n23_port, Z => n95);
   U121 : BUF_X1 port map( A => n24_port, Z => n92);
   U122 : CLKBUF_X1 port map( A => b(4), Z => n109_port);
   U123 : BUF_X1 port map( A => n13_port, Z => n107);
   U124 : NOR3_X1 port map( A1 => n87, A2 => s_r, A3 => n88, ZN => n23_port);
   U125 : NOR3_X1 port map( A1 => l_r, A2 => s_r, A3 => n88, ZN => n13_port);
   U126 : NOR2_X1 port map( A1 => n89, A2 => l_r, ZN => n24_port);
   U127 : INV_X1 port map( A => l_r, ZN => n87);
   U128 : INV_X1 port map( A => s_r, ZN => n89);
   U129 : NOR3_X1 port map( A1 => l_r, A2 => s_r, A3 => l_a, ZN => n20_port);
   U130 : NOR3_X1 port map( A1 => l_a, A2 => s_r, A3 => n87, ZN => n21_port);
   U131 : INV_X1 port map( A => l_a, ZN => n88);

end SYN_shifter_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4Adder_DATA_SIZE32_SPARSITY4_0 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end P4Adder_DATA_SIZE32_SPARSITY4_0;

architecture SYN_p4_adder_arch of P4Adder_DATA_SIZE32_SPARSITY4_0 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AdderSumGenerator_DATA_SIZE32_SPARSITY4_0
      port( a, b : in std_logic_vector (31 downto 0);  cin : in 
            std_logic_vector (7 downto 0);  sum : out std_logic_vector (31 
            downto 0));
   end component;
   
   component P4CarryGenerator_DATA_SIZE32_SPARSITY4_0
      port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  
            cout : out std_logic_vector (7 downto 0));
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, carry_1_port, n1, n2, n3 : std_logic;

begin
   
   CG0 : P4CarryGenerator_DATA_SIZE32_SPARSITY4_0 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => n2, a(27) 
                           => a(27), a(26) => a(26), a(25) => a(25), a(24) => 
                           a(24), a(23) => a(23), a(22) => a(22), a(21) => 
                           a(21), a(20) => a(20), a(19) => a(19), a(18) => 
                           a(18), a(17) => a(17), a(16) => a(16), a(15) => 
                           a(15), a(14) => a(14), a(13) => a(13), a(12) => 
                           a(12), a(11) => a(11), a(10) => a(10), a(9) => a(9),
                           a(8) => a(8), a(7) => a(7), a(6) => a(6), a(5) => 
                           a(5), a(4) => a(4), a(3) => a(3), a(2) => a(2), a(1)
                           => a(1), a(0) => a(0), b(31) => b(31), b(30) => 
                           b(30), b(29) => b(29), b(28) => b(28), b(27) => 
                           b(27), b(26) => b(26), b(25) => b(25), b(24) => 
                           b(24), b(23) => b(23), b(22) => b(22), b(21) => 
                           b(21), b(20) => b(20), b(19) => b(19), b(18) => 
                           b(18), b(17) => b(17), b(16) => b(16), b(15) => 
                           b(15), b(14) => b(14), b(13) => b(13), b(12) => 
                           b(12), b(11) => b(11), b(10) => b(10), b(9) => b(9),
                           b(8) => b(8), b(7) => b(7), b(6) => b(6), b(5) => 
                           b(5), b(4) => b(4), b(3) => b(3), b(2) => b(2), b(1)
                           => b(1), b(0) => b(0), cin => cin, cout(7) => cout, 
                           cout(6) => carry_7_port, cout(5) => carry_6_port, 
                           cout(4) => carry_5_port, cout(3) => carry_4_port, 
                           cout(2) => carry_3_port, cout(1) => carry_2_port, 
                           cout(0) => carry_1_port);
   SG0 : AdderSumGenerator_DATA_SIZE32_SPARSITY4_0 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => n1, a(0) => n3, b(31) => b(31), b(30) 
                           => b(30), b(29) => b(29), b(28) => b(28), b(27) => 
                           b(27), b(26) => b(26), b(25) => b(25), b(24) => 
                           b(24), b(23) => b(23), b(22) => b(22), b(21) => 
                           b(21), b(20) => b(20), b(19) => b(19), b(18) => 
                           b(18), b(17) => b(17), b(16) => b(16), b(15) => 
                           b(15), b(14) => b(14), b(13) => b(13), b(12) => 
                           b(12), b(11) => b(11), b(10) => b(10), b(9) => b(9),
                           b(8) => b(8), b(7) => b(7), b(6) => b(6), b(5) => 
                           b(5), b(4) => b(4), b(3) => b(3), b(2) => b(2), b(1)
                           => b(1), b(0) => b(0), cin(7) => carry_7_port, 
                           cin(6) => carry_6_port, cin(5) => carry_5_port, 
                           cin(4) => carry_4_port, cin(3) => carry_3_port, 
                           cin(2) => carry_2_port, cin(1) => carry_1_port, 
                           cin(0) => cin, sum(31) => s(31), sum(30) => s(30), 
                           sum(29) => s(29), sum(28) => s(28), sum(27) => s(27)
                           , sum(26) => s(26), sum(25) => s(25), sum(24) => 
                           s(24), sum(23) => s(23), sum(22) => s(22), sum(21) 
                           => s(21), sum(20) => s(20), sum(19) => s(19), 
                           sum(18) => s(18), sum(17) => s(17), sum(16) => s(16)
                           , sum(15) => s(15), sum(14) => s(14), sum(13) => 
                           s(13), sum(12) => s(12), sum(11) => s(11), sum(10) 
                           => s(10), sum(9) => s(9), sum(8) => s(8), sum(7) => 
                           s(7), sum(6) => s(6), sum(5) => s(5), sum(4) => s(4)
                           , sum(3) => s(3), sum(2) => s(2), sum(1) => s(1), 
                           sum(0) => s(0));
   U1 : CLKBUF_X1 port map( A => a(1), Z => n1);
   U2 : CLKBUF_X1 port map( A => a(28), Z => n2);
   U3 : CLKBUF_X1 port map( A => a(0), Z => n3);

end SYN_p4_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity StallGenerator_CWRD_SIZE20_DW01_inc_5 is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end StallGenerator_CWRD_SIZE20_DW01_inc_5;

architecture SYN_rpl of StallGenerator_CWRD_SIZE20_DW01_inc_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port : std_logic;

begin
   
   U1_1_30 : HA_X1 port map( A => A(30), B => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_1_29 : HA_X1 port map( A => A(29), B => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_1_28 : HA_X1 port map( A => A(28), B => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_1_27 : HA_X1 port map( A => A(27), B => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_1_26 : HA_X1 port map( A => A(26), B => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_1_25 : HA_X1 port map( A => A(25), B => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_1_24 : HA_X1 port map( A => A(24), B => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_1_23 : HA_X1 port map( A => A(23), B => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_1_22 : HA_X1 port map( A => A(22), B => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_1_21 : HA_X1 port map( A => A(21), B => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_1_20 : HA_X1 port map( A => A(20), B => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_1_19 : HA_X1 port map( A => A(19), B => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_1_18 : HA_X1 port map( A => A(18), B => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_1_17 : HA_X1 port map( A => A(17), B => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_1_16 : HA_X1 port map( A => A(16), B => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_1_15 : HA_X1 port map( A => A(15), B => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : XOR2_X1 port map( A => carry_31_port, B => A(31), Z => SUM(31));
   U2 : INV_X1 port map( A => A(0), ZN => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity StallGenerator_CWRD_SIZE20_DW01_inc_4 is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end StallGenerator_CWRD_SIZE20_DW01_inc_4;

architecture SYN_rpl of StallGenerator_CWRD_SIZE20_DW01_inc_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port : std_logic;

begin
   
   U1_1_30 : HA_X1 port map( A => A(30), B => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_1_29 : HA_X1 port map( A => A(29), B => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_1_28 : HA_X1 port map( A => A(28), B => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_1_27 : HA_X1 port map( A => A(27), B => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_1_26 : HA_X1 port map( A => A(26), B => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_1_25 : HA_X1 port map( A => A(25), B => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_1_24 : HA_X1 port map( A => A(24), B => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_1_23 : HA_X1 port map( A => A(23), B => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_1_22 : HA_X1 port map( A => A(22), B => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_1_21 : HA_X1 port map( A => A(21), B => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_1_20 : HA_X1 port map( A => A(20), B => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_1_19 : HA_X1 port map( A => A(19), B => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_1_18 : HA_X1 port map( A => A(18), B => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_1_17 : HA_X1 port map( A => A(17), B => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_1_16 : HA_X1 port map( A => A(16), B => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_1_15 : HA_X1 port map( A => A(15), B => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : XOR2_X1 port map( A => carry_31_port, B => A(31), Z => SUM(31));
   U2 : INV_X1 port map( A => A(0), ZN => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity StallGenerator_CWRD_SIZE20_DW01_inc_3 is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end StallGenerator_CWRD_SIZE20_DW01_inc_3;

architecture SYN_rpl of StallGenerator_CWRD_SIZE20_DW01_inc_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port : std_logic;

begin
   
   U1_1_30 : HA_X1 port map( A => A(30), B => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_1_29 : HA_X1 port map( A => A(29), B => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_1_28 : HA_X1 port map( A => A(28), B => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_1_27 : HA_X1 port map( A => A(27), B => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_1_26 : HA_X1 port map( A => A(26), B => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_1_25 : HA_X1 port map( A => A(25), B => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_1_24 : HA_X1 port map( A => A(24), B => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_1_23 : HA_X1 port map( A => A(23), B => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_1_22 : HA_X1 port map( A => A(22), B => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_1_21 : HA_X1 port map( A => A(21), B => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_1_20 : HA_X1 port map( A => A(20), B => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_1_19 : HA_X1 port map( A => A(19), B => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_1_18 : HA_X1 port map( A => A(18), B => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_1_17 : HA_X1 port map( A => A(17), B => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_1_16 : HA_X1 port map( A => A(16), B => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_1_15 : HA_X1 port map( A => A(15), B => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : XOR2_X1 port map( A => carry_31_port, B => A(31), Z => SUM(31));
   U2 : INV_X1 port map( A => A(0), ZN => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity StallGenerator_CWRD_SIZE20_DW01_inc_2 is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end StallGenerator_CWRD_SIZE20_DW01_inc_2;

architecture SYN_rpl of StallGenerator_CWRD_SIZE20_DW01_inc_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port : std_logic;

begin
   
   U1_1_30 : HA_X1 port map( A => A(30), B => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_1_29 : HA_X1 port map( A => A(29), B => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_1_28 : HA_X1 port map( A => A(28), B => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_1_27 : HA_X1 port map( A => A(27), B => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_1_26 : HA_X1 port map( A => A(26), B => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_1_25 : HA_X1 port map( A => A(25), B => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_1_24 : HA_X1 port map( A => A(24), B => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_1_23 : HA_X1 port map( A => A(23), B => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_1_22 : HA_X1 port map( A => A(22), B => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_1_21 : HA_X1 port map( A => A(21), B => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_1_20 : HA_X1 port map( A => A(20), B => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_1_19 : HA_X1 port map( A => A(19), B => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_1_18 : HA_X1 port map( A => A(18), B => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_1_17 : HA_X1 port map( A => A(17), B => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_1_16 : HA_X1 port map( A => A(16), B => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_1_15 : HA_X1 port map( A => A(15), B => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : XOR2_X1 port map( A => carry_31_port, B => A(31), Z => SUM(31));
   U2 : INV_X1 port map( A => A(0), ZN => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity StallGenerator_CWRD_SIZE20_DW01_inc_1 is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end StallGenerator_CWRD_SIZE20_DW01_inc_1;

architecture SYN_rpl of StallGenerator_CWRD_SIZE20_DW01_inc_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port : std_logic;

begin
   
   U1_1_30 : HA_X1 port map( A => A(30), B => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_1_29 : HA_X1 port map( A => A(29), B => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_1_28 : HA_X1 port map( A => A(28), B => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_1_27 : HA_X1 port map( A => A(27), B => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_1_26 : HA_X1 port map( A => A(26), B => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_1_25 : HA_X1 port map( A => A(25), B => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_1_24 : HA_X1 port map( A => A(24), B => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_1_23 : HA_X1 port map( A => A(23), B => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_1_22 : HA_X1 port map( A => A(22), B => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_1_21 : HA_X1 port map( A => A(21), B => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_1_20 : HA_X1 port map( A => A(20), B => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_1_19 : HA_X1 port map( A => A(19), B => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_1_18 : HA_X1 port map( A => A(18), B => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_1_17 : HA_X1 port map( A => A(17), B => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_1_16 : HA_X1 port map( A => A(16), B => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_1_15 : HA_X1 port map( A => A(15), B => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : XOR2_X1 port map( A => carry_31_port, B => A(31), Z => SUM(31));
   U2 : INV_X1 port map( A => A(0), ZN => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity StallGenerator_CWRD_SIZE20_DW01_inc_0 is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end StallGenerator_CWRD_SIZE20_DW01_inc_0;

architecture SYN_rpl of StallGenerator_CWRD_SIZE20_DW01_inc_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port : std_logic;

begin
   
   U1_1_30 : HA_X1 port map( A => A(30), B => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_1_29 : HA_X1 port map( A => A(29), B => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_1_28 : HA_X1 port map( A => A(28), B => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_1_27 : HA_X1 port map( A => A(27), B => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_1_26 : HA_X1 port map( A => A(26), B => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_1_25 : HA_X1 port map( A => A(25), B => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_1_24 : HA_X1 port map( A => A(24), B => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_1_23 : HA_X1 port map( A => A(23), B => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_1_22 : HA_X1 port map( A => A(22), B => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_1_21 : HA_X1 port map( A => A(21), B => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_1_20 : HA_X1 port map( A => A(20), B => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_1_19 : HA_X1 port map( A => A(19), B => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_1_18 : HA_X1 port map( A => A(18), B => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_1_17 : HA_X1 port map( A => A(17), B => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_1_16 : HA_X1 port map( A => A(16), B => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_1_15 : HA_X1 port map( A => A(15), B => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : XOR2_X1 port map( A => carry_31_port, B => A(31), Z => SUM(31));
   U2 : INV_X1 port map( A => A(0), ZN => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE32_3 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 0);
         dout : out std_logic_vector (31 downto 0));

end Reg_DATA_SIZE32_3;

architecture SYN_reg_arch of Reg_DATA_SIZE32_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99 : std_logic;

begin
   
   dout_reg_1_inst : DFFR_X1 port map( D => n63, CK => clk, RN => n97, Q => 
                           dout(1), QN => n31);
   dout_reg_2_inst : DFFR_X1 port map( D => n62, CK => clk, RN => n97, Q => 
                           dout(2), QN => n30);
   dout_reg_3_inst : DFFR_X1 port map( D => n61, CK => clk, RN => n97, Q => 
                           dout(3), QN => n29);
   dout_reg_4_inst : DFFR_X1 port map( D => n60, CK => clk, RN => n98, Q => 
                           dout(4), QN => n28);
   dout_reg_5_inst : DFFR_X1 port map( D => n59, CK => clk, RN => n98, Q => 
                           dout(5), QN => n27);
   dout_reg_6_inst : DFFR_X1 port map( D => n58, CK => clk, RN => n97, Q => 
                           dout(6), QN => n26);
   dout_reg_7_inst : DFFR_X1 port map( D => n57, CK => clk, RN => n98, Q => 
                           dout(7), QN => n25);
   dout_reg_8_inst : DFFR_X1 port map( D => n56, CK => clk, RN => n98, Q => 
                           dout(8), QN => n24);
   dout_reg_9_inst : DFFR_X1 port map( D => n55, CK => clk, RN => n99, Q => 
                           dout(9), QN => n23);
   dout_reg_10_inst : DFFR_X1 port map( D => n54, CK => clk, RN => n97, Q => 
                           dout(10), QN => n22);
   dout_reg_11_inst : DFFR_X1 port map( D => n53, CK => clk, RN => n97, Q => 
                           dout(11), QN => n21);
   dout_reg_12_inst : DFFR_X1 port map( D => n52, CK => clk, RN => n97, Q => 
                           dout(12), QN => n20);
   dout_reg_13_inst : DFFR_X1 port map( D => n51, CK => clk, RN => n97, Q => 
                           dout(13), QN => n19);
   dout_reg_14_inst : DFFR_X1 port map( D => n50, CK => clk, RN => n97, Q => 
                           dout(14), QN => n18);
   dout_reg_15_inst : DFFR_X1 port map( D => n49, CK => clk, RN => n98, Q => 
                           dout(15), QN => n17);
   dout_reg_16_inst : DFFR_X1 port map( D => n48, CK => clk, RN => n97, Q => 
                           dout(16), QN => n16);
   dout_reg_17_inst : DFFR_X1 port map( D => n47, CK => clk, RN => n97, Q => 
                           dout(17), QN => n15);
   dout_reg_18_inst : DFFR_X1 port map( D => n46, CK => clk, RN => n98, Q => 
                           dout(18), QN => n14);
   dout_reg_19_inst : DFFR_X1 port map( D => n45, CK => clk, RN => n97, Q => 
                           dout(19), QN => n13);
   dout_reg_20_inst : DFFR_X1 port map( D => n44, CK => clk, RN => n98, Q => 
                           dout(20), QN => n12);
   dout_reg_21_inst : DFFR_X1 port map( D => n43, CK => clk, RN => n98, Q => 
                           dout(21), QN => n11);
   dout_reg_22_inst : DFFR_X1 port map( D => n42, CK => clk, RN => n98, Q => 
                           dout(22), QN => n10);
   dout_reg_24_inst : DFFR_X1 port map( D => n40, CK => clk, RN => n99, Q => 
                           dout(24), QN => n8);
   dout_reg_25_inst : DFFR_X1 port map( D => n39, CK => clk, RN => n98, Q => 
                           dout(25), QN => n7);
   dout_reg_26_inst : DFFR_X1 port map( D => n38, CK => clk, RN => n98, Q => 
                           dout(26), QN => n6);
   dout_reg_27_inst : DFFR_X1 port map( D => n37, CK => clk, RN => n99, Q => 
                           dout(27), QN => n5);
   dout_reg_28_inst : DFFR_X1 port map( D => n36, CK => clk, RN => n99, Q => 
                           dout(28), QN => n4);
   dout_reg_29_inst : DFFR_X1 port map( D => n35, CK => clk, RN => n99, Q => 
                           dout(29), QN => n3);
   dout_reg_30_inst : DFFR_X1 port map( D => n34, CK => clk, RN => n99, Q => 
                           dout(30), QN => n2);
   dout_reg_31_inst : DFFR_X1 port map( D => n33, CK => clk, RN => n99, Q => 
                           dout(31), QN => n1);
   dout_reg_23_inst : DFFR_X1 port map( D => n41, CK => clk, RN => n98, Q => 
                           dout(23), QN => n9);
   dout_reg_0_inst : DFFR_X1 port map( D => n64, CK => clk, RN => n99, Q => 
                           dout(0), QN => n32);
   U2 : BUF_X1 port map( A => rst, Z => n98);
   U3 : BUF_X1 port map( A => rst, Z => n97);
   U4 : BUF_X1 port map( A => rst, Z => n99);
   U5 : OAI21_X1 port map( B1 => n1, B2 => en, A => n96, ZN => n33);
   U6 : NAND2_X1 port map( A1 => din(31), A2 => en, ZN => n96);
   U7 : OAI21_X1 port map( B1 => n2, B2 => en, A => n95, ZN => n34);
   U8 : NAND2_X1 port map( A1 => din(30), A2 => en, ZN => n95);
   U9 : OAI21_X1 port map( B1 => n3, B2 => en, A => n94, ZN => n35);
   U10 : NAND2_X1 port map( A1 => din(29), A2 => en, ZN => n94);
   U11 : OAI21_X1 port map( B1 => n4, B2 => en, A => n93, ZN => n36);
   U12 : NAND2_X1 port map( A1 => din(28), A2 => en, ZN => n93);
   U13 : OAI21_X1 port map( B1 => n5, B2 => en, A => n92, ZN => n37);
   U14 : NAND2_X1 port map( A1 => din(27), A2 => en, ZN => n92);
   U15 : OAI21_X1 port map( B1 => n6, B2 => en, A => n91, ZN => n38);
   U16 : NAND2_X1 port map( A1 => din(26), A2 => en, ZN => n91);
   U17 : OAI21_X1 port map( B1 => n7, B2 => en, A => n90, ZN => n39);
   U18 : NAND2_X1 port map( A1 => din(25), A2 => en, ZN => n90);
   U19 : OAI21_X1 port map( B1 => n8, B2 => en, A => n89, ZN => n40);
   U20 : NAND2_X1 port map( A1 => din(24), A2 => en, ZN => n89);
   U21 : OAI21_X1 port map( B1 => n9, B2 => en, A => n88, ZN => n41);
   U22 : NAND2_X1 port map( A1 => din(23), A2 => en, ZN => n88);
   U23 : OAI21_X1 port map( B1 => n10, B2 => en, A => n87, ZN => n42);
   U24 : NAND2_X1 port map( A1 => din(22), A2 => en, ZN => n87);
   U25 : OAI21_X1 port map( B1 => n11, B2 => en, A => n86, ZN => n43);
   U26 : NAND2_X1 port map( A1 => din(21), A2 => en, ZN => n86);
   U27 : OAI21_X1 port map( B1 => n12, B2 => en, A => n85, ZN => n44);
   U28 : NAND2_X1 port map( A1 => din(20), A2 => en, ZN => n85);
   U29 : OAI21_X1 port map( B1 => n13, B2 => en, A => n84, ZN => n45);
   U30 : NAND2_X1 port map( A1 => din(19), A2 => en, ZN => n84);
   U31 : OAI21_X1 port map( B1 => n14, B2 => en, A => n83, ZN => n46);
   U32 : NAND2_X1 port map( A1 => din(18), A2 => en, ZN => n83);
   U33 : OAI21_X1 port map( B1 => n15, B2 => en, A => n82, ZN => n47);
   U34 : NAND2_X1 port map( A1 => din(17), A2 => en, ZN => n82);
   U35 : OAI21_X1 port map( B1 => n16, B2 => en, A => n81, ZN => n48);
   U36 : NAND2_X1 port map( A1 => din(16), A2 => en, ZN => n81);
   U37 : OAI21_X1 port map( B1 => n17, B2 => en, A => n80, ZN => n49);
   U38 : NAND2_X1 port map( A1 => din(15), A2 => en, ZN => n80);
   U39 : OAI21_X1 port map( B1 => n18, B2 => en, A => n79, ZN => n50);
   U40 : NAND2_X1 port map( A1 => din(14), A2 => en, ZN => n79);
   U41 : OAI21_X1 port map( B1 => n19, B2 => en, A => n78, ZN => n51);
   U42 : NAND2_X1 port map( A1 => din(13), A2 => en, ZN => n78);
   U43 : OAI21_X1 port map( B1 => n20, B2 => en, A => n77, ZN => n52);
   U44 : NAND2_X1 port map( A1 => din(12), A2 => en, ZN => n77);
   U45 : OAI21_X1 port map( B1 => n21, B2 => en, A => n76, ZN => n53);
   U46 : NAND2_X1 port map( A1 => din(11), A2 => en, ZN => n76);
   U47 : OAI21_X1 port map( B1 => n22, B2 => en, A => n75, ZN => n54);
   U48 : NAND2_X1 port map( A1 => din(10), A2 => en, ZN => n75);
   U49 : OAI21_X1 port map( B1 => n23, B2 => en, A => n74, ZN => n55);
   U50 : NAND2_X1 port map( A1 => din(9), A2 => en, ZN => n74);
   U51 : OAI21_X1 port map( B1 => n24, B2 => en, A => n73, ZN => n56);
   U52 : NAND2_X1 port map( A1 => din(8), A2 => en, ZN => n73);
   U53 : OAI21_X1 port map( B1 => n25, B2 => en, A => n72, ZN => n57);
   U54 : NAND2_X1 port map( A1 => din(7), A2 => en, ZN => n72);
   U55 : OAI21_X1 port map( B1 => n26, B2 => en, A => n71, ZN => n58);
   U56 : NAND2_X1 port map( A1 => din(6), A2 => en, ZN => n71);
   U57 : OAI21_X1 port map( B1 => n27, B2 => en, A => n70, ZN => n59);
   U58 : NAND2_X1 port map( A1 => din(5), A2 => en, ZN => n70);
   U59 : OAI21_X1 port map( B1 => n28, B2 => en, A => n69, ZN => n60);
   U60 : NAND2_X1 port map( A1 => din(4), A2 => en, ZN => n69);
   U61 : OAI21_X1 port map( B1 => n29, B2 => en, A => n68, ZN => n61);
   U62 : NAND2_X1 port map( A1 => din(3), A2 => en, ZN => n68);
   U63 : OAI21_X1 port map( B1 => n30, B2 => en, A => n67, ZN => n62);
   U64 : NAND2_X1 port map( A1 => din(2), A2 => en, ZN => n67);
   U65 : OAI21_X1 port map( B1 => n31, B2 => en, A => n66, ZN => n63);
   U66 : NAND2_X1 port map( A1 => din(1), A2 => en, ZN => n66);
   U67 : OAI21_X1 port map( B1 => n32, B2 => en, A => n65, ZN => n64);
   U68 : NAND2_X1 port map( A1 => en, A2 => din(0), ZN => n65);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux4_DATA_SIZE32 is

   port( sel : in std_logic_vector (1 downto 0);  din0, din1, din2, din3 : in 
         std_logic_vector (31 downto 0);  dout : out std_logic_vector (31 
         downto 0));

end Mux4_DATA_SIZE32;

architecture SYN_mux4_arch of Mux4_DATA_SIZE32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, 
      n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61
      , n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, 
      n76, n77, n78, n79, n80, n81, n82, n83, n84 : std_logic;

begin
   
   U3 : BUF_X1 port map( A => n8, Z => n74);
   U4 : BUF_X1 port map( A => n8, Z => n73);
   U5 : BUF_X1 port map( A => n8, Z => n75);
   U6 : BUF_X1 port map( A => n7, Z => n77);
   U7 : BUF_X1 port map( A => n5, Z => n83);
   U8 : BUF_X1 port map( A => n6, Z => n80);
   U9 : NOR2_X1 port map( A1 => n71, A2 => n72, ZN => n8);
   U10 : BUF_X1 port map( A => n7, Z => n76);
   U11 : BUF_X1 port map( A => n5, Z => n82);
   U12 : BUF_X1 port map( A => n6, Z => n79);
   U13 : BUF_X1 port map( A => n7, Z => n78);
   U14 : BUF_X1 port map( A => n5, Z => n84);
   U15 : BUF_X1 port map( A => n6, Z => n81);
   U16 : NOR2_X1 port map( A1 => sel(0), A2 => sel(1), ZN => n7);
   U17 : NOR2_X1 port map( A1 => n71, A2 => sel(1), ZN => n6);
   U18 : NOR2_X1 port map( A1 => n72, A2 => sel(0), ZN => n5);
   U19 : INV_X1 port map( A => sel(0), ZN => n71);
   U20 : INV_X1 port map( A => sel(1), ZN => n72);
   U21 : AOI22_X1 port map( A1 => din0(30), A2 => n76, B1 => din3(30), B2 => 
                           n73, ZN => n59);
   U22 : AOI22_X1 port map( A1 => din0(31), A2 => n78, B1 => din3(31), B2 => 
                           n75, ZN => n3);
   U23 : AOI22_X1 port map( A1 => din0(29), A2 => n76, B1 => din3(29), B2 => 
                           n73, ZN => n61);
   U24 : AOI22_X1 port map( A1 => din2(29), A2 => n82, B1 => din1(29), B2 => 
                           n79, ZN => n62);
   U25 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => dout(23));
   U26 : AOI22_X1 port map( A1 => din0(23), A2 => n78, B1 => din3(23), B2 => 
                           n75, ZN => n11);
   U27 : AOI22_X1 port map( A1 => din2(23), A2 => n84, B1 => din1(23), B2 => 
                           n81, ZN => n12);
   U28 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => dout(16));
   U29 : AOI22_X1 port map( A1 => din0(16), A2 => n77, B1 => din3(16), B2 => 
                           n74, ZN => n25);
   U30 : AOI22_X1 port map( A1 => din2(16), A2 => n83, B1 => din1(16), B2 => 
                           n80, ZN => n26);
   U31 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => dout(17));
   U32 : AOI22_X1 port map( A1 => din0(17), A2 => n77, B1 => din3(17), B2 => 
                           n74, ZN => n23);
   U33 : AOI22_X1 port map( A1 => din2(17), A2 => n83, B1 => din1(17), B2 => 
                           n80, ZN => n24);
   U34 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => dout(6));
   U35 : AOI22_X1 port map( A1 => din2(6), A2 => n83, B1 => din1(6), B2 => n80,
                           ZN => n46);
   U36 : AOI22_X1 port map( A1 => din0(6), A2 => n77, B1 => din3(6), B2 => n74,
                           ZN => n45);
   U37 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => dout(7));
   U38 : AOI22_X1 port map( A1 => din2(7), A2 => n83, B1 => din1(7), B2 => n80,
                           ZN => n44);
   U39 : AOI22_X1 port map( A1 => din0(7), A2 => n77, B1 => din3(7), B2 => n74,
                           ZN => n43);
   U40 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => dout(8));
   U41 : AOI22_X1 port map( A1 => din2(8), A2 => n83, B1 => din1(8), B2 => n80,
                           ZN => n42);
   U42 : AOI22_X1 port map( A1 => din0(8), A2 => n77, B1 => din3(8), B2 => n74,
                           ZN => n41);
   U43 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => dout(9));
   U44 : AOI22_X1 port map( A1 => din2(9), A2 => n83, B1 => din1(9), B2 => n80,
                           ZN => n40);
   U45 : AOI22_X1 port map( A1 => din0(9), A2 => n77, B1 => din3(9), B2 => n74,
                           ZN => n39);
   U46 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => dout(10));
   U47 : AOI22_X1 port map( A1 => din2(10), A2 => n83, B1 => din1(10), B2 => 
                           n80, ZN => n38);
   U48 : AOI22_X1 port map( A1 => din0(10), A2 => n77, B1 => din3(10), B2 => 
                           n74, ZN => n37);
   U49 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => dout(11));
   U50 : AOI22_X1 port map( A1 => din2(11), A2 => n83, B1 => din1(11), B2 => 
                           n80, ZN => n36);
   U51 : AOI22_X1 port map( A1 => din0(11), A2 => n77, B1 => din3(11), B2 => 
                           n74, ZN => n35);
   U52 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => dout(12));
   U53 : AOI22_X1 port map( A1 => din0(12), A2 => n77, B1 => din3(12), B2 => 
                           n74, ZN => n33);
   U54 : AOI22_X1 port map( A1 => din2(12), A2 => n83, B1 => din1(12), B2 => 
                           n80, ZN => n34);
   U55 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => dout(13));
   U56 : AOI22_X1 port map( A1 => din0(13), A2 => n77, B1 => din3(13), B2 => 
                           n74, ZN => n31);
   U57 : AOI22_X1 port map( A1 => din2(13), A2 => n83, B1 => din1(13), B2 => 
                           n80, ZN => n32);
   U58 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => dout(14));
   U59 : AOI22_X1 port map( A1 => din0(14), A2 => n77, B1 => din3(14), B2 => 
                           n74, ZN => n29);
   U60 : AOI22_X1 port map( A1 => din2(14), A2 => n83, B1 => din1(14), B2 => 
                           n80, ZN => n30);
   U61 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => dout(15));
   U62 : AOI22_X1 port map( A1 => din0(15), A2 => n77, B1 => din3(15), B2 => 
                           n74, ZN => n27);
   U63 : AOI22_X1 port map( A1 => din2(15), A2 => n83, B1 => din1(15), B2 => 
                           n80, ZN => n28);
   U64 : NAND2_X1 port map( A1 => n64, A2 => n63, ZN => dout(28));
   U65 : AOI22_X1 port map( A1 => din0(28), A2 => n76, B1 => din3(28), B2 => 
                           n73, ZN => n63);
   U66 : AOI22_X1 port map( A1 => din2(28), A2 => n82, B1 => din1(28), B2 => 
                           n79, ZN => n64);
   U67 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => dout(27));
   U68 : AOI22_X1 port map( A1 => din0(27), A2 => n76, B1 => din3(27), B2 => 
                           n73, ZN => n65);
   U69 : AOI22_X1 port map( A1 => din2(27), A2 => n82, B1 => din1(27), B2 => 
                           n79, ZN => n66);
   U70 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => dout(25));
   U71 : AOI22_X1 port map( A1 => din0(25), A2 => n76, B1 => din3(25), B2 => 
                           n73, ZN => n69);
   U72 : AOI22_X1 port map( A1 => din2(25), A2 => n82, B1 => din1(25), B2 => 
                           n79, ZN => n70);
   U73 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => dout(26));
   U74 : AOI22_X1 port map( A1 => din0(26), A2 => n76, B1 => din3(26), B2 => 
                           n73, ZN => n67);
   U75 : AOI22_X1 port map( A1 => din2(26), A2 => n82, B1 => din1(26), B2 => 
                           n79, ZN => n68);
   U76 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => dout(1));
   U77 : AOI22_X1 port map( A1 => din2(1), A2 => n82, B1 => din1(1), B2 => n79,
                           ZN => n56);
   U78 : AOI22_X1 port map( A1 => din0(1), A2 => n76, B1 => din3(1), B2 => n73,
                           ZN => n55);
   U79 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => dout(2));
   U80 : AOI22_X1 port map( A1 => din2(2), A2 => n82, B1 => din1(2), B2 => n79,
                           ZN => n54);
   U81 : AOI22_X1 port map( A1 => din0(2), A2 => n76, B1 => din3(2), B2 => n73,
                           ZN => n53);
   U82 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => dout(3));
   U83 : AOI22_X1 port map( A1 => din2(3), A2 => n82, B1 => din1(3), B2 => n79,
                           ZN => n52);
   U84 : AOI22_X1 port map( A1 => din0(3), A2 => n76, B1 => din3(3), B2 => n73,
                           ZN => n51);
   U85 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => dout(4));
   U86 : AOI22_X1 port map( A1 => din2(4), A2 => n82, B1 => din1(4), B2 => n79,
                           ZN => n50);
   U87 : AOI22_X1 port map( A1 => din0(4), A2 => n76, B1 => din3(4), B2 => n73,
                           ZN => n49);
   U88 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => dout(5));
   U89 : AOI22_X1 port map( A1 => din2(5), A2 => n82, B1 => din1(5), B2 => n79,
                           ZN => n48);
   U90 : AOI22_X1 port map( A1 => din0(5), A2 => n76, B1 => din3(5), B2 => n73,
                           ZN => n47);
   U91 : NAND2_X1 port map( A1 => n9, A2 => n10, ZN => dout(24));
   U92 : AOI22_X1 port map( A1 => din0(24), A2 => n78, B1 => din3(24), B2 => 
                           n75, ZN => n9);
   U93 : AOI22_X1 port map( A1 => din2(24), A2 => n84, B1 => din1(24), B2 => 
                           n81, ZN => n10);
   U94 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => dout(18));
   U95 : AOI22_X1 port map( A1 => din0(18), A2 => n78, B1 => din3(18), B2 => 
                           n75, ZN => n21);
   U96 : AOI22_X1 port map( A1 => din2(18), A2 => n84, B1 => din1(18), B2 => 
                           n81, ZN => n22);
   U97 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => dout(19));
   U98 : AOI22_X1 port map( A1 => din0(19), A2 => n78, B1 => din3(19), B2 => 
                           n75, ZN => n19);
   U99 : AOI22_X1 port map( A1 => din2(19), A2 => n84, B1 => din1(19), B2 => 
                           n81, ZN => n20);
   U100 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => dout(20));
   U101 : AOI22_X1 port map( A1 => din0(20), A2 => n78, B1 => din3(20), B2 => 
                           n75, ZN => n17);
   U102 : AOI22_X1 port map( A1 => din2(20), A2 => n84, B1 => din1(20), B2 => 
                           n81, ZN => n18);
   U103 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => dout(21));
   U104 : AOI22_X1 port map( A1 => din0(21), A2 => n78, B1 => din3(21), B2 => 
                           n75, ZN => n15);
   U105 : AOI22_X1 port map( A1 => din2(21), A2 => n84, B1 => din1(21), B2 => 
                           n81, ZN => n16);
   U106 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => dout(22));
   U107 : AOI22_X1 port map( A1 => din0(22), A2 => n78, B1 => din3(22), B2 => 
                           n75, ZN => n13);
   U108 : AOI22_X1 port map( A1 => din2(22), A2 => n84, B1 => din1(22), B2 => 
                           n81, ZN => n14);
   U109 : AOI22_X1 port map( A1 => din2(0), A2 => n82, B1 => din1(0), B2 => n79
                           , ZN => n58);
   U110 : NAND2_X1 port map( A1 => n60, A2 => n59, ZN => dout(30));
   U111 : AOI22_X1 port map( A1 => din2(30), A2 => n82, B1 => din1(30), B2 => 
                           n79, ZN => n60);
   U112 : NAND2_X1 port map( A1 => n62, A2 => n61, ZN => dout(29));
   U113 : NAND2_X1 port map( A1 => n4, A2 => n3, ZN => dout(31));
   U114 : AOI22_X1 port map( A1 => din2(31), A2 => n84, B1 => din1(31), B2 => 
                           n81, ZN => n4);
   U115 : AOI22_X1 port map( A1 => din0(0), A2 => n76, B1 => din3(0), B2 => n73
                           , ZN => n57);
   U116 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => dout(0));

end SYN_mux4_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Div_DATA_SIZE32_DIV_STAGE34_SQRT_STAGE18 is

   port( rst, clk, en, lock, sign, func : in std_logic;  a, b : in 
         std_logic_vector (31 downto 0);  o : out std_logic_vector (31 downto 
         0));

end Div_DATA_SIZE32_DIV_STAGE34_SQRT_STAGE18;

architecture SYN_div_arch of Div_DATA_SIZE32_DIV_STAGE34_SQRT_STAGE18 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component Div_DATA_SIZE32_DIV_STAGE34_SQRT_STAGE18_DW01_inc_0
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component AddSub_DATA_SIZE32_2
      port( as : in std_logic;  a, b : in std_logic_vector (31 downto 0);  re :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;
   
   component Sipo_DATA_SIZE32
      port( rst, en, clk, din : in std_logic;  dout : out std_logic_vector (31 
            downto 0));
   end component;
   
   component Reg_DATA_SIZE64
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (63 downto 
            0);  dout : out std_logic_vector (63 downto 0));
   end component;
   
   component AddSub_DATA_SIZE64
      port( as : in std_logic;  a, b : in std_logic_vector (63 downto 0);  re :
            out std_logic_vector (63 downto 0);  cout : out std_logic);
   end component;
   
   component Mux_DATA_SIZE64
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (63 downto 0)
            ;  dout : out std_logic_vector (63 downto 0));
   end component;
   
   component AddSub_DATA_SIZE32_3
      port( as : in std_logic;  a, b : in std_logic_vector (31 downto 0);  re :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;
   
   component AddSub_DATA_SIZE32_0
      port( as : in std_logic;  a, b : in std_logic_vector (31 downto 0);  re :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic0_port, a_mod_63_port, a_mod_62_port, a_mod_61_port, 
      a_mod_60_port, a_mod_59_port, a_mod_58_port, a_mod_57_port, a_mod_56_port
      , a_mod_55_port, a_mod_54_port, a_mod_53_port, a_mod_52_port, 
      a_mod_51_port, a_mod_50_port, a_mod_49_port, a_mod_48_port, a_mod_47_port
      , a_mod_46_port, a_mod_45_port, a_mod_44_port, a_mod_43_port, 
      a_mod_42_port, a_mod_41_port, a_mod_40_port, a_mod_39_port, a_mod_38_port
      , a_mod_37_port, a_mod_36_port, a_mod_35_port, a_mod_34_port, 
      a_mod_33_port, a_mod_32_port, a_mod_27_port, a_mod_26_port, a_mod_25_port
      , a_mod_24_port, a_mod_23_port, a_mod_22_port, a_mod_21_port, 
      a_mod_20_port, a_mod_19_port, a_mod_18_port, a_mod_17_port, a_mod_16_port
      , a_mod_15_port, a_mod_14_port, a_mod_13_port, a_mod_12_port, 
      a_mod_11_port, a_mod_10_port, a_mod_9_port, a_mod_8_port, a_mod_7_port, 
      a_mod_6_port, a_mod_5_port, a_mod_4_port, a_mod_3_port, a_mod_2_port, 
      a_mod_1_port, a_mod_0_port, a_adj_31_port, a_adj_30_port, a_adj_29_port, 
      a_adj_28_port, a_adj_27_port, a_adj_26_port, a_adj_25_port, a_adj_24_port
      , a_adj_23_port, a_adj_22_port, a_adj_21_port, a_adj_20_port, 
      a_adj_19_port, a_adj_18_port, a_adj_17_port, a_adj_16_port, a_adj_15_port
      , a_adj_14_port, a_adj_13_port, a_adj_12_port, a_adj_11_port, 
      a_adj_10_port, a_adj_9_port, a_adj_8_port, a_adj_7_port, a_adj_6_port, 
      a_adj_5_port, a_adj_4_port, a_adj_3_port, a_adj_2_port, a_adj_1_port, 
      a_adj_0_port, b_adj_31_port, b_adj_30_port, b_adj_29_port, b_adj_28_port,
      b_adj_27_port, b_adj_26_port, b_adj_25_port, b_adj_24_port, b_adj_23_port
      , b_adj_22_port, b_adj_21_port, b_adj_20_port, b_adj_19_port, 
      b_adj_18_port, b_adj_17_port, b_adj_16_port, b_adj_15_port, b_adj_14_port
      , b_adj_13_port, b_adj_12_port, b_adj_11_port, b_adj_10_port, 
      b_adj_9_port, b_adj_8_port, b_adj_7_port, b_adj_6_port, b_adj_5_port, 
      b_adj_4_port, b_adj_3_port, b_adj_2_port, b_adj_1_port, b_adj_0_port, 
      r_63_port, r_62_port, r_61_port, r_60_port, r_59_port, r_58_port, 
      r_57_port, r_56_port, r_55_port, r_54_port, r_53_port, r_52_port, 
      r_51_port, r_50_port, r_49_port, r_48_port, r_47_port, r_46_port, 
      r_45_port, r_44_port, r_43_port, r_42_port, r_41_port, r_40_port, 
      r_39_port, r_38_port, r_37_port, r_36_port, r_35_port, r_34_port, 
      r_33_port, r_32_port, r_31_port, r_30_port, r_29_port, r_28_port, 
      r_27_port, r_26_port, r_25_port, r_24_port, r_23_port, r_22_port, 
      r_21_port, r_20_port, r_19_port, r_18_port, r_17_port, r_16_port, 
      r_15_port, r_14_port, r_13_port, r_12_port, r_11_port, r_10_port, 
      r_9_port, r_8_port, r_7_port, r_6_port, r_5_port, r_4_port, r_3_port, 
      r_2_port, r_1_port, r_0_port, a_mux_63_port, a_mux_62_port, a_mux_61_port
      , a_mux_60_port, a_mux_59_port, a_mux_58_port, a_mux_57_port, 
      a_mux_56_port, a_mux_55_port, a_mux_54_port, a_mux_53_port, a_mux_52_port
      , a_mux_51_port, a_mux_50_port, a_mux_49_port, a_mux_48_port, 
      a_mux_47_port, a_mux_46_port, a_mux_45_port, a_mux_44_port, a_mux_43_port
      , a_mux_42_port, a_mux_41_port, a_mux_40_port, a_mux_39_port, 
      a_mux_38_port, a_mux_37_port, a_mux_36_port, a_mux_35_port, a_mux_34_port
      , a_mux_33_port, a_mux_32_port, a_mux_31_port, a_mux_30_port, 
      a_mux_29_port, a_mux_28_port, a_mux_27_port, a_mux_26_port, a_mux_25_port
      , a_mux_24_port, a_mux_23_port, a_mux_22_port, a_mux_21_port, 
      a_mux_20_port, a_mux_19_port, a_mux_18_port, a_mux_17_port, a_mux_16_port
      , a_mux_15_port, a_mux_14_port, a_mux_13_port, a_mux_12_port, 
      a_mux_11_port, a_mux_10_port, a_mux_9_port, a_mux_8_port, a_mux_7_port, 
      a_mux_6_port, a_mux_5_port, a_mux_4_port, a_mux_3_port, a_mux_2_port, 
      a_mux_1_port, a_mux_0_port, not_r_sign, a_shf_1_port, q_31_port, 
      q_30_port, b_shf_sqrt_63_port, b_shf_sqrt_62_port, b_shf_sqrt_61_port, 
      b_shf_sqrt_60_port, b_shf_sqrt_59_port, b_shf_sqrt_58_port, 
      b_shf_sqrt_57_port, b_shf_sqrt_56_port, b_shf_sqrt_55_port, 
      b_shf_sqrt_54_port, b_shf_sqrt_53_port, b_shf_sqrt_52_port, 
      b_shf_sqrt_51_port, b_shf_sqrt_50_port, b_shf_sqrt_49_port, 
      b_shf_sqrt_48_port, b_shf_sqrt_47_port, b_shf_sqrt_46_port, 
      b_shf_sqrt_45_port, b_shf_sqrt_44_port, b_shf_sqrt_43_port, 
      b_shf_sqrt_42_port, b_shf_sqrt_41_port, b_shf_sqrt_40_port, 
      b_shf_sqrt_39_port, b_shf_sqrt_38_port, b_shf_sqrt_37_port, 
      b_shf_sqrt_36_port, b_shf_sqrt_35_port, b_shf_sqrt_34_port, b_shf_63_port
      , b_shf_62_port, b_shf_61_port, b_shf_60_port, b_shf_59_port, 
      b_shf_58_port, b_shf_57_port, b_shf_56_port, b_shf_55_port, b_shf_54_port
      , b_shf_53_port, b_shf_52_port, b_shf_51_port, b_shf_50_port, 
      b_shf_49_port, b_shf_48_port, b_shf_47_port, b_shf_46_port, b_shf_45_port
      , b_shf_44_port, b_shf_43_port, b_shf_42_port, b_shf_41_port, 
      b_shf_40_port, b_shf_39_port, b_shf_38_port, b_shf_37_port, b_shf_36_port
      , b_shf_35_port, b_shf_34_port, b_shf_33_port, b_shf_32_port, 
      b_shf_31_port, b_shf_30_port, b_shf_29_port, b_shf_28_port, b_shf_27_port
      , b_shf_26_port, b_shf_25_port, b_shf_24_port, b_shf_23_port, 
      b_shf_22_port, b_shf_21_port, b_shf_20_port, b_shf_19_port, b_shf_18_port
      , b_shf_17_port, b_shf_16_port, b_shf_15_port, b_shf_14_port, 
      b_shf_13_port, b_shf_12_port, b_shf_11_port, b_shf_10_port, b_shf_9_port,
      b_shf_8_port, b_shf_7_port, b_shf_6_port, b_shf_5_port, b_shf_4_port, 
      b_shf_3_port, b_shf_2_port, b_shf_1_port, b_shf_0_port, r_es_63_port, 
      r_es_62_port, r_es_61_port, r_es_60_port, r_es_59_port, r_es_58_port, 
      r_es_57_port, r_es_56_port, r_es_55_port, r_es_54_port, r_es_53_port, 
      r_es_52_port, r_es_51_port, r_es_50_port, r_es_49_port, r_es_48_port, 
      r_es_47_port, r_es_46_port, r_es_45_port, r_es_44_port, r_es_43_port, 
      r_es_42_port, r_es_41_port, r_es_40_port, r_es_39_port, r_es_38_port, 
      r_es_37_port, r_es_36_port, r_es_35_port, r_es_34_port, r_es_33_port, 
      r_es_32_port, r_es_31_port, r_es_30_port, r_es_29_port, r_es_28_port, 
      r_es_27_port, r_es_26_port, r_es_25_port, r_es_24_port, r_es_23_port, 
      r_es_22_port, r_es_21_port, r_es_20_port, r_es_19_port, r_es_18_port, 
      r_es_17_port, r_es_16_port, r_es_15_port, r_es_14_port, r_es_13_port, 
      r_es_12_port, r_es_11_port, r_es_10_port, r_es_9_port, r_es_8_port, 
      r_es_7_port, r_es_6_port, r_es_5_port, r_es_4_port, r_es_3_port, 
      r_es_2_port, r_es_1_port, r_es_0_port, not_r_es_sign, n_state_31_port, 
      n_state_30_port, n_state_29_port, n_state_28_port, n_state_27_port, 
      n_state_26_port, n_state_25_port, n_state_24_port, n_state_23_port, 
      n_state_22_port, n_state_21_port, n_state_20_port, n_state_19_port, 
      n_state_18_port, n_state_17_port, n_state_16_port, n_state_15_port, 
      n_state_14_port, n_state_13_port, n_state_12_port, n_state_11_port, 
      n_state_10_port, n_state_9_port, n_state_8_port, n_state_7_port, 
      n_state_6_port, n_state_5_port, n_state_4_port, n_state_3_port, 
      n_state_2_port, n_state_1_port, c_state_31_port, c_state_29_port, 
      c_state_28_port, c_state_27_port, c_state_26_port, c_state_24_port, 
      c_state_23_port, c_state_22_port, c_state_21_port, c_state_20_port, 
      c_state_19_port, c_state_17_port, c_state_16_port, c_state_15_port, 
      c_state_14_port, c_state_13_port, c_state_12_port, c_state_11_port, 
      c_state_10_port, c_state_9_port, c_state_8_port, c_state_7_port, 
      c_state_6_port, c_state_5_port, c_state_4_port, c_state_3_port, 
      c_state_2_port, c_state_1_port, c_state_0_port, N17, N18, N19, N20, N21, 
      N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36
      , N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, net3927, 
      net3928, net3929, net3930, n297, n298, n299, n300, n301, n302, n303, n304
      , n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
      n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, 
      n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, 
      n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, 
      n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n372, n373, 
      n374, n71, n72, n73, n76, n77, n78, n80, n81, n82, net108616, net108617, 
      net108618, net108619, net108620, net108621, net108622, net108623, 
      net108624, net108625, net108626, net108627, net108628, net108629, 
      net108630, net108631, net108632, net108633, net108634, net108635, 
      net108636, net108637, net108638, net108639, net108640, net108641, 
      net108642, net108643, net108644, net108645, net108646, net108650, 
      net108651, net108652, net108653, net108654, net108655, net108656, 
      net108657, net108658, net108659, net108660, net108661, net108662, 
      net108663, net108664, net108665, net108666, net108667, net108668, 
      net108669, net108670, net108671, net108672, net108673, net108674, 
      net108675, net108676, net108677, net108678, net108680, net108681, 
      net108685, net108686, net108687, n224, n225, n226, n227, n228, n229, n230
      , n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n87, 
      n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, 
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, 
      n222, n223, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, 
      n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, 
      n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, 
      n288, n289, n290, n291, n292, n293, n294, n295, n296, n363, n364, n365, 
      n366, n367, n368, n369, n370, n371, n375, n376, n377, n378, n379, n380, 
      n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, 
      net164131, net164132 : std_logic;

begin
   
   X_Logic0_port <= '0';
   c_state_reg_0_inst : DFFR_X1 port map( D => n259, CK => clk, RN => n173, Q 
                           => c_state_0_port, QN => n362);
   c_state_reg_10_inst : DFFR_X1 port map( D => n_state_10_port, CK => clk, RN 
                           => n172, Q => c_state_10_port, QN => n91);
   c_state_reg_1_inst : DFFR_X1 port map( D => n_state_1_port, CK => clk, RN =>
                           n173, Q => c_state_1_port, QN => n373);
   c_state_reg_2_inst : DFFR_X1 port map( D => n_state_2_port, CK => clk, RN =>
                           n173, Q => c_state_2_port, QN => n77);
   c_state_reg_3_inst : DFFR_X1 port map( D => n_state_3_port, CK => clk, RN =>
                           n173, Q => c_state_3_port, QN => n78);
   c_state_reg_4_inst : DFFR_X1 port map( D => n_state_4_port, CK => clk, RN =>
                           n173, Q => c_state_4_port, QN => n76);
   c_state_reg_5_inst : DFFR_X1 port map( D => n_state_5_port, CK => clk, RN =>
                           n173, Q => c_state_5_port, QN => n82);
   c_state_reg_6_inst : DFFR_X1 port map( D => n_state_6_port, CK => clk, RN =>
                           n173, Q => c_state_6_port, QN => n100);
   c_state_reg_7_inst : DFFR_X1 port map( D => n_state_7_port, CK => clk, RN =>
                           n173, Q => c_state_7_port, QN => n80);
   c_state_reg_8_inst : DFFR_X1 port map( D => n_state_8_port, CK => clk, RN =>
                           n173, Q => c_state_8_port, QN => n81);
   c_state_reg_9_inst : DFFR_X1 port map( D => n_state_9_port, CK => clk, RN =>
                           n173, Q => c_state_9_port, QN => n95);
   c_state_reg_11_inst : DFFR_X1 port map( D => n_state_11_port, CK => clk, RN 
                           => n172, Q => c_state_11_port, QN => n92);
   c_state_reg_12_inst : DFFR_X1 port map( D => n_state_12_port, CK => clk, RN 
                           => n172, Q => c_state_12_port, QN => net108687);
   c_state_reg_13_inst : DFFR_X1 port map( D => n_state_13_port, CK => clk, RN 
                           => n172, Q => c_state_13_port, QN => n101);
   c_state_reg_14_inst : DFFR_X1 port map( D => n_state_14_port, CK => clk, RN 
                           => n172, Q => c_state_14_port, QN => n96);
   c_state_reg_15_inst : DFFR_X1 port map( D => n_state_15_port, CK => clk, RN 
                           => n172, Q => c_state_15_port, QN => n73);
   c_state_reg_16_inst : DFFR_X1 port map( D => n_state_16_port, CK => clk, RN 
                           => n172, Q => c_state_16_port, QN => net108686);
   c_state_reg_17_inst : DFFR_X1 port map( D => n_state_17_port, CK => clk, RN 
                           => n172, Q => c_state_17_port, QN => net108685);
   c_state_reg_18_inst : DFFR_X1 port map( D => n_state_18_port, CK => clk, RN 
                           => n172, Q => n186, QN => n146);
   c_state_reg_19_inst : DFFR_X1 port map( D => n_state_19_port, CK => clk, RN 
                           => n172, Q => c_state_19_port, QN => n372);
   c_state_reg_20_inst : DFFR_X1 port map( D => n_state_20_port, CK => clk, RN 
                           => n172, Q => c_state_20_port, QN => n374);
   c_state_reg_21_inst : DFFR_X1 port map( D => n_state_21_port, CK => clk, RN 
                           => n172, Q => c_state_21_port, QN => n89);
   c_state_reg_22_inst : DFFR_X1 port map( D => n_state_22_port, CK => clk, RN 
                           => n172, Q => c_state_22_port, QN => n98);
   c_state_reg_23_inst : DFFR_X1 port map( D => n_state_23_port, CK => clk, RN 
                           => n172, Q => c_state_23_port, QN => n93);
   c_state_reg_24_inst : DFFR_X1 port map( D => n_state_24_port, CK => clk, RN 
                           => n172, Q => c_state_24_port, QN => n90);
   c_state_reg_25_inst : DFFR_X1 port map( D => n_state_25_port, CK => clk, RN 
                           => n172, Q => n178, QN => net164132);
   c_state_reg_26_inst : DFFR_X1 port map( D => n_state_26_port, CK => clk, RN 
                           => n173, Q => c_state_26_port, QN => n99);
   c_state_reg_27_inst : DFFR_X1 port map( D => n_state_27_port, CK => clk, RN 
                           => n173, Q => c_state_27_port, QN => n94);
   c_state_reg_28_inst : DFFR_X1 port map( D => n_state_28_port, CK => clk, RN 
                           => n173, Q => c_state_28_port, QN => net108681);
   c_state_reg_29_inst : DFFR_X1 port map( D => n_state_29_port, CK => clk, RN 
                           => n173, Q => c_state_29_port, QN => net108680);
   c_state_reg_30_inst : DFFR_X1 port map( D => n_state_30_port, CK => clk, RN 
                           => n173, Q => n180, QN => net164131);
   c_state_reg_31_inst : DFFR_X1 port map( D => n_state_31_port, CK => clk, RN 
                           => n173, Q => c_state_31_port, QN => n72);
   a_mod_reg_0_inst : DFF_X1 port map( D => n361, CK => clk, Q => a_mod_0_port,
                           QN => net108678);
   a_mod_reg_1_inst : DFF_X1 port map( D => n360, CK => clk, Q => a_mod_1_port,
                           QN => net108677);
   a_mod_reg_2_inst : DFF_X1 port map( D => n359, CK => clk, Q => a_mod_2_port,
                           QN => net108676);
   a_mod_reg_3_inst : DFF_X1 port map( D => n358, CK => clk, Q => a_mod_3_port,
                           QN => net108675);
   a_mod_reg_4_inst : DFF_X1 port map( D => n357, CK => clk, Q => a_mod_4_port,
                           QN => net108674);
   a_mod_reg_5_inst : DFF_X1 port map( D => n356, CK => clk, Q => a_mod_5_port,
                           QN => net108673);
   a_mod_reg_6_inst : DFF_X1 port map( D => n355, CK => clk, Q => a_mod_6_port,
                           QN => net108672);
   a_mod_reg_7_inst : DFF_X1 port map( D => n354, CK => clk, Q => a_mod_7_port,
                           QN => net108671);
   a_mod_reg_8_inst : DFF_X1 port map( D => n353, CK => clk, Q => a_mod_8_port,
                           QN => net108670);
   a_mod_reg_9_inst : DFF_X1 port map( D => n352, CK => clk, Q => a_mod_9_port,
                           QN => net108669);
   a_mod_reg_10_inst : DFF_X1 port map( D => n351, CK => clk, Q => 
                           a_mod_10_port, QN => net108668);
   a_mod_reg_11_inst : DFF_X1 port map( D => n350, CK => clk, Q => 
                           a_mod_11_port, QN => net108667);
   a_mod_reg_12_inst : DFF_X1 port map( D => n349, CK => clk, Q => 
                           a_mod_12_port, QN => net108666);
   a_mod_reg_13_inst : DFF_X1 port map( D => n348, CK => clk, Q => 
                           a_mod_13_port, QN => net108665);
   a_mod_reg_14_inst : DFF_X1 port map( D => n347, CK => clk, Q => 
                           a_mod_14_port, QN => net108664);
   a_mod_reg_15_inst : DFF_X1 port map( D => n346, CK => clk, Q => 
                           a_mod_15_port, QN => net108663);
   a_mod_reg_16_inst : DFF_X1 port map( D => n345, CK => clk, Q => 
                           a_mod_16_port, QN => net108662);
   a_mod_reg_17_inst : DFF_X1 port map( D => n344, CK => clk, Q => 
                           a_mod_17_port, QN => net108661);
   a_mod_reg_18_inst : DFF_X1 port map( D => n343, CK => clk, Q => 
                           a_mod_18_port, QN => net108660);
   a_mod_reg_19_inst : DFF_X1 port map( D => n342, CK => clk, Q => 
                           a_mod_19_port, QN => net108659);
   a_mod_reg_20_inst : DFF_X1 port map( D => n341, CK => clk, Q => 
                           a_mod_20_port, QN => net108658);
   a_mod_reg_21_inst : DFF_X1 port map( D => n340, CK => clk, Q => 
                           a_mod_21_port, QN => net108657);
   a_mod_reg_22_inst : DFF_X1 port map( D => n339, CK => clk, Q => 
                           a_mod_22_port, QN => net108656);
   a_mod_reg_23_inst : DFF_X1 port map( D => n338, CK => clk, Q => 
                           a_mod_23_port, QN => net108655);
   a_mod_reg_24_inst : DFF_X1 port map( D => n337, CK => clk, Q => 
                           a_mod_24_port, QN => net108654);
   a_mod_reg_25_inst : DFF_X1 port map( D => n336, CK => clk, Q => 
                           a_mod_25_port, QN => net108653);
   a_mod_reg_26_inst : DFF_X1 port map( D => n335, CK => clk, Q => 
                           a_mod_26_port, QN => net108652);
   a_mod_reg_27_inst : DFF_X1 port map( D => n334, CK => clk, Q => 
                           a_mod_27_port, QN => net108651);
   a_mod_reg_28_inst : DFF_X1 port map( D => n333, CK => clk, Q => n221, QN => 
                           net108650);
   b_mod_reg_32_inst : DFF_X1 port map( D => n329, CK => clk, Q => n129, QN => 
                           n71);
   b_mod_reg_33_inst : DFF_X1 port map( D => n328, CK => clk, Q => n97, QN => 
                           net108646);
   b_mod_reg_34_inst : DFF_X1 port map( D => n327, CK => clk, Q => n128, QN => 
                           net108645);
   b_mod_reg_35_inst : DFF_X1 port map( D => n326, CK => clk, Q => n127, QN => 
                           net108644);
   b_mod_reg_36_inst : DFF_X1 port map( D => n325, CK => clk, Q => n126, QN => 
                           net108643);
   b_mod_reg_37_inst : DFF_X1 port map( D => n324, CK => clk, Q => n125, QN => 
                           net108642);
   b_mod_reg_38_inst : DFF_X1 port map( D => n323, CK => clk, Q => n124, QN => 
                           net108641);
   b_mod_reg_39_inst : DFF_X1 port map( D => n322, CK => clk, Q => n123, QN => 
                           net108640);
   b_mod_reg_40_inst : DFF_X1 port map( D => n321, CK => clk, Q => n122, QN => 
                           net108639);
   b_mod_reg_41_inst : DFF_X1 port map( D => n320, CK => clk, Q => n121, QN => 
                           net108638);
   b_mod_reg_42_inst : DFF_X1 port map( D => n319, CK => clk, Q => n120, QN => 
                           net108637);
   b_mod_reg_43_inst : DFF_X1 port map( D => n318, CK => clk, Q => n119, QN => 
                           net108636);
   b_mod_reg_44_inst : DFF_X1 port map( D => n317, CK => clk, Q => n118, QN => 
                           net108635);
   b_mod_reg_45_inst : DFF_X1 port map( D => n316, CK => clk, Q => n117, QN => 
                           net108634);
   b_mod_reg_46_inst : DFF_X1 port map( D => n315, CK => clk, Q => n116, QN => 
                           net108633);
   b_mod_reg_47_inst : DFF_X1 port map( D => n314, CK => clk, Q => n115, QN => 
                           net108632);
   b_mod_reg_48_inst : DFF_X1 port map( D => n313, CK => clk, Q => n114, QN => 
                           net108631);
   b_mod_reg_49_inst : DFF_X1 port map( D => n312, CK => clk, Q => n113, QN => 
                           net108630);
   b_mod_reg_50_inst : DFF_X1 port map( D => n311, CK => clk, Q => n112, QN => 
                           net108629);
   b_mod_reg_51_inst : DFF_X1 port map( D => n310, CK => clk, Q => n111, QN => 
                           net108628);
   b_mod_reg_52_inst : DFF_X1 port map( D => n309, CK => clk, Q => n110, QN => 
                           net108627);
   b_mod_reg_53_inst : DFF_X1 port map( D => n308, CK => clk, Q => n109, QN => 
                           net108626);
   b_mod_reg_54_inst : DFF_X1 port map( D => n307, CK => clk, Q => n108, QN => 
                           net108625);
   b_mod_reg_55_inst : DFF_X1 port map( D => n306, CK => clk, Q => n107, QN => 
                           net108624);
   b_mod_reg_56_inst : DFF_X1 port map( D => n305, CK => clk, Q => n106, QN => 
                           net108623);
   b_mod_reg_57_inst : DFF_X1 port map( D => n304, CK => clk, Q => n105, QN => 
                           net108622);
   b_mod_reg_58_inst : DFF_X1 port map( D => n303, CK => clk, Q => n104, QN => 
                           net108621);
   b_mod_reg_59_inst : DFF_X1 port map( D => n302, CK => clk, Q => n103, QN => 
                           net108620);
   b_mod_reg_60_inst : DFF_X1 port map( D => n301, CK => clk, Q => n217, QN => 
                           net108619);
   b_mod_reg_61_inst : DFF_X1 port map( D => n300, CK => clk, Q => n216, QN => 
                           net108618);
   b_shf_31_port <= '0';
   b_shf_30_port <= '0';
   b_shf_29_port <= '0';
   b_shf_28_port <= '0';
   b_shf_27_port <= '0';
   b_shf_26_port <= '0';
   b_shf_25_port <= '0';
   b_shf_24_port <= '0';
   b_shf_23_port <= '0';
   b_shf_22_port <= '0';
   b_shf_21_port <= '0';
   b_shf_20_port <= '0';
   b_shf_19_port <= '0';
   b_shf_18_port <= '0';
   b_shf_17_port <= '0';
   b_shf_16_port <= '0';
   b_shf_15_port <= '0';
   b_shf_14_port <= '0';
   b_shf_13_port <= '0';
   b_shf_12_port <= '0';
   b_shf_11_port <= '0';
   b_shf_10_port <= '0';
   b_shf_9_port <= '0';
   b_shf_8_port <= '0';
   b_shf_7_port <= '0';
   b_shf_6_port <= '0';
   b_shf_5_port <= '0';
   b_shf_4_port <= '0';
   b_shf_3_port <= '0';
   b_shf_2_port <= '0';
   b_shf_1_port <= '0';
   b_shf_0_port <= '0';
   a_mod_63_port <= '0';
   a_mod_62_port <= '0';
   a_mod_61_port <= '0';
   a_mod_60_port <= '0';
   a_mod_59_port <= '0';
   a_mod_58_port <= '0';
   a_mod_57_port <= '0';
   a_mod_56_port <= '0';
   a_mod_55_port <= '0';
   a_mod_54_port <= '0';
   a_mod_53_port <= '0';
   a_mod_52_port <= '0';
   a_mod_51_port <= '0';
   a_mod_50_port <= '0';
   a_mod_49_port <= '0';
   a_mod_48_port <= '0';
   a_mod_47_port <= '0';
   a_mod_46_port <= '0';
   a_mod_45_port <= '0';
   a_mod_44_port <= '0';
   a_mod_43_port <= '0';
   a_mod_42_port <= '0';
   a_mod_41_port <= '0';
   a_mod_40_port <= '0';
   a_mod_39_port <= '0';
   a_mod_38_port <= '0';
   a_mod_37_port <= '0';
   a_mod_36_port <= '0';
   a_mod_35_port <= '0';
   a_mod_34_port <= '0';
   a_mod_33_port <= '0';
   a_mod_32_port <= '0';
   ADJUST0a : AddSub_DATA_SIZE32_0 port map( as => n141, a(31) => X_Logic0_port
                           , a(30) => X_Logic0_port, a(29) => X_Logic0_port, 
                           a(28) => X_Logic0_port, a(27) => X_Logic0_port, 
                           a(26) => X_Logic0_port, a(25) => X_Logic0_port, 
                           a(24) => X_Logic0_port, a(23) => X_Logic0_port, 
                           a(22) => X_Logic0_port, a(21) => X_Logic0_port, 
                           a(20) => X_Logic0_port, a(19) => X_Logic0_port, 
                           a(18) => X_Logic0_port, a(17) => X_Logic0_port, 
                           a(16) => X_Logic0_port, a(15) => X_Logic0_port, 
                           a(14) => X_Logic0_port, a(13) => X_Logic0_port, 
                           a(12) => X_Logic0_port, a(11) => X_Logic0_port, 
                           a(10) => X_Logic0_port, a(9) => X_Logic0_port, a(8) 
                           => X_Logic0_port, a(7) => X_Logic0_port, a(6) => 
                           X_Logic0_port, a(5) => X_Logic0_port, a(4) => 
                           X_Logic0_port, a(3) => X_Logic0_port, a(2) => 
                           X_Logic0_port, a(1) => X_Logic0_port, a(0) => 
                           X_Logic0_port, b(31) => a(31), b(30) => a(30), b(29)
                           => a(29), b(28) => a(28), b(27) => a(27), b(26) => 
                           a(26), b(25) => a(25), b(24) => a(24), b(23) => 
                           a(23), b(22) => a(22), b(21) => a(21), b(20) => 
                           a(20), b(19) => a(19), b(18) => a(18), b(17) => 
                           a(17), b(16) => a(16), b(15) => a(15), b(14) => 
                           a(14), b(13) => a(13), b(12) => a(12), b(11) => 
                           a(11), b(10) => a(10), b(9) => a(9), b(8) => a(8), 
                           b(7) => a(7), b(6) => a(6), b(5) => a(5), b(4) => 
                           a(4), b(3) => a(3), b(2) => a(2), b(1) => a(1), b(0)
                           => a(0), re(31) => a_adj_31_port, re(30) => 
                           a_adj_30_port, re(29) => a_adj_29_port, re(28) => 
                           a_adj_28_port, re(27) => a_adj_27_port, re(26) => 
                           a_adj_26_port, re(25) => a_adj_25_port, re(24) => 
                           a_adj_24_port, re(23) => a_adj_23_port, re(22) => 
                           a_adj_22_port, re(21) => a_adj_21_port, re(20) => 
                           a_adj_20_port, re(19) => a_adj_19_port, re(18) => 
                           a_adj_18_port, re(17) => a_adj_17_port, re(16) => 
                           a_adj_16_port, re(15) => a_adj_15_port, re(14) => 
                           a_adj_14_port, re(13) => a_adj_13_port, re(12) => 
                           a_adj_12_port, re(11) => a_adj_11_port, re(10) => 
                           a_adj_10_port, re(9) => a_adj_9_port, re(8) => 
                           a_adj_8_port, re(7) => a_adj_7_port, re(6) => 
                           a_adj_6_port, re(5) => a_adj_5_port, re(4) => 
                           a_adj_4_port, re(3) => a_adj_3_port, re(2) => 
                           a_adj_2_port, re(1) => a_adj_1_port, re(0) => 
                           a_adj_0_port, cout => net3930);
   ADJUST0b : AddSub_DATA_SIZE32_3 port map( as => n145, a(31) => X_Logic0_port
                           , a(30) => X_Logic0_port, a(29) => X_Logic0_port, 
                           a(28) => X_Logic0_port, a(27) => X_Logic0_port, 
                           a(26) => X_Logic0_port, a(25) => X_Logic0_port, 
                           a(24) => X_Logic0_port, a(23) => X_Logic0_port, 
                           a(22) => X_Logic0_port, a(21) => X_Logic0_port, 
                           a(20) => X_Logic0_port, a(19) => X_Logic0_port, 
                           a(18) => X_Logic0_port, a(17) => X_Logic0_port, 
                           a(16) => X_Logic0_port, a(15) => X_Logic0_port, 
                           a(14) => X_Logic0_port, a(13) => X_Logic0_port, 
                           a(12) => X_Logic0_port, a(11) => X_Logic0_port, 
                           a(10) => X_Logic0_port, a(9) => X_Logic0_port, a(8) 
                           => X_Logic0_port, a(7) => X_Logic0_port, a(6) => 
                           X_Logic0_port, a(5) => X_Logic0_port, a(4) => 
                           X_Logic0_port, a(3) => X_Logic0_port, a(2) => 
                           X_Logic0_port, a(1) => X_Logic0_port, a(0) => 
                           X_Logic0_port, b(31) => b(31), b(30) => b(30), b(29)
                           => b(29), b(28) => b(28), b(27) => b(27), b(26) => 
                           b(26), b(25) => b(25), b(24) => b(24), b(23) => 
                           b(23), b(22) => b(22), b(21) => b(21), b(20) => 
                           b(20), b(19) => b(19), b(18) => b(18), b(17) => 
                           b(17), b(16) => b(16), b(15) => b(15), b(14) => 
                           b(14), b(13) => b(13), b(12) => b(12), b(11) => 
                           b(11), b(10) => b(10), b(9) => b(9), b(8) => b(8), 
                           b(7) => b(7), b(6) => b(6), b(5) => b(5), b(4) => 
                           b(4), b(3) => b(3), b(2) => b(2), b(1) => b(1), b(0)
                           => b(0), re(31) => b_adj_31_port, re(30) => 
                           b_adj_30_port, re(29) => b_adj_29_port, re(28) => 
                           b_adj_28_port, re(27) => b_adj_27_port, re(26) => 
                           b_adj_26_port, re(25) => b_adj_25_port, re(24) => 
                           b_adj_24_port, re(23) => b_adj_23_port, re(22) => 
                           b_adj_22_port, re(21) => b_adj_21_port, re(20) => 
                           b_adj_20_port, re(19) => b_adj_19_port, re(18) => 
                           b_adj_18_port, re(17) => b_adj_17_port, re(16) => 
                           b_adj_16_port, re(15) => b_adj_15_port, re(14) => 
                           b_adj_14_port, re(13) => b_adj_13_port, re(12) => 
                           b_adj_12_port, re(11) => b_adj_11_port, re(10) => 
                           b_adj_10_port, re(9) => b_adj_9_port, re(8) => 
                           b_adj_8_port, re(7) => b_adj_7_port, re(6) => 
                           b_adj_6_port, re(5) => b_adj_5_port, re(4) => 
                           b_adj_4_port, re(3) => b_adj_3_port, re(2) => 
                           b_adj_2_port, re(1) => b_adj_1_port, re(0) => 
                           b_adj_0_port, cout => net3929);
   MUXa : Mux_DATA_SIZE64 port map( sel => n149, din0(63) => a_mod_63_port, 
                           din0(62) => a_mod_62_port, din0(61) => a_mod_61_port
                           , din0(60) => a_mod_60_port, din0(59) => 
                           a_mod_59_port, din0(58) => a_mod_58_port, din0(57) 
                           => a_mod_57_port, din0(56) => a_mod_56_port, 
                           din0(55) => a_mod_55_port, din0(54) => a_mod_54_port
                           , din0(53) => a_mod_53_port, din0(52) => 
                           a_mod_52_port, din0(51) => a_mod_51_port, din0(50) 
                           => a_mod_50_port, din0(49) => a_mod_49_port, 
                           din0(48) => a_mod_48_port, din0(47) => a_mod_47_port
                           , din0(46) => a_mod_46_port, din0(45) => 
                           a_mod_45_port, din0(44) => a_mod_44_port, din0(43) 
                           => a_mod_43_port, din0(42) => a_mod_42_port, 
                           din0(41) => a_mod_41_port, din0(40) => a_mod_40_port
                           , din0(39) => a_mod_39_port, din0(38) => 
                           a_mod_38_port, din0(37) => a_mod_37_port, din0(36) 
                           => a_mod_36_port, din0(35) => a_mod_35_port, 
                           din0(34) => a_mod_34_port, din0(33) => a_mod_33_port
                           , din0(32) => a_mod_32_port, din0(31) => n218, 
                           din0(30) => n219, din0(29) => n220, din0(28) => n221
                           , din0(27) => a_mod_27_port, din0(26) => 
                           a_mod_26_port, din0(25) => a_mod_25_port, din0(24) 
                           => a_mod_24_port, din0(23) => a_mod_23_port, 
                           din0(22) => a_mod_22_port, din0(21) => a_mod_21_port
                           , din0(20) => a_mod_20_port, din0(19) => 
                           a_mod_19_port, din0(18) => a_mod_18_port, din0(17) 
                           => a_mod_17_port, din0(16) => a_mod_16_port, 
                           din0(15) => a_mod_15_port, din0(14) => a_mod_14_port
                           , din0(13) => a_mod_13_port, din0(12) => 
                           a_mod_12_port, din0(11) => a_mod_11_port, din0(10) 
                           => a_mod_10_port, din0(9) => a_mod_9_port, din0(8) 
                           => a_mod_8_port, din0(7) => a_mod_7_port, din0(6) =>
                           a_mod_6_port, din0(5) => a_mod_5_port, din0(4) => 
                           a_mod_4_port, din0(3) => a_mod_3_port, din0(2) => 
                           a_mod_2_port, din0(1) => a_mod_1_port, din0(0) => 
                           a_mod_0_port, din1(63) => r_63_port, din1(62) => 
                           r_62_port, din1(61) => r_61_port, din1(60) => 
                           r_60_port, din1(59) => r_59_port, din1(58) => 
                           r_58_port, din1(57) => r_57_port, din1(56) => 
                           r_56_port, din1(55) => r_55_port, din1(54) => 
                           r_54_port, din1(53) => r_53_port, din1(52) => 
                           r_52_port, din1(51) => r_51_port, din1(50) => 
                           r_50_port, din1(49) => r_49_port, din1(48) => 
                           r_48_port, din1(47) => r_47_port, din1(46) => 
                           r_46_port, din1(45) => r_45_port, din1(44) => 
                           r_44_port, din1(43) => r_43_port, din1(42) => 
                           r_42_port, din1(41) => r_41_port, din1(40) => 
                           r_40_port, din1(39) => r_39_port, din1(38) => 
                           r_38_port, din1(37) => r_37_port, din1(36) => 
                           r_36_port, din1(35) => r_35_port, din1(34) => 
                           r_34_port, din1(33) => r_33_port, din1(32) => 
                           r_32_port, din1(31) => r_31_port, din1(30) => 
                           r_30_port, din1(29) => r_29_port, din1(28) => 
                           r_28_port, din1(27) => r_27_port, din1(26) => 
                           r_26_port, din1(25) => r_25_port, din1(24) => 
                           r_24_port, din1(23) => r_23_port, din1(22) => 
                           r_22_port, din1(21) => r_21_port, din1(20) => 
                           r_20_port, din1(19) => r_19_port, din1(18) => 
                           r_18_port, din1(17) => r_17_port, din1(16) => 
                           r_16_port, din1(15) => r_15_port, din1(14) => 
                           r_14_port, din1(13) => r_13_port, din1(12) => 
                           r_12_port, din1(11) => r_11_port, din1(10) => 
                           r_10_port, din1(9) => r_9_port, din1(8) => r_8_port,
                           din1(7) => r_7_port, din1(6) => r_6_port, din1(5) =>
                           r_5_port, din1(4) => r_4_port, din1(3) => r_3_port, 
                           din1(2) => r_2_port, din1(1) => r_1_port, din1(0) =>
                           r_0_port, dout(63) => a_mux_63_port, dout(62) => 
                           a_mux_62_port, dout(61) => a_mux_61_port, dout(60) 
                           => a_mux_60_port, dout(59) => a_mux_59_port, 
                           dout(58) => a_mux_58_port, dout(57) => a_mux_57_port
                           , dout(56) => a_mux_56_port, dout(55) => 
                           a_mux_55_port, dout(54) => a_mux_54_port, dout(53) 
                           => a_mux_53_port, dout(52) => a_mux_52_port, 
                           dout(51) => a_mux_51_port, dout(50) => a_mux_50_port
                           , dout(49) => a_mux_49_port, dout(48) => 
                           a_mux_48_port, dout(47) => a_mux_47_port, dout(46) 
                           => a_mux_46_port, dout(45) => a_mux_45_port, 
                           dout(44) => a_mux_44_port, dout(43) => a_mux_43_port
                           , dout(42) => a_mux_42_port, dout(41) => 
                           a_mux_41_port, dout(40) => a_mux_40_port, dout(39) 
                           => a_mux_39_port, dout(38) => a_mux_38_port, 
                           dout(37) => a_mux_37_port, dout(36) => a_mux_36_port
                           , dout(35) => a_mux_35_port, dout(34) => 
                           a_mux_34_port, dout(33) => a_mux_33_port, dout(32) 
                           => a_mux_32_port, dout(31) => a_mux_31_port, 
                           dout(30) => a_mux_30_port, dout(29) => a_mux_29_port
                           , dout(28) => a_mux_28_port, dout(27) => 
                           a_mux_27_port, dout(26) => a_mux_26_port, dout(25) 
                           => a_mux_25_port, dout(24) => a_mux_24_port, 
                           dout(23) => a_mux_23_port, dout(22) => a_mux_22_port
                           , dout(21) => a_mux_21_port, dout(20) => 
                           a_mux_20_port, dout(19) => a_mux_19_port, dout(18) 
                           => a_mux_18_port, dout(17) => a_mux_17_port, 
                           dout(16) => a_mux_16_port, dout(15) => a_mux_15_port
                           , dout(14) => a_mux_14_port, dout(13) => 
                           a_mux_13_port, dout(12) => a_mux_12_port, dout(11) 
                           => a_mux_11_port, dout(10) => a_mux_10_port, dout(9)
                           => a_mux_9_port, dout(8) => a_mux_8_port, dout(7) =>
                           a_mux_7_port, dout(6) => a_mux_6_port, dout(5) => 
                           a_mux_5_port, dout(4) => a_mux_4_port, dout(3) => 
                           a_mux_3_port, dout(2) => a_mux_2_port, dout(1) => 
                           a_mux_1_port, dout(0) => a_mux_0_port);
   ADD0 : AddSub_DATA_SIZE64 port map( as => not_r_sign, a(63) => n260, a(62) 
                           => n261, a(61) => n262, a(60) => n263, a(59) => n264
                           , a(58) => n265, a(57) => n266, a(56) => n267, a(55)
                           => n268, a(54) => n269, a(53) => n270, a(52) => n271
                           , a(51) => n272, a(50) => n273, a(49) => n274, a(48)
                           => n275, a(47) => n276, a(46) => n277, a(45) => n278
                           , a(44) => n279, a(43) => n280, a(42) => n281, a(41)
                           => n282, a(40) => n283, a(39) => n284, a(38) => n285
                           , a(37) => n286, a(36) => n287, a(35) => n288, a(34)
                           => n289, a(33) => n290, a(32) => n291, a(31) => n292
                           , a(30) => n293, a(29) => n294, a(28) => n295, a(27)
                           => n296, a(26) => n363, a(25) => n364, a(24) => n365
                           , a(23) => n366, a(22) => n367, a(21) => n368, a(20)
                           => n369, a(19) => n370, a(18) => n371, a(17) => n375
                           , a(16) => n376, a(15) => n377, a(14) => n378, a(13)
                           => n379, a(12) => n380, a(11) => n381, a(10) => n382
                           , a(9) => n383, a(8) => n384, a(7) => n385, a(6) => 
                           n386, a(5) => n387, a(4) => n388, a(3) => n389, a(2)
                           => n390, a(1) => a_shf_1_port, a(0) => X_Logic0_port
                           , b(63) => b_shf_63_port, b(62) => b_shf_62_port, 
                           b(61) => b_shf_61_port, b(60) => b_shf_60_port, 
                           b(59) => b_shf_59_port, b(58) => b_shf_58_port, 
                           b(57) => b_shf_57_port, b(56) => b_shf_56_port, 
                           b(55) => b_shf_55_port, b(54) => b_shf_54_port, 
                           b(53) => b_shf_53_port, b(52) => b_shf_52_port, 
                           b(51) => b_shf_51_port, b(50) => b_shf_50_port, 
                           b(49) => b_shf_49_port, b(48) => b_shf_48_port, 
                           b(47) => b_shf_47_port, b(46) => b_shf_46_port, 
                           b(45) => b_shf_45_port, b(44) => b_shf_44_port, 
                           b(43) => b_shf_43_port, b(42) => b_shf_42_port, 
                           b(41) => b_shf_41_port, b(40) => b_shf_40_port, 
                           b(39) => b_shf_39_port, b(38) => b_shf_38_port, 
                           b(37) => b_shf_37_port, b(36) => b_shf_36_port, 
                           b(35) => b_shf_35_port, b(34) => b_shf_34_port, 
                           b(33) => b_shf_33_port, b(32) => b_shf_32_port, 
                           b(31) => b_shf_31_port, b(30) => b_shf_30_port, 
                           b(29) => b_shf_29_port, b(28) => b_shf_28_port, 
                           b(27) => b_shf_27_port, b(26) => b_shf_26_port, 
                           b(25) => b_shf_25_port, b(24) => b_shf_24_port, 
                           b(23) => b_shf_23_port, b(22) => b_shf_22_port, 
                           b(21) => b_shf_21_port, b(20) => b_shf_20_port, 
                           b(19) => b_shf_19_port, b(18) => b_shf_18_port, 
                           b(17) => b_shf_17_port, b(16) => b_shf_16_port, 
                           b(15) => b_shf_15_port, b(14) => b_shf_14_port, 
                           b(13) => b_shf_13_port, b(12) => b_shf_12_port, 
                           b(11) => b_shf_11_port, b(10) => b_shf_10_port, b(9)
                           => b_shf_9_port, b(8) => b_shf_8_port, b(7) => 
                           b_shf_7_port, b(6) => b_shf_6_port, b(5) => 
                           b_shf_5_port, b(4) => b_shf_4_port, b(3) => 
                           b_shf_3_port, b(2) => b_shf_2_port, b(1) => 
                           b_shf_1_port, b(0) => b_shf_0_port, re(63) => 
                           r_es_63_port, re(62) => r_es_62_port, re(61) => 
                           r_es_61_port, re(60) => r_es_60_port, re(59) => 
                           r_es_59_port, re(58) => r_es_58_port, re(57) => 
                           r_es_57_port, re(56) => r_es_56_port, re(55) => 
                           r_es_55_port, re(54) => r_es_54_port, re(53) => 
                           r_es_53_port, re(52) => r_es_52_port, re(51) => 
                           r_es_51_port, re(50) => r_es_50_port, re(49) => 
                           r_es_49_port, re(48) => r_es_48_port, re(47) => 
                           r_es_47_port, re(46) => r_es_46_port, re(45) => 
                           r_es_45_port, re(44) => r_es_44_port, re(43) => 
                           r_es_43_port, re(42) => r_es_42_port, re(41) => 
                           r_es_41_port, re(40) => r_es_40_port, re(39) => 
                           r_es_39_port, re(38) => r_es_38_port, re(37) => 
                           r_es_37_port, re(36) => r_es_36_port, re(35) => 
                           r_es_35_port, re(34) => r_es_34_port, re(33) => 
                           r_es_33_port, re(32) => r_es_32_port, re(31) => 
                           r_es_31_port, re(30) => r_es_30_port, re(29) => 
                           r_es_29_port, re(28) => r_es_28_port, re(27) => 
                           r_es_27_port, re(26) => r_es_26_port, re(25) => 
                           r_es_25_port, re(24) => r_es_24_port, re(23) => 
                           r_es_23_port, re(22) => r_es_22_port, re(21) => 
                           r_es_21_port, re(20) => r_es_20_port, re(19) => 
                           r_es_19_port, re(18) => r_es_18_port, re(17) => 
                           r_es_17_port, re(16) => r_es_16_port, re(15) => 
                           r_es_15_port, re(14) => r_es_14_port, re(13) => 
                           r_es_13_port, re(12) => r_es_12_port, re(11) => 
                           r_es_11_port, re(10) => r_es_10_port, re(9) => 
                           r_es_9_port, re(8) => r_es_8_port, re(7) => 
                           r_es_7_port, re(6) => r_es_6_port, re(5) => 
                           r_es_5_port, re(4) => r_es_4_port, re(3) => 
                           r_es_3_port, re(2) => r_es_2_port, re(1) => 
                           r_es_1_port, re(0) => r_es_0_port, cout => net3928);
   REG_R : Reg_DATA_SIZE64 port map( rst => n152, en => n163, clk => clk, 
                           din(63) => r_es_63_port, din(62) => r_es_62_port, 
                           din(61) => r_es_61_port, din(60) => r_es_60_port, 
                           din(59) => r_es_59_port, din(58) => r_es_58_port, 
                           din(57) => r_es_57_port, din(56) => r_es_56_port, 
                           din(55) => r_es_55_port, din(54) => r_es_54_port, 
                           din(53) => r_es_53_port, din(52) => r_es_52_port, 
                           din(51) => r_es_51_port, din(50) => r_es_50_port, 
                           din(49) => r_es_49_port, din(48) => r_es_48_port, 
                           din(47) => r_es_47_port, din(46) => r_es_46_port, 
                           din(45) => r_es_45_port, din(44) => r_es_44_port, 
                           din(43) => r_es_43_port, din(42) => r_es_42_port, 
                           din(41) => r_es_41_port, din(40) => r_es_40_port, 
                           din(39) => r_es_39_port, din(38) => r_es_38_port, 
                           din(37) => r_es_37_port, din(36) => r_es_36_port, 
                           din(35) => r_es_35_port, din(34) => r_es_34_port, 
                           din(33) => r_es_33_port, din(32) => r_es_32_port, 
                           din(31) => r_es_31_port, din(30) => r_es_30_port, 
                           din(29) => r_es_29_port, din(28) => r_es_28_port, 
                           din(27) => r_es_27_port, din(26) => r_es_26_port, 
                           din(25) => r_es_25_port, din(24) => r_es_24_port, 
                           din(23) => r_es_23_port, din(22) => r_es_22_port, 
                           din(21) => r_es_21_port, din(20) => r_es_20_port, 
                           din(19) => r_es_19_port, din(18) => r_es_18_port, 
                           din(17) => r_es_17_port, din(16) => r_es_16_port, 
                           din(15) => r_es_15_port, din(14) => r_es_14_port, 
                           din(13) => r_es_13_port, din(12) => r_es_12_port, 
                           din(11) => r_es_11_port, din(10) => r_es_10_port, 
                           din(9) => r_es_9_port, din(8) => r_es_8_port, din(7)
                           => r_es_7_port, din(6) => r_es_6_port, din(5) => 
                           r_es_5_port, din(4) => r_es_4_port, din(3) => 
                           r_es_3_port, din(2) => r_es_2_port, din(1) => 
                           r_es_1_port, din(0) => r_es_0_port, dout(63) => 
                           r_63_port, dout(62) => r_62_port, dout(61) => 
                           r_61_port, dout(60) => r_60_port, dout(59) => 
                           r_59_port, dout(58) => r_58_port, dout(57) => 
                           r_57_port, dout(56) => r_56_port, dout(55) => 
                           r_55_port, dout(54) => r_54_port, dout(53) => 
                           r_53_port, dout(52) => r_52_port, dout(51) => 
                           r_51_port, dout(50) => r_50_port, dout(49) => 
                           r_49_port, dout(48) => r_48_port, dout(47) => 
                           r_47_port, dout(46) => r_46_port, dout(45) => 
                           r_45_port, dout(44) => r_44_port, dout(43) => 
                           r_43_port, dout(42) => r_42_port, dout(41) => 
                           r_41_port, dout(40) => r_40_port, dout(39) => 
                           r_39_port, dout(38) => r_38_port, dout(37) => 
                           r_37_port, dout(36) => r_36_port, dout(35) => 
                           r_35_port, dout(34) => r_34_port, dout(33) => 
                           r_33_port, dout(32) => r_32_port, dout(31) => 
                           r_31_port, dout(30) => r_30_port, dout(29) => 
                           r_29_port, dout(28) => r_28_port, dout(27) => 
                           r_27_port, dout(26) => r_26_port, dout(25) => 
                           r_25_port, dout(24) => r_24_port, dout(23) => 
                           r_23_port, dout(22) => r_22_port, dout(21) => 
                           r_21_port, dout(20) => r_20_port, dout(19) => 
                           r_19_port, dout(18) => r_18_port, dout(17) => 
                           r_17_port, dout(16) => r_16_port, dout(15) => 
                           r_15_port, dout(14) => r_14_port, dout(13) => 
                           r_13_port, dout(12) => r_12_port, dout(11) => 
                           r_11_port, dout(10) => r_10_port, dout(9) => 
                           r_9_port, dout(8) => r_8_port, dout(7) => r_7_port, 
                           dout(6) => r_6_port, dout(5) => r_5_port, dout(4) =>
                           r_4_port, dout(3) => r_3_port, dout(2) => r_2_port, 
                           dout(1) => r_1_port, dout(0) => r_0_port);
   REG_Q : Sipo_DATA_SIZE32 port map( rst => n152, en => n163, clk => clk, din 
                           => not_r_es_sign, dout(31) => q_31_port, dout(30) =>
                           q_30_port, dout(29) => b_shf_sqrt_63_port, dout(28) 
                           => b_shf_sqrt_62_port, dout(27) => 
                           b_shf_sqrt_61_port, dout(26) => b_shf_sqrt_60_port, 
                           dout(25) => b_shf_sqrt_59_port, dout(24) => 
                           b_shf_sqrt_58_port, dout(23) => b_shf_sqrt_57_port, 
                           dout(22) => b_shf_sqrt_56_port, dout(21) => 
                           b_shf_sqrt_55_port, dout(20) => b_shf_sqrt_54_port, 
                           dout(19) => b_shf_sqrt_53_port, dout(18) => 
                           b_shf_sqrt_52_port, dout(17) => b_shf_sqrt_51_port, 
                           dout(16) => b_shf_sqrt_50_port, dout(15) => 
                           b_shf_sqrt_49_port, dout(14) => b_shf_sqrt_48_port, 
                           dout(13) => b_shf_sqrt_47_port, dout(12) => 
                           b_shf_sqrt_46_port, dout(11) => b_shf_sqrt_45_port, 
                           dout(10) => b_shf_sqrt_44_port, dout(9) => 
                           b_shf_sqrt_43_port, dout(8) => b_shf_sqrt_42_port, 
                           dout(7) => b_shf_sqrt_41_port, dout(6) => 
                           b_shf_sqrt_40_port, dout(5) => b_shf_sqrt_39_port, 
                           dout(4) => b_shf_sqrt_38_port, dout(3) => 
                           b_shf_sqrt_37_port, dout(2) => b_shf_sqrt_36_port, 
                           dout(1) => b_shf_sqrt_35_port, dout(0) => 
                           b_shf_sqrt_34_port);
   ADJUST : AddSub_DATA_SIZE32_2 port map( as => n213, a(31) => X_Logic0_port, 
                           a(30) => X_Logic0_port, a(29) => X_Logic0_port, 
                           a(28) => X_Logic0_port, a(27) => X_Logic0_port, 
                           a(26) => X_Logic0_port, a(25) => X_Logic0_port, 
                           a(24) => X_Logic0_port, a(23) => X_Logic0_port, 
                           a(22) => X_Logic0_port, a(21) => X_Logic0_port, 
                           a(20) => X_Logic0_port, a(19) => X_Logic0_port, 
                           a(18) => X_Logic0_port, a(17) => X_Logic0_port, 
                           a(16) => X_Logic0_port, a(15) => X_Logic0_port, 
                           a(14) => X_Logic0_port, a(13) => X_Logic0_port, 
                           a(12) => X_Logic0_port, a(11) => X_Logic0_port, 
                           a(10) => X_Logic0_port, a(9) => X_Logic0_port, a(8) 
                           => X_Logic0_port, a(7) => X_Logic0_port, a(6) => 
                           X_Logic0_port, a(5) => X_Logic0_port, a(4) => 
                           X_Logic0_port, a(3) => X_Logic0_port, a(2) => 
                           X_Logic0_port, a(1) => X_Logic0_port, a(0) => 
                           X_Logic0_port, b(31) => q_31_port, b(30) => 
                           q_30_port, b(29) => b_shf_sqrt_63_port, b(28) => 
                           b_shf_sqrt_62_port, b(27) => b_shf_sqrt_61_port, 
                           b(26) => b_shf_sqrt_60_port, b(25) => 
                           b_shf_sqrt_59_port, b(24) => b_shf_sqrt_58_port, 
                           b(23) => b_shf_sqrt_57_port, b(22) => 
                           b_shf_sqrt_56_port, b(21) => b_shf_sqrt_55_port, 
                           b(20) => b_shf_sqrt_54_port, b(19) => 
                           b_shf_sqrt_53_port, b(18) => b_shf_sqrt_52_port, 
                           b(17) => b_shf_sqrt_51_port, b(16) => 
                           b_shf_sqrt_50_port, b(15) => b_shf_sqrt_49_port, 
                           b(14) => b_shf_sqrt_48_port, b(13) => 
                           b_shf_sqrt_47_port, b(12) => b_shf_sqrt_46_port, 
                           b(11) => b_shf_sqrt_45_port, b(10) => 
                           b_shf_sqrt_44_port, b(9) => b_shf_sqrt_43_port, b(8)
                           => b_shf_sqrt_42_port, b(7) => b_shf_sqrt_41_port, 
                           b(6) => b_shf_sqrt_40_port, b(5) => 
                           b_shf_sqrt_39_port, b(4) => b_shf_sqrt_38_port, b(3)
                           => b_shf_sqrt_37_port, b(2) => b_shf_sqrt_36_port, 
                           b(1) => b_shf_sqrt_35_port, b(0) => 
                           b_shf_sqrt_34_port, re(31) => o(31), re(30) => o(30)
                           , re(29) => o(29), re(28) => o(28), re(27) => o(27),
                           re(26) => o(26), re(25) => o(25), re(24) => o(24), 
                           re(23) => o(23), re(22) => o(22), re(21) => o(21), 
                           re(20) => o(20), re(19) => o(19), re(18) => o(18), 
                           re(17) => o(17), re(16) => o(16), re(15) => o(15), 
                           re(14) => o(14), re(13) => o(13), re(12) => o(12), 
                           re(11) => o(11), re(10) => o(10), re(9) => o(9), 
                           re(8) => o(8), re(7) => o(7), re(6) => o(6), re(5) 
                           => o(5), re(4) => o(4), re(3) => o(3), re(2) => o(2)
                           , re(1) => o(1), re(0) => o(0), cout => net3927);
   add_197 : Div_DATA_SIZE32_DIV_STAGE34_SQRT_STAGE18_DW01_inc_0 port map( 
                           A(31) => c_state_31_port, A(30) => n180, A(29) => 
                           c_state_29_port, A(28) => c_state_28_port, A(27) => 
                           c_state_27_port, A(26) => c_state_26_port, A(25) => 
                           n178, A(24) => c_state_24_port, A(23) => 
                           c_state_23_port, A(22) => c_state_22_port, A(21) => 
                           c_state_21_port, A(20) => c_state_20_port, A(19) => 
                           c_state_19_port, A(18) => n186, A(17) => 
                           c_state_17_port, A(16) => c_state_16_port, A(15) => 
                           c_state_15_port, A(14) => c_state_14_port, A(13) => 
                           c_state_13_port, A(12) => c_state_12_port, A(11) => 
                           c_state_11_port, A(10) => c_state_10_port, A(9) => 
                           c_state_9_port, A(8) => c_state_8_port, A(7) => 
                           c_state_7_port, A(6) => c_state_6_port, A(5) => 
                           c_state_5_port, A(4) => c_state_4_port, A(3) => 
                           c_state_3_port, A(2) => c_state_2_port, A(1) => 
                           c_state_1_port, A(0) => c_state_0_port, SUM(31) => 
                           N48, SUM(30) => N47, SUM(29) => N46, SUM(28) => N45,
                           SUM(27) => N44, SUM(26) => N43, SUM(25) => N42, 
                           SUM(24) => N41, SUM(23) => N40, SUM(22) => N39, 
                           SUM(21) => N38, SUM(20) => N37, SUM(19) => N36, 
                           SUM(18) => N35, SUM(17) => N34, SUM(16) => N33, 
                           SUM(15) => N32, SUM(14) => N31, SUM(13) => N30, 
                           SUM(12) => N29, SUM(11) => N28, SUM(10) => N27, 
                           SUM(9) => N26, SUM(8) => N25, SUM(7) => N24, SUM(6) 
                           => N23, SUM(5) => N22, SUM(4) => N21, SUM(3) => N20,
                           SUM(2) => N19, SUM(1) => N18, SUM(0) => N17);
   inv_q_flag_mod_reg : DFF_X1 port map( D => n297, CK => clk, Q => n213, QN =>
                           n87);
   a_mod_reg_30_inst : DFF_X1 port map( D => n331, CK => clk, Q => n219, QN => 
                           n142);
   a_mod_reg_29_inst : DFF_X1 port map( D => n332, CK => clk, Q => n220, QN => 
                           n140);
   a_mod_reg_31_inst : DFF_X1 port map( D => n330, CK => clk, Q => n218, QN => 
                           n136);
   b_mod_reg_63_inst : DFF_X1 port map( D => n298, CK => clk, Q => n214, QN => 
                           net108616);
   b_mod_reg_62_inst : DFF_X1 port map( D => n299, CK => clk, Q => n215, QN => 
                           net108617);
   U3 : AND2_X1 port map( A1 => n134, A2 => n135, ZN => n190);
   U4 : MUX2_X1 port map( A => a_mux_1_port, B => a_mux_0_port, S => n168, Z =>
                           n390);
   U5 : BUF_X1 port map( A => n169, Z => n157);
   U6 : NAND2_X1 port map( A1 => n215, A2 => n163, ZN => n131);
   U7 : NAND2_X1 port map( A1 => n214, A2 => n163, ZN => n133);
   U8 : INV_X1 port map( A => n87, ZN => n88);
   U9 : OR2_X1 port map( A1 => n195, A2 => n193, ZN => n102);
   U10 : BUF_X1 port map( A => n391, Z => n163);
   U11 : NAND2_X1 port map( A1 => b_adj_30_port, A2 => n167, ZN => n130);
   U12 : NAND2_X1 port map( A1 => n130, A2 => n131, ZN => n299);
   U13 : NAND2_X1 port map( A1 => b_adj_31_port, A2 => n165, ZN => n132);
   U14 : NAND2_X1 port map( A1 => n132, A2 => n133, ZN => n298);
   U15 : AND3_X1 port map( A1 => sign, A2 => a(31), A3 => n171, ZN => n141);
   U16 : AND2_X1 port map( A1 => n183, A2 => n182, ZN => n134);
   U17 : AND2_X1 port map( A1 => n189, A2 => n188, ZN => n135);
   U18 : AND3_X2 port map( A1 => sign, A2 => b(31), A3 => n158, ZN => n145);
   U19 : MUX2_X1 port map( A => a_adj_28_port, B => n221, S => n164, Z => n333)
                           ;
   U20 : CLKBUF_X1 port map( A => n145, Z => n137);
   U21 : INV_X1 port map( A => n141, ZN => n210);
   U22 : CLKBUF_X1 port map( A => n149, Z => n138);
   U23 : INV_X1 port map( A => n137, ZN => n211);
   U24 : NAND3_X1 port map( A1 => n190, A2 => n191, A3 => n192, ZN => n139);
   U25 : MUX2_X1 port map( A => a_adj_31_port, B => n218, S => n164, Z => n330)
                           ;
   U26 : NAND2_X1 port map( A1 => b_adj_29_port, A2 => n166, ZN => n143);
   U27 : NAND2_X1 port map( A1 => n216, A2 => n163, ZN => n144);
   U28 : NAND2_X1 port map( A1 => n143, A2 => n144, ZN => n300);
   U29 : INV_X1 port map( A => n146, ZN => n147);
   U30 : INV_X2 port map( A => n159, ZN => n169);
   U31 : OAI21_X1 port map( B1 => c_state_4_port, B2 => n170, A => 
                           c_state_5_port, ZN => n148);
   U32 : INV_X1 port map( A => n138, ZN => n199);
   U33 : AND3_X2 port map( A1 => n197, A2 => n201, A3 => n204, ZN => n149);
   U34 : CLKBUF_X1 port map( A => n139, Z => n150);
   U35 : NOR2_X1 port map( A1 => n139, A2 => n102, ZN => n223);
   U36 : CLKBUF_X1 port map( A => n169, Z => n153);
   U37 : CLKBUF_X1 port map( A => n169, Z => n154);
   U38 : CLKBUF_X1 port map( A => n169, Z => n155);
   U39 : CLKBUF_X1 port map( A => n223, Z => n151);
   U40 : BUF_X2 port map( A => n169, Z => n156);
   U41 : INV_X1 port map( A => n164, ZN => n165);
   U42 : INV_X1 port map( A => n164, ZN => n166);
   U43 : INV_X1 port map( A => n164, ZN => n167);
   U44 : BUF_X1 port map( A => n258, Z => n160);
   U45 : BUF_X1 port map( A => n258, Z => n161);
   U46 : BUF_X1 port map( A => n258, Z => n162);
   U47 : AND2_X1 port map( A1 => n172, A2 => n163, ZN => n152);
   U48 : AND2_X1 port map( A1 => n171, A2 => a_mux_0_port, ZN => a_shf_1_port);
   U49 : AND2_X1 port map( A1 => N46, A2 => n160, ZN => n_state_29_port);
   U50 : AND2_X1 port map( A1 => N45, A2 => n160, ZN => n_state_28_port);
   U51 : AND2_X1 port map( A1 => N47, A2 => n160, ZN => n_state_30_port);
   U52 : AND2_X1 port map( A1 => N44, A2 => n161, ZN => n_state_27_port);
   U53 : AND2_X1 port map( A1 => N43, A2 => n161, ZN => n_state_26_port);
   U54 : AND2_X1 port map( A1 => N42, A2 => n161, ZN => n_state_25_port);
   U55 : AND2_X1 port map( A1 => N41, A2 => n161, ZN => n_state_24_port);
   U56 : AND2_X1 port map( A1 => N40, A2 => n161, ZN => n_state_23_port);
   U57 : AND2_X1 port map( A1 => N39, A2 => n161, ZN => n_state_22_port);
   U58 : BUF_X1 port map( A => rst, Z => n172);
   U59 : BUF_X1 port map( A => n391, Z => n164);
   U60 : AND2_X1 port map( A1 => N37, A2 => n161, ZN => n_state_20_port);
   U61 : AND2_X1 port map( A1 => N36, A2 => n161, ZN => n_state_19_port);
   U62 : AND2_X1 port map( A1 => N34, A2 => n161, ZN => n_state_17_port);
   U63 : AND2_X1 port map( A1 => N33, A2 => n162, ZN => n_state_16_port);
   U64 : AND2_X1 port map( A1 => N32, A2 => n162, ZN => n_state_15_port);
   U65 : AND2_X1 port map( A1 => N29, A2 => n162, ZN => n_state_12_port);
   U66 : AND2_X1 port map( A1 => N25, A2 => n160, ZN => n_state_8_port);
   U67 : AND2_X1 port map( A1 => N24, A2 => n160, ZN => n_state_7_port);
   U68 : AND2_X1 port map( A1 => N22, A2 => n160, ZN => n_state_5_port);
   U69 : AND2_X1 port map( A1 => N20, A2 => n160, ZN => n_state_3_port);
   U70 : AND2_X1 port map( A1 => N19, A2 => n160, ZN => n_state_2_port);
   U71 : AND2_X1 port map( A1 => N18, A2 => n161, ZN => n_state_1_port);
   U72 : AND2_X1 port map( A1 => N38, A2 => n161, ZN => n_state_21_port);
   U73 : AND2_X1 port map( A1 => N35, A2 => n161, ZN => n_state_18_port);
   U74 : AND2_X1 port map( A1 => N31, A2 => n162, ZN => n_state_14_port);
   U75 : AND2_X1 port map( A1 => N30, A2 => n162, ZN => n_state_13_port);
   U76 : AND2_X1 port map( A1 => N28, A2 => n162, ZN => n_state_11_port);
   U77 : AND2_X1 port map( A1 => N26, A2 => n160, ZN => n_state_9_port);
   U78 : AND2_X1 port map( A1 => N23, A2 => n160, ZN => n_state_6_port);
   U79 : AND2_X1 port map( A1 => N21, A2 => n160, ZN => n_state_4_port);
   U80 : AND2_X1 port map( A1 => N27, A2 => n162, ZN => n_state_10_port);
   U81 : BUF_X1 port map( A => rst, Z => n173);
   U82 : OAI21_X1 port map( B1 => net108644, B2 => n154, A => n252, ZN => 
                           b_shf_35_port);
   U83 : NAND2_X1 port map( A1 => b_shf_sqrt_35_port, A2 => n153, ZN => n252);
   U84 : OAI21_X1 port map( B1 => net108643, B2 => n154, A => n251, ZN => 
                           b_shf_36_port);
   U85 : NAND2_X1 port map( A1 => b_shf_sqrt_36_port, A2 => n153, ZN => n251);
   U86 : OAI21_X1 port map( B1 => net108619, B2 => n169, A => n227, ZN => 
                           b_shf_60_port);
   U87 : NAND2_X1 port map( A1 => b_shf_sqrt_60_port, A2 => n153, ZN => n227);
   U88 : NAND2_X1 port map( A1 => b_shf_sqrt_34_port, A2 => n153, ZN => n253);
   U89 : OAI21_X1 port map( B1 => net108642, B2 => n154, A => n250, ZN => 
                           b_shf_37_port);
   U90 : NAND2_X1 port map( A1 => b_shf_sqrt_37_port, A2 => n168, ZN => n250);
   U91 : OAI21_X1 port map( B1 => net108639, B2 => n169, A => n247, ZN => 
                           b_shf_40_port);
   U92 : NAND2_X1 port map( A1 => b_shf_sqrt_40_port, A2 => n168, ZN => n247);
   U93 : OAI21_X1 port map( B1 => net108634, B2 => n168, A => n242, ZN => 
                           b_shf_45_port);
   U94 : NAND2_X1 port map( A1 => b_shf_sqrt_45_port, A2 => n169, ZN => n242);
   U95 : OAI21_X1 port map( B1 => net108635, B2 => n169, A => n243, ZN => 
                           b_shf_44_port);
   U96 : NAND2_X1 port map( A1 => b_shf_sqrt_44_port, A2 => n154, ZN => n243);
   U97 : OAI21_X1 port map( B1 => net108631, B2 => n154, A => n239, ZN => 
                           b_shf_48_port);
   U98 : NAND2_X1 port map( A1 => b_shf_sqrt_48_port, A2 => n154, ZN => n239);
   U99 : OAI21_X1 port map( B1 => net108637, B2 => n155, A => n245, ZN => 
                           b_shf_42_port);
   U100 : NAND2_X1 port map( A1 => b_shf_sqrt_42_port, A2 => n154, ZN => n245);
   U101 : OAI21_X1 port map( B1 => net108629, B2 => n155, A => n237, ZN => 
                           b_shf_50_port);
   U102 : NAND2_X1 port map( A1 => b_shf_sqrt_50_port, A2 => n153, ZN => n237);
   U103 : OAI21_X1 port map( B1 => net108640, B2 => n154, A => n248, ZN => 
                           b_shf_39_port);
   U104 : NAND2_X1 port map( A1 => b_shf_sqrt_39_port, A2 => n168, ZN => n248);
   U105 : OAI21_X1 port map( B1 => net108636, B2 => n169, A => n244, ZN => 
                           b_shf_43_port);
   U106 : NAND2_X1 port map( A1 => b_shf_sqrt_43_port, A2 => n154, ZN => n244);
   U107 : OAI21_X1 port map( B1 => net108628, B2 => n154, A => n236, ZN => 
                           b_shf_51_port);
   U108 : NAND2_X1 port map( A1 => b_shf_sqrt_51_port, A2 => n153, ZN => n236);
   U109 : OAI21_X1 port map( B1 => net108627, B2 => n154, A => n235, ZN => 
                           b_shf_52_port);
   U110 : NAND2_X1 port map( A1 => b_shf_sqrt_52_port, A2 => n153, ZN => n235);
   U111 : OAI21_X1 port map( B1 => net108623, B2 => n169, A => n231, ZN => 
                           b_shf_56_port);
   U112 : NAND2_X1 port map( A1 => b_shf_sqrt_56_port, A2 => n168, ZN => n231);
   U113 : OAI21_X1 port map( B1 => net108633, B2 => n154, A => n241, ZN => 
                           b_shf_46_port);
   U114 : NAND2_X1 port map( A1 => b_shf_sqrt_46_port, A2 => n154, ZN => n241);
   U115 : OAI21_X1 port map( B1 => net108632, B2 => n168, A => n240, ZN => 
                           b_shf_47_port);
   U116 : NAND2_X1 port map( A1 => b_shf_sqrt_47_port, A2 => n168, ZN => n240);
   U117 : OAI21_X1 port map( B1 => net108638, B2 => n154, A => n246, ZN => 
                           b_shf_41_port);
   U118 : NAND2_X1 port map( A1 => b_shf_sqrt_41_port, A2 => n168, ZN => n246);
   U119 : OAI21_X1 port map( B1 => net108641, B2 => n154, A => n249, ZN => 
                           b_shf_38_port);
   U120 : NAND2_X1 port map( A1 => b_shf_sqrt_38_port, A2 => n153, ZN => n249);
   U121 : OAI21_X1 port map( B1 => net108630, B2 => n169, A => n238, ZN => 
                           b_shf_49_port);
   U122 : NAND2_X1 port map( A1 => b_shf_sqrt_49_port, A2 => n154, ZN => n238);
   U123 : NAND2_X1 port map( A1 => n76, A2 => n82, ZN => n193);
   U124 : OR2_X1 port map( A1 => n205, A2 => c_state_31_port, ZN => n196);
   U125 : OAI21_X1 port map( B1 => c_state_4_port, B2 => n170, A => 
                           c_state_5_port, ZN => n201);
   U126 : AND2_X1 port map( A1 => N48, A2 => n160, ZN => n_state_31_port);
   U127 : OAI21_X1 port map( B1 => net108618, B2 => n155, A => n226, ZN => 
                           b_shf_61_port);
   U128 : NAND2_X1 port map( A1 => b_shf_sqrt_61_port, A2 => n153, ZN => n226);
   U129 : OAI21_X1 port map( B1 => net108625, B2 => n154, A => n233, ZN => 
                           b_shf_54_port);
   U130 : NAND2_X1 port map( A1 => b_shf_sqrt_54_port, A2 => n169, ZN => n233);
   U131 : OAI21_X1 port map( B1 => net108621, B2 => n155, A => n229, ZN => 
                           b_shf_58_port);
   U132 : NAND2_X1 port map( A1 => b_shf_sqrt_58_port, A2 => n169, ZN => n229);
   U133 : OAI21_X1 port map( B1 => net108624, B2 => n169, A => n232, ZN => 
                           b_shf_55_port);
   U134 : NAND2_X1 port map( A1 => b_shf_sqrt_55_port, A2 => n168, ZN => n232);
   U135 : OAI21_X1 port map( B1 => net108626, B2 => n153, A => n234, ZN => 
                           b_shf_53_port);
   U136 : NAND2_X1 port map( A1 => b_shf_sqrt_53_port, A2 => n153, ZN => n234);
   U137 : OAI21_X1 port map( B1 => net108622, B2 => n154, A => n230, ZN => 
                           b_shf_57_port);
   U138 : NAND2_X1 port map( A1 => b_shf_sqrt_57_port, A2 => n153, ZN => n230);
   U139 : OAI21_X1 port map( B1 => net108616, B2 => n154, A => n224, ZN => 
                           b_shf_63_port);
   U140 : NAND2_X1 port map( A1 => b_shf_sqrt_63_port, A2 => n153, ZN => n224);
   U141 : OAI21_X1 port map( B1 => net108617, B2 => n168, A => n225, ZN => 
                           b_shf_62_port);
   U142 : NAND2_X1 port map( A1 => b_shf_sqrt_62_port, A2 => n153, ZN => n225);
   U143 : OAI21_X1 port map( B1 => net108620, B2 => n154, A => n228, ZN => 
                           b_shf_59_port);
   U144 : NAND2_X1 port map( A1 => b_shf_sqrt_59_port, A2 => n154, ZN => n228);
   U145 : AND2_X1 port map( A1 => c_state_0_port, A2 => n82, ZN => n202);
   U146 : OAI22_X1 port map( A1 => n257, A2 => n256, B1 => n255, B2 => n254, ZN
                           => n259);
   U147 : OAI21_X1 port map( B1 => n209, B2 => c_state_31_port, A => n208, ZN 
                           => n257);
   U148 : OAI21_X1 port map( B1 => n198, B2 => n362, A => n199, ZN => n391);
   U149 : INV_X1 port map( A => n168, ZN => n159);
   U150 : INV_X1 port map( A => func, ZN => n158);
   U151 : INV_X1 port map( A => func, ZN => n171);
   U152 : NAND2_X1 port map( A1 => func, A2 => c_state_4_port, ZN => n203);
   U153 : OAI21_X1 port map( B1 => net108645, B2 => n157, A => n253, ZN => 
                           b_shf_34_port);
   U154 : INV_X1 port map( A => n171, ZN => n168);
   U155 : INV_X1 port map( A => n158, ZN => n170);
   U156 : INV_X1 port map( A => r_es_63_port, ZN => not_r_es_sign);
   U157 : NAND3_X1 port map( A1 => n373, A2 => n77, A3 => n78, ZN => n195);
   U158 : NAND3_X1 port map( A1 => n98, A2 => n93, A3 => n89, ZN => n175);
   U159 : NAND3_X1 port map( A1 => n99, A2 => n94, A3 => n90, ZN => n174);
   U160 : NOR2_X1 port map( A1 => n175, A2 => n174, ZN => n192);
   U161 : NAND3_X1 port map( A1 => n100, A2 => n95, A3 => n91, ZN => n177);
   U162 : NAND3_X1 port map( A1 => n101, A2 => n96, A3 => n92, ZN => n176);
   U163 : NOR2_X1 port map( A1 => n177, A2 => n176, ZN => n191);
   U164 : NAND2_X1 port map( A1 => n372, A2 => n374, ZN => n179);
   U165 : NOR2_X1 port map( A1 => n179, A2 => n178, ZN => n183);
   U166 : NAND2_X1 port map( A1 => net108681, A2 => net108680, ZN => n181);
   U167 : NOR2_X1 port map( A1 => n181, A2 => n180, ZN => n182);
   U168 : NAND2_X1 port map( A1 => net108687, A2 => n73, ZN => n185);
   U169 : NAND2_X1 port map( A1 => n80, A2 => n81, ZN => n184);
   U170 : NOR2_X1 port map( A1 => n185, A2 => n184, ZN => n189);
   U171 : NAND2_X1 port map( A1 => net108686, A2 => net108685, ZN => n187);
   U172 : NOR2_X1 port map( A1 => n187, A2 => n147, ZN => n188);
   U173 : NAND3_X1 port map( A1 => n190, A2 => n191, A3 => n192, ZN => n205);
   U174 : NAND2_X1 port map( A1 => n72, A2 => n223, ZN => n198);
   U175 : NAND2_X1 port map( A1 => n82, A2 => n203, ZN => n194);
   U176 : NAND2_X1 port map( A1 => n195, A2 => n194, ZN => n204);
   U177 : NOR2_X1 port map( A1 => n196, A2 => n223, ZN => n197);
   U178 : NAND2_X1 port map( A1 => n71, A2 => n159, ZN => b_shf_32_port);
   U179 : MUX2_X1 port map( A => n97, B => a_mux_63_port, S => n155, Z => 
                           b_shf_33_port);
   U180 : MUX2_X1 port map( A => a_mux_2_port, B => a_mux_1_port, S => n169, Z 
                           => n389);
   U181 : MUX2_X1 port map( A => a_mux_3_port, B => a_mux_2_port, S => n169, Z 
                           => n388);
   U182 : MUX2_X1 port map( A => a_mux_4_port, B => a_mux_3_port, S => n169, Z 
                           => n387);
   U183 : MUX2_X1 port map( A => a_mux_5_port, B => a_mux_4_port, S => n168, Z 
                           => n386);
   U184 : MUX2_X1 port map( A => a_mux_6_port, B => a_mux_5_port, S => n168, Z 
                           => n385);
   U185 : MUX2_X1 port map( A => a_mux_7_port, B => a_mux_6_port, S => n157, Z 
                           => n384);
   U186 : MUX2_X1 port map( A => a_mux_8_port, B => a_mux_7_port, S => n157, Z 
                           => n383);
   U187 : MUX2_X1 port map( A => a_mux_9_port, B => a_mux_8_port, S => n157, Z 
                           => n382);
   U188 : MUX2_X1 port map( A => a_mux_10_port, B => a_mux_9_port, S => n156, Z
                           => n381);
   U189 : MUX2_X1 port map( A => a_mux_11_port, B => a_mux_10_port, S => n156, 
                           Z => n380);
   U190 : MUX2_X1 port map( A => a_mux_12_port, B => a_mux_11_port, S => n156, 
                           Z => n379);
   U191 : MUX2_X1 port map( A => a_mux_13_port, B => a_mux_12_port, S => n156, 
                           Z => n378);
   U192 : MUX2_X1 port map( A => a_mux_14_port, B => a_mux_13_port, S => n156, 
                           Z => n377);
   U193 : MUX2_X1 port map( A => a_mux_15_port, B => a_mux_14_port, S => n156, 
                           Z => n376);
   U194 : MUX2_X1 port map( A => a_mux_16_port, B => a_mux_15_port, S => n156, 
                           Z => n375);
   U195 : MUX2_X1 port map( A => a_mux_17_port, B => a_mux_16_port, S => n156, 
                           Z => n371);
   U196 : MUX2_X1 port map( A => a_mux_18_port, B => a_mux_17_port, S => n156, 
                           Z => n370);
   U197 : MUX2_X1 port map( A => a_mux_19_port, B => a_mux_18_port, S => n156, 
                           Z => n369);
   U198 : MUX2_X1 port map( A => a_mux_20_port, B => a_mux_19_port, S => n157, 
                           Z => n368);
   U199 : MUX2_X1 port map( A => a_mux_21_port, B => a_mux_20_port, S => n156, 
                           Z => n367);
   U200 : MUX2_X1 port map( A => a_mux_22_port, B => a_mux_21_port, S => n156, 
                           Z => n366);
   U201 : MUX2_X1 port map( A => a_mux_23_port, B => a_mux_22_port, S => n156, 
                           Z => n365);
   U202 : MUX2_X1 port map( A => a_mux_24_port, B => a_mux_23_port, S => n155, 
                           Z => n364);
   U203 : MUX2_X1 port map( A => a_mux_25_port, B => a_mux_24_port, S => n155, 
                           Z => n363);
   U204 : MUX2_X1 port map( A => a_mux_26_port, B => a_mux_25_port, S => n155, 
                           Z => n296);
   U205 : MUX2_X1 port map( A => a_mux_27_port, B => a_mux_26_port, S => n168, 
                           Z => n295);
   U206 : MUX2_X1 port map( A => a_mux_28_port, B => a_mux_27_port, S => n168, 
                           Z => n294);
   U207 : MUX2_X1 port map( A => a_mux_29_port, B => a_mux_28_port, S => n168, 
                           Z => n293);
   U208 : MUX2_X1 port map( A => a_mux_30_port, B => a_mux_29_port, S => n155, 
                           Z => n292);
   U209 : MUX2_X1 port map( A => a_mux_31_port, B => a_mux_30_port, S => n156, 
                           Z => n291);
   U210 : MUX2_X1 port map( A => a_mux_32_port, B => a_mux_31_port, S => n156, 
                           Z => n290);
   U211 : MUX2_X1 port map( A => a_mux_33_port, B => a_mux_32_port, S => n156, 
                           Z => n289);
   U212 : MUX2_X1 port map( A => a_mux_34_port, B => a_mux_33_port, S => n155, 
                           Z => n288);
   U213 : MUX2_X1 port map( A => a_mux_35_port, B => a_mux_34_port, S => n155, 
                           Z => n287);
   U214 : MUX2_X1 port map( A => a_mux_36_port, B => a_mux_35_port, S => n168, 
                           Z => n286);
   U215 : MUX2_X1 port map( A => a_mux_37_port, B => a_mux_36_port, S => n155, 
                           Z => n285);
   U216 : MUX2_X1 port map( A => a_mux_38_port, B => a_mux_37_port, S => n155, 
                           Z => n284);
   U217 : MUX2_X1 port map( A => a_mux_39_port, B => a_mux_38_port, S => n168, 
                           Z => n283);
   U218 : MUX2_X1 port map( A => a_mux_40_port, B => a_mux_39_port, S => n168, 
                           Z => n282);
   U219 : MUX2_X1 port map( A => a_mux_41_port, B => a_mux_40_port, S => n156, 
                           Z => n281);
   U220 : MUX2_X1 port map( A => a_mux_42_port, B => a_mux_41_port, S => n155, 
                           Z => n280);
   U221 : MUX2_X1 port map( A => a_mux_43_port, B => a_mux_42_port, S => n169, 
                           Z => n279);
   U222 : MUX2_X1 port map( A => a_mux_44_port, B => a_mux_43_port, S => n155, 
                           Z => n278);
   U223 : MUX2_X1 port map( A => a_mux_45_port, B => a_mux_44_port, S => n169, 
                           Z => n277);
   U224 : MUX2_X1 port map( A => a_mux_46_port, B => a_mux_45_port, S => n156, 
                           Z => n276);
   U225 : MUX2_X1 port map( A => a_mux_47_port, B => a_mux_46_port, S => n169, 
                           Z => n275);
   U226 : MUX2_X1 port map( A => a_mux_48_port, B => a_mux_47_port, S => n155, 
                           Z => n274);
   U227 : MUX2_X1 port map( A => a_mux_49_port, B => a_mux_48_port, S => n168, 
                           Z => n273);
   U228 : MUX2_X1 port map( A => a_mux_50_port, B => a_mux_49_port, S => n154, 
                           Z => n272);
   U229 : MUX2_X1 port map( A => a_mux_51_port, B => a_mux_50_port, S => n157, 
                           Z => n271);
   U230 : MUX2_X1 port map( A => a_mux_52_port, B => a_mux_51_port, S => n168, 
                           Z => n270);
   U231 : MUX2_X1 port map( A => a_mux_53_port, B => a_mux_52_port, S => n153, 
                           Z => n269);
   U232 : MUX2_X1 port map( A => a_mux_54_port, B => a_mux_53_port, S => n157, 
                           Z => n268);
   U233 : MUX2_X1 port map( A => a_mux_55_port, B => a_mux_54_port, S => n154, 
                           Z => n267);
   U234 : MUX2_X1 port map( A => a_mux_56_port, B => a_mux_55_port, S => n154, 
                           Z => n266);
   U235 : MUX2_X1 port map( A => a_mux_57_port, B => a_mux_56_port, S => n168, 
                           Z => n265);
   U236 : MUX2_X1 port map( A => a_mux_58_port, B => a_mux_57_port, S => n154, 
                           Z => n264);
   U237 : MUX2_X1 port map( A => a_mux_59_port, B => a_mux_58_port, S => n168, 
                           Z => n263);
   U238 : MUX2_X1 port map( A => a_mux_60_port, B => a_mux_59_port, S => n153, 
                           Z => n262);
   U239 : MUX2_X1 port map( A => a_mux_61_port, B => a_mux_60_port, S => n157, 
                           Z => n261);
   U240 : MUX2_X1 port map( A => a_mux_62_port, B => a_mux_61_port, S => n169, 
                           Z => n260);
   U241 : INV_X1 port map( A => a_mux_63_port, ZN => not_r_sign);
   U242 : NOR2_X1 port map( A1 => n151, A2 => c_state_0_port, ZN => n200);
   U243 : AOI22_X1 port map( A1 => n203, A2 => n202, B1 => n148, B2 => n200, ZN
                           => n207);
   U244 : INV_X1 port map( A => n204, ZN => n206);
   U245 : NOR3_X1 port map( A1 => n207, A2 => n206, A3 => n150, ZN => n209);
   U246 : NAND2_X1 port map( A1 => en, A2 => lock, ZN => n208);
   U247 : INV_X1 port map( A => n257, ZN => n258);
   U248 : OAI22_X1 port map( A1 => n211, A2 => a(31), B1 => n210, B2 => b(31), 
                           ZN => n212);
   U249 : MUX2_X1 port map( A => n88, B => n212, S => n165, Z => n297);
   U250 : MUX2_X1 port map( A => n217, B => b_adj_28_port, S => n166, Z => n301
                           );
   U251 : MUX2_X1 port map( A => n103, B => b_adj_27_port, S => n166, Z => n302
                           );
   U252 : MUX2_X1 port map( A => n104, B => b_adj_26_port, S => n167, Z => n303
                           );
   U253 : MUX2_X1 port map( A => n105, B => b_adj_25_port, S => n166, Z => n304
                           );
   U254 : MUX2_X1 port map( A => n106, B => b_adj_24_port, S => n165, Z => n305
                           );
   U255 : MUX2_X1 port map( A => n107, B => b_adj_23_port, S => n166, Z => n306
                           );
   U256 : MUX2_X1 port map( A => n108, B => b_adj_22_port, S => n167, Z => n307
                           );
   U257 : MUX2_X1 port map( A => n109, B => b_adj_21_port, S => n165, Z => n308
                           );
   U258 : MUX2_X1 port map( A => n110, B => b_adj_20_port, S => n167, Z => n309
                           );
   U259 : MUX2_X1 port map( A => n111, B => b_adj_19_port, S => n166, Z => n310
                           );
   U260 : MUX2_X1 port map( A => n112, B => b_adj_18_port, S => n165, Z => n311
                           );
   U261 : MUX2_X1 port map( A => n113, B => b_adj_17_port, S => n167, Z => n312
                           );
   U262 : MUX2_X1 port map( A => n114, B => b_adj_16_port, S => n166, Z => n313
                           );
   U263 : MUX2_X1 port map( A => n115, B => b_adj_15_port, S => n165, Z => n314
                           );
   U264 : MUX2_X1 port map( A => n116, B => b_adj_14_port, S => n167, Z => n315
                           );
   U265 : MUX2_X1 port map( A => n117, B => b_adj_13_port, S => n166, Z => n316
                           );
   U266 : MUX2_X1 port map( A => n118, B => b_adj_12_port, S => n165, Z => n317
                           );
   U267 : MUX2_X1 port map( A => n119, B => b_adj_11_port, S => n167, Z => n318
                           );
   U268 : MUX2_X1 port map( A => n120, B => b_adj_10_port, S => n166, Z => n319
                           );
   U269 : MUX2_X1 port map( A => n121, B => b_adj_9_port, S => n165, Z => n320)
                           ;
   U270 : MUX2_X1 port map( A => n122, B => b_adj_8_port, S => n165, Z => n321)
                           ;
   U271 : MUX2_X1 port map( A => n123, B => b_adj_7_port, S => n165, Z => n322)
                           ;
   U272 : MUX2_X1 port map( A => n124, B => b_adj_6_port, S => n165, Z => n323)
                           ;
   U273 : MUX2_X1 port map( A => n125, B => b_adj_5_port, S => n165, Z => n324)
                           ;
   U274 : MUX2_X1 port map( A => n126, B => b_adj_4_port, S => n165, Z => n325)
                           ;
   U275 : MUX2_X1 port map( A => n127, B => b_adj_3_port, S => n165, Z => n326)
                           ;
   U276 : MUX2_X1 port map( A => n128, B => b_adj_2_port, S => n165, Z => n327)
                           ;
   U277 : MUX2_X1 port map( A => n97, B => b_adj_1_port, S => n165, Z => n328);
   U278 : MUX2_X1 port map( A => n129, B => b_adj_0_port, S => n165, Z => n329)
                           ;
   U279 : MUX2_X1 port map( A => n219, B => a_adj_30_port, S => n165, Z => n331
                           );
   U280 : MUX2_X1 port map( A => n220, B => a_adj_29_port, S => n165, Z => n332
                           );
   U281 : MUX2_X1 port map( A => a_mod_27_port, B => a_adj_27_port, S => n166, 
                           Z => n334);
   U282 : MUX2_X1 port map( A => a_mod_26_port, B => a_adj_26_port, S => n166, 
                           Z => n335);
   U283 : MUX2_X1 port map( A => a_mod_25_port, B => a_adj_25_port, S => n166, 
                           Z => n336);
   U284 : MUX2_X1 port map( A => a_mod_24_port, B => a_adj_24_port, S => n166, 
                           Z => n337);
   U285 : MUX2_X1 port map( A => a_mod_23_port, B => a_adj_23_port, S => n166, 
                           Z => n338);
   U286 : MUX2_X1 port map( A => a_mod_22_port, B => a_adj_22_port, S => n166, 
                           Z => n339);
   U287 : MUX2_X1 port map( A => a_mod_21_port, B => a_adj_21_port, S => n166, 
                           Z => n340);
   U288 : MUX2_X1 port map( A => a_mod_20_port, B => a_adj_20_port, S => n166, 
                           Z => n341);
   U289 : MUX2_X1 port map( A => a_mod_19_port, B => a_adj_19_port, S => n166, 
                           Z => n342);
   U290 : MUX2_X1 port map( A => a_mod_18_port, B => a_adj_18_port, S => n166, 
                           Z => n343);
   U291 : MUX2_X1 port map( A => a_mod_17_port, B => a_adj_17_port, S => n166, 
                           Z => n344);
   U292 : MUX2_X1 port map( A => a_mod_16_port, B => a_adj_16_port, S => n167, 
                           Z => n345);
   U293 : MUX2_X1 port map( A => a_mod_15_port, B => a_adj_15_port, S => n167, 
                           Z => n346);
   U294 : MUX2_X1 port map( A => a_mod_14_port, B => a_adj_14_port, S => n167, 
                           Z => n347);
   U295 : MUX2_X1 port map( A => a_mod_13_port, B => a_adj_13_port, S => n167, 
                           Z => n348);
   U296 : MUX2_X1 port map( A => a_mod_12_port, B => a_adj_12_port, S => n167, 
                           Z => n349);
   U297 : MUX2_X1 port map( A => a_mod_11_port, B => a_adj_11_port, S => n167, 
                           Z => n350);
   U298 : MUX2_X1 port map( A => a_mod_10_port, B => a_adj_10_port, S => n167, 
                           Z => n351);
   U299 : MUX2_X1 port map( A => a_mod_9_port, B => a_adj_9_port, S => n167, Z 
                           => n352);
   U300 : MUX2_X1 port map( A => a_mod_8_port, B => a_adj_8_port, S => n167, Z 
                           => n353);
   U301 : MUX2_X1 port map( A => a_mod_7_port, B => a_adj_7_port, S => n167, Z 
                           => n354);
   U302 : MUX2_X1 port map( A => a_mod_6_port, B => a_adj_6_port, S => n167, Z 
                           => n355);
   U303 : MUX2_X1 port map( A => a_mod_5_port, B => a_adj_5_port, S => n167, Z 
                           => n356);
   U304 : MUX2_X1 port map( A => a_mod_4_port, B => a_adj_4_port, S => n166, Z 
                           => n357);
   U305 : MUX2_X1 port map( A => a_mod_3_port, B => a_adj_3_port, S => n165, Z 
                           => n358);
   U306 : MUX2_X1 port map( A => a_mod_2_port, B => a_adj_2_port, S => n165, Z 
                           => n359);
   U307 : MUX2_X1 port map( A => a_mod_1_port, B => a_adj_1_port, S => n167, Z 
                           => n360);
   U308 : MUX2_X1 port map( A => a_mod_0_port, B => a_adj_0_port, S => n167, Z 
                           => n361);
   U309 : INV_X1 port map( A => N17, ZN => n256);
   U310 : INV_X1 port map( A => lock, ZN => n222);
   U311 : NAND2_X1 port map( A1 => n362, A2 => n222, ZN => n255);
   U312 : NAND3_X1 port map( A1 => en, A2 => n72, A3 => n151, ZN => n254);

end SYN_div_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mul_DATA_SIZE16_STAGE10 is

   port( rst, clk, en, lock, sign : in std_logic;  a, b : in std_logic_vector 
         (15 downto 0);  o : out std_logic_vector (31 downto 0));

end Mul_DATA_SIZE16_STAGE10;

architecture SYN_mul_arch_struct of Mul_DATA_SIZE16_STAGE10 is

   component BoothMul_DATA_SIZE16_STAGE10
      port( rst, clk, en, lock, sign : in std_logic;  a, b : in 
            std_logic_vector (15 downto 0);  o : out std_logic_vector (31 
            downto 0));
   end component;

begin
   
   BM0 : BoothMul_DATA_SIZE16_STAGE10 port map( rst => rst, clk => clk, en => 
                           en, lock => lock, sign => sign, a(15) => a(15), 
                           a(14) => a(14), a(13) => a(13), a(12) => a(12), 
                           a(11) => a(11), a(10) => a(10), a(9) => a(9), a(8) 
                           => a(8), a(7) => a(7), a(6) => a(6), a(5) => a(5), 
                           a(4) => a(4), a(3) => a(3), a(2) => a(2), a(1) => 
                           a(1), a(0) => a(0), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           o(31) => o(31), o(30) => o(30), o(29) => o(29), 
                           o(28) => o(28), o(27) => o(27), o(26) => o(26), 
                           o(25) => o(25), o(24) => o(24), o(23) => o(23), 
                           o(22) => o(22), o(21) => o(21), o(20) => o(20), 
                           o(19) => o(19), o(18) => o(18), o(17) => o(17), 
                           o(16) => o(16), o(15) => o(15), o(14) => o(14), 
                           o(13) => o(13), o(12) => o(12), o(11) => o(11), 
                           o(10) => o(10), o(9) => o(9), o(8) => o(8), o(7) => 
                           o(7), o(6) => o(6), o(5) => o(5), o(4) => o(4), o(3)
                           => o(3), o(2) => o(2), o(1) => o(1), o(0) => o(0));

end SYN_mul_arch_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Alu_DATA_SIZE32 is

   port( f : in std_logic_vector (4 downto 0);  a, b : in std_logic_vector (31 
         downto 0);  o : out std_logic_vector (31 downto 0));

end Alu_DATA_SIZE32;

architecture SYN_alu_arch of Alu_DATA_SIZE32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component Shifter_DATA_SIZE32
      port( l_r, l_a, s_r : in std_logic;  a, b : in std_logic_vector (31 
            downto 0);  o : out std_logic_vector (31 downto 0));
   end component;
   
   component Adder_DATA_SIZE32_6
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal X_Logic0_port, b_new_31_port, b_new_30_port, b_new_29_port, 
      b_new_28_port, b_new_27_port, b_new_26_port, b_new_25_port, b_new_24_port
      , b_new_23_port, b_new_22_port, b_new_21_port, b_new_20_port, 
      b_new_19_port, b_new_18_port, b_new_17_port, b_new_16_port, b_new_15_port
      , b_new_14_port, b_new_13_port, b_new_12_port, b_new_11_port, 
      b_new_10_port, b_new_9_port, b_new_8_port, b_new_7_port, b_new_6_port, 
      b_new_5_port, b_new_4_port, b_new_3_port, b_new_2_port, b_new_1_port, 
      b_new_0_port, ado_31_port, ado_30_port, ado_29_port, ado_28_port, 
      ado_27_port, ado_26_port, ado_25_port, ado_24_port, ado_23_port, 
      ado_22_port, ado_21_port, ado_20_port, ado_19_port, ado_18_port, 
      ado_17_port, ado_16_port, ado_15_port, ado_14_port, ado_13_port, 
      ado_12_port, ado_11_port, ado_10_port, ado_9_port, ado_8_port, ado_7_port
      , ado_6_port, ado_5_port, ado_4_port, ado_3_port, ado_2_port, ado_1_port,
      ado_0_port, c_f, sho_31_port, sho_30_port, sho_29_port, sho_28_port, 
      sho_27_port, sho_26_port, sho_25_port, sho_24_port, sho_23_port, 
      sho_22_port, sho_21_port, sho_20_port, sho_19_port, sho_18_port, 
      sho_17_port, sho_16_port, sho_15_port, sho_14_port, sho_13_port, 
      sho_12_port, sho_11_port, sho_10_port, sho_9_port, sho_8_port, sho_7_port
      , sho_6_port, sho_5_port, sho_4_port, sho_3_port, sho_2_port, sho_1_port,
      sho_0_port, n72, n74, n75, n76, n77, n79, n80, n81, n82, n84, n85, n86, 
      n87, n89, n90, n91, n92, n94, n95, n96, n97, n99, n100, n101, n102, n104,
      n105, n107, n109, n110, n112, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n124, n125, n127, n128, n129, n130, n131, n132, n134, n135, 
      n136, n137, n139, n140, n141, n142, n144, n145, n146, n147, n149, n150, 
      n151, n152, n154, n155, n156, n157, n159, n160, n161, n162, n164, n165, 
      n166, n167, n169, n170, n171, n172, n174, n175, n176, n177, n179, n180, 
      n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, 
      n194, n195, n196, n197, n199, n200, n201, n202, n204, n205, n206, n207, 
      n209, n210, n211, n212, n214, n215, n216, n217, n219, n220, n221, n222, 
      n224, n225, n226, n227, n229, n230, n231, n232, n234, n235, n236, n238, 
      n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, 
      n251, n252, n253, n254, n255, n260, n261, n262, n263, n264, n265, n266, 
      n233, n237, n256, n257, n258, n259, n267, n268, n269, n270, n271, n272, 
      n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, 
      n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, 
      n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, 
      n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, 
      n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, 
      n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, 
      n345, n346 : std_logic;

begin
   
   X_Logic0_port <= '0';
   U229 : NAND3_X1 port map( A1 => n286, A2 => n320, A3 => b(9), ZN => n74);
   U230 : NAND3_X1 port map( A1 => n288, A2 => n318, A3 => b(8), ZN => n84);
   U231 : NAND3_X1 port map( A1 => n287, A2 => n316, A3 => b(7), ZN => n89);
   U232 : NAND3_X1 port map( A1 => n286, A2 => n314, A3 => b(6), ZN => n94);
   U233 : NAND3_X1 port map( A1 => n286, A2 => n312, A3 => b(5), ZN => n99);
   U234 : NAND3_X1 port map( A1 => n288, A2 => n310, A3 => b(4), ZN => n104);
   U235 : NAND3_X1 port map( A1 => n288, A2 => n308, A3 => b(3), ZN => n109);
   U236 : NAND3_X1 port map( A1 => n288, A2 => n345, A3 => b(31), ZN => n114);
   U237 : NAND3_X1 port map( A1 => n288, A2 => n118, A3 => b(30), ZN => n119);
   U238 : NAND3_X1 port map( A1 => n288, A2 => n306, A3 => n298, ZN => n124);
   U239 : NAND3_X1 port map( A1 => n288, A2 => n128, A3 => b(29), ZN => n129);
   U240 : NAND3_X1 port map( A1 => n288, A2 => n275, A3 => b(28), ZN => n134);
   U241 : NAND3_X1 port map( A1 => n288, A2 => n344, A3 => b(27), ZN => n139);
   U242 : NAND3_X1 port map( A1 => n288, A2 => n343, A3 => b(26), ZN => n144);
   U243 : NAND3_X1 port map( A1 => n288, A2 => n342, A3 => b(25), ZN => n149);
   U244 : NAND3_X1 port map( A1 => n288, A2 => n341, A3 => b(24), ZN => n154);
   U245 : NAND3_X1 port map( A1 => n288, A2 => n339, A3 => b(23), ZN => n159);
   U246 : NAND3_X1 port map( A1 => n288, A2 => n337, A3 => b(22), ZN => n164);
   U247 : NAND3_X1 port map( A1 => n288, A2 => n336, A3 => b(21), ZN => n169);
   U248 : NAND3_X1 port map( A1 => n288, A2 => n334, A3 => b(20), ZN => n174);
   U249 : NAND3_X1 port map( A1 => n288, A2 => n304, A3 => n296, ZN => n179);
   U250 : NAND3_X1 port map( A1 => n288, A2 => n183, A3 => b(19), ZN => n184);
   U251 : NAND3_X1 port map( A1 => n288, A2 => n188, A3 => b(18), ZN => n189);
   U252 : NAND3_X1 port map( A1 => n288, A2 => n193, A3 => b(17), ZN => n194);
   U253 : NAND3_X1 port map( A1 => n288, A2 => n333, A3 => b(16), ZN => n199);
   U254 : NAND3_X1 port map( A1 => n287, A2 => n332, A3 => b(15), ZN => n204);
   U255 : NAND3_X1 port map( A1 => n287, A2 => n330, A3 => b(14), ZN => n209);
   U256 : NAND3_X1 port map( A1 => n287, A2 => n328, A3 => b(13), ZN => n214);
   U257 : NAND3_X1 port map( A1 => n287, A2 => n326, A3 => b(12), ZN => n219);
   U258 : NAND3_X1 port map( A1 => n287, A2 => n324, A3 => b(11), ZN => n224);
   U259 : NAND3_X1 port map( A1 => n287, A2 => n322, A3 => b(10), ZN => n229);
   U260 : OAI33_X1 port map( A1 => n257, A2 => n269, A3 => n248, B1 => n238, B2
                           => f(0), B3 => n252, ZN => n249);
   U262 : XOR2_X1 port map( A => b(31), B => n273, Z => b_new_31_port);
   ADD0 : Adder_DATA_SIZE32_6 port map( cin => n346, a(31) => a(31), a(30) => 
                           a(30), a(29) => a(29), a(28) => n274, a(27) => a(27)
                           , a(26) => a(26), a(25) => a(25), a(24) => n340, 
                           a(23) => n338, a(22) => a(22), a(21) => n335, a(20) 
                           => a(20), a(19) => a(19), a(18) => a(18), a(17) => 
                           a(17), a(16) => a(16), a(15) => n331, a(14) => n329,
                           a(13) => n327, a(12) => n325, a(11) => n323, a(10) 
                           => n321, a(9) => n319, a(8) => n317, a(7) => n315, 
                           a(6) => n313, a(5) => n311, a(4) => n309, a(3) => 
                           n307, a(2) => n305, a(1) => a(1), a(0) => n302, 
                           b(31) => b_new_31_port, b(30) => b_new_30_port, 
                           b(29) => b_new_29_port, b(28) => b_new_28_port, 
                           b(27) => b_new_27_port, b(26) => b_new_26_port, 
                           b(25) => b_new_25_port, b(24) => b_new_24_port, 
                           b(23) => b_new_23_port, b(22) => b_new_22_port, 
                           b(21) => b_new_21_port, b(20) => b_new_20_port, 
                           b(19) => b_new_19_port, b(18) => b_new_18_port, 
                           b(17) => b_new_17_port, b(16) => b_new_16_port, 
                           b(15) => b_new_15_port, b(14) => b_new_14_port, 
                           b(13) => b_new_13_port, b(12) => b_new_12_port, 
                           b(11) => b_new_11_port, b(10) => b_new_10_port, b(9)
                           => b_new_9_port, b(8) => b_new_8_port, b(7) => 
                           b_new_7_port, b(6) => b_new_6_port, b(5) => 
                           b_new_5_port, b(4) => b_new_4_port, b(3) => 
                           b_new_3_port, b(2) => b_new_2_port, b(1) => 
                           b_new_1_port, b(0) => b_new_0_port, s(31) => 
                           ado_31_port, s(30) => ado_30_port, s(29) => 
                           ado_29_port, s(28) => ado_28_port, s(27) => 
                           ado_27_port, s(26) => ado_26_port, s(25) => 
                           ado_25_port, s(24) => ado_24_port, s(23) => 
                           ado_23_port, s(22) => ado_22_port, s(21) => 
                           ado_21_port, s(20) => ado_20_port, s(19) => 
                           ado_19_port, s(18) => ado_18_port, s(17) => 
                           ado_17_port, s(16) => ado_16_port, s(15) => 
                           ado_15_port, s(14) => ado_14_port, s(13) => 
                           ado_13_port, s(12) => ado_12_port, s(11) => 
                           ado_11_port, s(10) => ado_10_port, s(9) => 
                           ado_9_port, s(8) => ado_8_port, s(7) => ado_7_port, 
                           s(6) => ado_6_port, s(5) => ado_5_port, s(4) => 
                           ado_4_port, s(3) => ado_3_port, s(2) => ado_2_port, 
                           s(1) => ado_1_port, s(0) => ado_0_port, cout => c_f)
                           ;
   SHF0 : Shifter_DATA_SIZE32 port map( l_r => f(0), l_a => f(1), s_r => 
                           X_Logic0_port, a(31) => a(31), a(30) => a(30), a(29)
                           => a(29), a(28) => n274, a(27) => a(27), a(26) => 
                           a(26), a(25) => a(25), a(24) => n340, a(23) => n338,
                           a(22) => a(22), a(21) => n335, a(20) => a(20), a(19)
                           => a(19), a(18) => a(18), a(17) => a(17), a(16) => 
                           a(16), a(15) => n331, a(14) => n329, a(13) => n327, 
                           a(12) => n325, a(11) => n323, a(10) => n321, a(9) =>
                           n319, a(8) => n317, a(7) => n315, a(6) => n313, a(5)
                           => n311, a(4) => n309, a(3) => n307, a(2) => n305, 
                           a(1) => a(1), a(0) => n302, b(31) => b(31), b(30) =>
                           b(30), b(29) => b(29), b(28) => b(28), b(27) => 
                           b(27), b(26) => b(26), b(25) => b(25), b(24) => 
                           b(24), b(23) => b(23), b(22) => b(22), b(21) => 
                           b(21), b(20) => b(20), b(19) => b(19), b(18) => 
                           b(18), b(17) => b(17), b(16) => b(16), b(15) => 
                           b(15), b(14) => b(14), b(13) => b(13), b(12) => 
                           b(12), b(11) => b(11), b(10) => b(10), b(9) => b(9),
                           b(8) => b(8), b(7) => b(7), b(6) => b(6), b(5) => 
                           b(5), b(4) => b(4), b(3) => b(3), b(2) => n298, b(1)
                           => n296, b(0) => n270, o(31) => sho_31_port, o(30) 
                           => sho_30_port, o(29) => sho_29_port, o(28) => 
                           sho_28_port, o(27) => sho_27_port, o(26) => 
                           sho_26_port, o(25) => sho_25_port, o(24) => 
                           sho_24_port, o(23) => sho_23_port, o(22) => 
                           sho_22_port, o(21) => sho_21_port, o(20) => 
                           sho_20_port, o(19) => sho_19_port, o(18) => 
                           sho_18_port, o(17) => sho_17_port, o(16) => 
                           sho_16_port, o(15) => sho_15_port, o(14) => 
                           sho_14_port, o(13) => sho_13_port, o(12) => 
                           sho_12_port, o(11) => sho_11_port, o(10) => 
                           sho_10_port, o(9) => sho_9_port, o(8) => sho_8_port,
                           o(7) => sho_7_port, o(6) => sho_6_port, o(5) => 
                           sho_5_port, o(4) => sho_4_port, o(3) => sho_3_port, 
                           o(2) => sho_2_port, o(1) => sho_1_port, o(0) => 
                           sho_0_port);
   U2 : NOR4_X1 port map( A1 => ado_28_port, A2 => ado_29_port, A3 => 
                           ado_2_port, A4 => ado_30_port, ZN => n278);
   U3 : INV_X1 port map( A => n269, ZN => n256);
   U4 : INV_X1 port map( A => n328, ZN => n327);
   U5 : INV_X1 port map( A => n330, ZN => n329);
   U6 : CLKBUF_X1 port map( A => f(4), Z => n346);
   U7 : CLKBUF_X1 port map( A => n266, Z => n267);
   U8 : AND2_X1 port map( A1 => n277, A2 => n268, ZN => n233);
   U9 : AND2_X1 port map( A1 => n278, A2 => n233, ZN => n255);
   U10 : INV_X1 port map( A => n267, ZN => n237);
   U11 : XNOR2_X1 port map( A => n251, B => n256, ZN => n250);
   U12 : AOI22_X1 port map( A1 => c_f, A2 => f(2), B1 => n253, B2 => n238, ZN 
                           => n257);
   U13 : CLKBUF_X1 port map( A => f(4), Z => n258);
   U14 : CLKBUF_X1 port map( A => n346, Z => n259);
   U15 : AND2_X1 port map( A1 => n279, A2 => n271, ZN => n268);
   U16 : INV_X1 port map( A => f(0), ZN => n269);
   U17 : XNOR2_X1 port map( A => n267, B => n264, ZN => n253);
   U18 : CLKBUF_X1 port map( A => b(0), Z => n270);
   U19 : XOR2_X1 port map( A => b(0), B => f(4), Z => b_new_0_port);
   U20 : XNOR2_X1 port map( A => n346, B => n231, ZN => b_new_10_port);
   U21 : XNOR2_X1 port map( A => n259, B => n201, ZN => b_new_16_port);
   U22 : XNOR2_X1 port map( A => n346, B => n196, ZN => b_new_17_port);
   U23 : XNOR2_X1 port map( A => n259, B => n206, ZN => b_new_15_port);
   U24 : AOI22_X1 port map( A1 => sho_29_port, A2 => n293, B1 => ado_29_port, 
                           B2 => n290, ZN => n130);
   U25 : AOI22_X1 port map( A1 => sho_27_port, A2 => n293, B1 => ado_27_port, 
                           B2 => n290, ZN => n140);
   U26 : AOI22_X1 port map( A1 => sho_26_port, A2 => n293, B1 => ado_26_port, 
                           B2 => n290, ZN => n145);
   U27 : AOI22_X1 port map( A1 => sho_25_port, A2 => n293, B1 => ado_25_port, 
                           B2 => n290, ZN => n150);
   U28 : AOI22_X1 port map( A1 => sho_21_port, A2 => n293, B1 => ado_21_port, 
                           B2 => n290, ZN => n170);
   U29 : AOI22_X1 port map( A1 => sho_22_port, A2 => n293, B1 => ado_22_port, 
                           B2 => n290, ZN => n165);
   U30 : AOI22_X1 port map( A1 => sho_23_port, A2 => n293, B1 => ado_23_port, 
                           B2 => n290, ZN => n160);
   U31 : AOI22_X1 port map( A1 => sho_13_port, A2 => n292, B1 => ado_13_port, 
                           B2 => n289, ZN => n215);
   U32 : AOI22_X1 port map( A1 => sho_14_port, A2 => n292, B1 => ado_14_port, 
                           B2 => n289, ZN => n210);
   U33 : AOI22_X1 port map( A1 => sho_15_port, A2 => n292, B1 => ado_15_port, 
                           B2 => n289, ZN => n205);
   U34 : AOI22_X1 port map( A1 => sho_17_port, A2 => n292, B1 => ado_17_port, 
                           B2 => n289, ZN => n195);
   U35 : AOI22_X1 port map( A1 => sho_18_port, A2 => n292, B1 => ado_18_port, 
                           B2 => n289, ZN => n190);
   U36 : AOI22_X1 port map( A1 => sho_19_port, A2 => n292, B1 => ado_19_port, 
                           B2 => n289, ZN => n185);
   U37 : OR4_X1 port map( A1 => ado_17_port, A2 => ado_18_port, A3 => 
                           ado_19_port, A4 => ado_1_port, ZN => n261);
   U38 : INV_X1 port map( A => n299, ZN => n298);
   U39 : BUF_X1 port map( A => n80, Z => n283);
   U40 : BUF_X1 port map( A => n80, Z => n284);
   U41 : BUF_X1 port map( A => n80, Z => n285);
   U42 : NOR4_X1 port map( A1 => ado_24_port, A2 => ado_25_port, A3 => 
                           ado_26_port, A4 => ado_27_port, ZN => n279);
   U43 : AOI22_X1 port map( A1 => sho_31_port, A2 => n294, B1 => n237, B2 => 
                           n291, ZN => n115);
   U44 : AOI22_X1 port map( A1 => sho_28_port, A2 => n293, B1 => ado_28_port, 
                           B2 => n290, ZN => n135);
   U45 : AOI22_X1 port map( A1 => sho_30_port, A2 => n293, B1 => ado_30_port, 
                           B2 => n290, ZN => n120);
   U46 : AOI22_X1 port map( A1 => sho_24_port, A2 => n293, B1 => ado_24_port, 
                           B2 => n290, ZN => n155);
   U47 : AOI22_X1 port map( A1 => sho_20_port, A2 => n293, B1 => ado_20_port, 
                           B2 => n290, ZN => n175);
   U48 : AOI22_X1 port map( A1 => sho_12_port, A2 => n292, B1 => ado_12_port, 
                           B2 => n289, ZN => n220);
   U49 : AOI22_X1 port map( A1 => sho_16_port, A2 => n292, B1 => ado_16_port, 
                           B2 => n289, ZN => n200);
   U50 : AOI221_X1 port map( B1 => n286, B2 => n295, C1 => n270, C2 => n283, A 
                           => n280, ZN => n232);
   U51 : AOI22_X1 port map( A1 => sho_0_port, A2 => n292, B1 => ado_0_port, B2 
                           => n289, ZN => n235);
   U52 : OAI211_X1 port map( C1 => n177, C2 => n304, A => n179, B => n180, ZN 
                           => o(1));
   U53 : AOI221_X1 port map( B1 => n286, B2 => n297, C1 => n296, C2 => n283, A 
                           => n280, ZN => n177);
   U54 : AOI22_X1 port map( A1 => sho_1_port, A2 => n292, B1 => ado_1_port, B2 
                           => n289, ZN => n180);
   U55 : OAI211_X1 port map( C1 => n122, C2 => n306, A => n124, B => n125, ZN 
                           => o(2));
   U56 : AOI221_X1 port map( B1 => n286, B2 => n299, C1 => n298, C2 => n284, A 
                           => n281, ZN => n122);
   U57 : AOI22_X1 port map( A1 => sho_2_port, A2 => n293, B1 => ado_2_port, B2 
                           => n290, ZN => n125);
   U58 : OAI211_X1 port map( C1 => n227, C2 => n322, A => n229, B => n230, ZN 
                           => o(10));
   U59 : AOI221_X1 port map( B1 => n286, B2 => n231, C1 => b(10), C2 => n283, A
                           => n280, ZN => n227);
   U60 : AOI22_X1 port map( A1 => sho_10_port, A2 => n292, B1 => ado_10_port, 
                           B2 => n289, ZN => n230);
   U61 : OAI211_X1 port map( C1 => n222, C2 => n324, A => n224, B => n225, ZN 
                           => o(11));
   U62 : AOI221_X1 port map( B1 => n286, B2 => n226, C1 => b(11), C2 => n283, A
                           => n280, ZN => n222);
   U63 : AOI22_X1 port map( A1 => sho_11_port, A2 => n292, B1 => ado_11_port, 
                           B2 => n289, ZN => n225);
   U64 : OAI211_X1 port map( C1 => n107, C2 => n308, A => n109, B => n110, ZN 
                           => o(3));
   U65 : AOI221_X1 port map( B1 => n287, B2 => n300, C1 => b(3), C2 => n285, A 
                           => n282, ZN => n107);
   U66 : AOI22_X1 port map( A1 => sho_3_port, A2 => n294, B1 => ado_3_port, B2 
                           => n291, ZN => n110);
   U67 : OAI211_X1 port map( C1 => n102, C2 => n310, A => n104, B => n105, ZN 
                           => o(4));
   U68 : AOI221_X1 port map( B1 => n287, B2 => n301, C1 => b(4), C2 => n285, A 
                           => n282, ZN => n102);
   U69 : AOI22_X1 port map( A1 => sho_4_port, A2 => n294, B1 => ado_4_port, B2 
                           => n291, ZN => n105);
   U70 : OAI211_X1 port map( C1 => n97, C2 => n312, A => n99, B => n100, ZN => 
                           o(5));
   U71 : AOI221_X1 port map( B1 => n287, B2 => n101, C1 => b(5), C2 => n285, A 
                           => n282, ZN => n97);
   U72 : AOI22_X1 port map( A1 => sho_5_port, A2 => n294, B1 => ado_5_port, B2 
                           => n291, ZN => n100);
   U73 : OAI211_X1 port map( C1 => n92, C2 => n314, A => n94, B => n95, ZN => 
                           o(6));
   U74 : AOI221_X1 port map( B1 => n287, B2 => n96, C1 => b(6), C2 => n285, A 
                           => n282, ZN => n92);
   U75 : AOI22_X1 port map( A1 => sho_6_port, A2 => n294, B1 => ado_6_port, B2 
                           => n291, ZN => n95);
   U76 : OAI211_X1 port map( C1 => n87, C2 => n316, A => n89, B => n90, ZN => 
                           o(7));
   U77 : AOI221_X1 port map( B1 => n287, B2 => n91, C1 => b(7), C2 => n285, A 
                           => n282, ZN => n87);
   U78 : AOI22_X1 port map( A1 => sho_7_port, A2 => n294, B1 => ado_7_port, B2 
                           => n291, ZN => n90);
   U79 : OAI211_X1 port map( C1 => n82, C2 => n318, A => n84, B => n85, ZN => 
                           o(8));
   U80 : AOI221_X1 port map( B1 => n287, B2 => n86, C1 => b(8), C2 => n285, A 
                           => n282, ZN => n82);
   U81 : AOI22_X1 port map( A1 => sho_8_port, A2 => n294, B1 => ado_8_port, B2 
                           => n291, ZN => n85);
   U82 : OAI211_X1 port map( C1 => n72, C2 => n320, A => n74, B => n75, ZN => 
                           o(9));
   U83 : AOI221_X1 port map( B1 => n287, B2 => n79, C1 => n285, C2 => b(9), A 
                           => n282, ZN => n72);
   U84 : AOI22_X1 port map( A1 => sho_9_port, A2 => n294, B1 => ado_9_port, B2 
                           => n291, ZN => n75);
   U85 : NOR4_X1 port map( A1 => n260, A2 => n261, A3 => n262, A4 => n263, ZN 
                           => n254);
   U86 : OR4_X1 port map( A1 => ado_0_port, A2 => ado_10_port, A3 => 
                           ado_11_port, A4 => ado_12_port, ZN => n263);
   U87 : OR4_X1 port map( A1 => ado_13_port, A2 => ado_14_port, A3 => 
                           ado_15_port, A4 => ado_16_port, ZN => n262);
   U88 : OR4_X1 port map( A1 => ado_20_port, A2 => ado_21_port, A3 => 
                           ado_22_port, A4 => ado_23_port, ZN => n260);
   U89 : INV_X1 port map( A => b(2), ZN => n299);
   U90 : INV_X1 port map( A => b(1), ZN => n297);
   U91 : INV_X1 port map( A => b(10), ZN => n231);
   U92 : INV_X1 port map( A => b(15), ZN => n206);
   U93 : INV_X1 port map( A => b(13), ZN => n216);
   U94 : INV_X1 port map( A => b(7), ZN => n91);
   U95 : INV_X1 port map( A => b(11), ZN => n226);
   U96 : INV_X1 port map( A => b(9), ZN => n79);
   U97 : INV_X1 port map( A => b(17), ZN => n196);
   U98 : INV_X1 port map( A => b(16), ZN => n201);
   U99 : INV_X1 port map( A => b(12), ZN => n221);
   U100 : INV_X1 port map( A => b(6), ZN => n96);
   U101 : INV_X1 port map( A => b(8), ZN => n86);
   U102 : INV_X1 port map( A => b(5), ZN => n101);
   U103 : INV_X1 port map( A => b(14), ZN => n211);
   U104 : INV_X1 port map( A => b(18), ZN => n191);
   U105 : INV_X1 port map( A => b(19), ZN => n186);
   U106 : INV_X1 port map( A => b(23), ZN => n161);
   U107 : INV_X1 port map( A => b(25), ZN => n151);
   U108 : INV_X1 port map( A => b(24), ZN => n156);
   U109 : INV_X1 port map( A => b(22), ZN => n166);
   U110 : INV_X1 port map( A => b(21), ZN => n171);
   U111 : INV_X1 port map( A => b(20), ZN => n176);
   U112 : INV_X1 port map( A => b(28), ZN => n136);
   U113 : INV_X1 port map( A => b(29), ZN => n131);
   U114 : NOR4_X1 port map( A1 => ado_6_port, A2 => ado_7_port, A3 => 
                           ado_8_port, A4 => ado_9_port, ZN => n271);
   U115 : INV_X1 port map( A => b_new_31_port, ZN => n265);
   U116 : INV_X1 port map( A => n272, ZN => n288);
   U117 : INV_X1 port map( A => n272, ZN => n287);
   U118 : NOR3_X1 port map( A1 => n236, A2 => n259, A3 => n269, ZN => n80);
   U119 : AOI221_X1 port map( B1 => n287, B2 => n116, C1 => b(31), C2 => n285, 
                           A => n282, ZN => n112);
   U120 : INV_X1 port map( A => b(31), ZN => n116);
   U121 : AOI221_X1 port map( B1 => n286, B2 => n221, C1 => b(12), C2 => n283, 
                           A => n280, ZN => n217);
   U122 : AOI221_X1 port map( B1 => n286, B2 => n216, C1 => b(13), C2 => n283, 
                           A => n280, ZN => n212);
   U123 : AOI221_X1 port map( B1 => n286, B2 => n211, C1 => b(14), C2 => n283, 
                           A => n280, ZN => n207);
   U124 : AOI221_X1 port map( B1 => n286, B2 => n206, C1 => b(15), C2 => n283, 
                           A => n280, ZN => n202);
   U125 : AOI221_X1 port map( B1 => n286, B2 => n201, C1 => b(16), C2 => n283, 
                           A => n280, ZN => n197);
   U126 : AOI221_X1 port map( B1 => n286, B2 => n196, C1 => b(17), C2 => n283, 
                           A => n280, ZN => n192);
   U127 : AOI221_X1 port map( B1 => n286, B2 => n191, C1 => b(18), C2 => n283, 
                           A => n280, ZN => n187);
   U128 : AOI221_X1 port map( B1 => n286, B2 => n186, C1 => b(19), C2 => n283, 
                           A => n280, ZN => n182);
   U129 : AOI221_X1 port map( B1 => n286, B2 => n176, C1 => b(20), C2 => n284, 
                           A => n281, ZN => n172);
   U130 : AOI221_X1 port map( B1 => n287, B2 => n171, C1 => b(21), C2 => n284, 
                           A => n281, ZN => n167);
   U131 : AOI221_X1 port map( B1 => n286, B2 => n166, C1 => b(22), C2 => n284, 
                           A => n281, ZN => n162);
   U132 : AOI221_X1 port map( B1 => n287, B2 => n161, C1 => b(23), C2 => n284, 
                           A => n281, ZN => n157);
   U133 : AOI221_X1 port map( B1 => n287, B2 => n156, C1 => b(24), C2 => n284, 
                           A => n281, ZN => n152);
   U134 : AOI221_X1 port map( B1 => n287, B2 => n151, C1 => b(25), C2 => n284, 
                           A => n281, ZN => n147);
   U135 : AOI221_X1 port map( B1 => n287, B2 => n146, C1 => b(26), C2 => n284, 
                           A => n281, ZN => n142);
   U136 : AOI221_X1 port map( B1 => n286, B2 => n141, C1 => b(27), C2 => n284, 
                           A => n281, ZN => n137);
   U137 : AOI221_X1 port map( B1 => n286, B2 => n136, C1 => b(28), C2 => n284, 
                           A => n281, ZN => n132);
   U138 : AOI221_X1 port map( B1 => n287, B2 => n131, C1 => b(29), C2 => n284, 
                           A => n281, ZN => n127);
   U139 : AOI221_X1 port map( B1 => n288, B2 => n121, C1 => b(30), C2 => n284, 
                           A => n281, ZN => n117);
   U140 : BUF_X1 port map( A => n76, Z => n292);
   U141 : BUF_X1 port map( A => n76, Z => n293);
   U142 : BUF_X1 port map( A => n81, Z => n280);
   U143 : BUF_X1 port map( A => n81, Z => n281);
   U144 : BUF_X1 port map( A => n77, Z => n289);
   U145 : BUF_X1 port map( A => n77, Z => n290);
   U146 : BUF_X1 port map( A => n76, Z => n294);
   U147 : BUF_X1 port map( A => n81, Z => n282);
   U148 : BUF_X1 port map( A => n77, Z => n291);
   U149 : NOR2_X1 port map( A1 => n302, A2 => n272, ZN => n240);
   U150 : INV_X1 port map( A => b(30), ZN => n121);
   U151 : INV_X1 port map( A => b(26), ZN => n146);
   U152 : INV_X1 port map( A => b(27), ZN => n141);
   U153 : INV_X1 port map( A => n341, ZN => n340);
   U154 : INV_X1 port map( A => n332, ZN => n331);
   U155 : INV_X1 port map( A => n308, ZN => n307);
   U156 : INV_X1 port map( A => n339, ZN => n338);
   U157 : INV_X1 port map( A => n312, ZN => n311);
   U158 : INV_X1 port map( A => n326, ZN => n325);
   U159 : OAI211_X1 port map( C1 => n117, C2 => n118, A => n119, B => n120, ZN 
                           => o(30));
   U160 : OAI211_X1 port map( C1 => n112, C2 => n345, A => n114, B => n115, ZN 
                           => o(31));
   U161 : OAI211_X1 port map( C1 => n127, C2 => n128, A => n129, B => n130, ZN 
                           => o(29));
   U162 : OAI211_X1 port map( C1 => n157, C2 => n339, A => n159, B => n160, ZN 
                           => o(23));
   U163 : OAI211_X1 port map( C1 => n197, C2 => n333, A => n199, B => n200, ZN 
                           => o(16));
   U164 : OAI211_X1 port map( C1 => n192, C2 => n193, A => n194, B => n195, ZN 
                           => o(17));
   U165 : OAI211_X1 port map( C1 => n217, C2 => n326, A => n219, B => n220, ZN 
                           => o(12));
   U166 : OAI211_X1 port map( C1 => n212, C2 => n328, A => n214, B => n215, ZN 
                           => o(13));
   U167 : OAI211_X1 port map( C1 => n207, C2 => n330, A => n209, B => n210, ZN 
                           => o(14));
   U168 : OAI211_X1 port map( C1 => n202, C2 => n332, A => n204, B => n205, ZN 
                           => o(15));
   U169 : OAI211_X1 port map( C1 => n132, C2 => n275, A => n134, B => n135, ZN 
                           => o(28));
   U170 : OAI211_X1 port map( C1 => n137, C2 => n344, A => n139, B => n140, ZN 
                           => o(27));
   U171 : OAI211_X1 port map( C1 => n147, C2 => n342, A => n149, B => n150, ZN 
                           => o(25));
   U172 : OAI211_X1 port map( C1 => n142, C2 => n343, A => n144, B => n145, ZN 
                           => o(26));
   U173 : OAI211_X1 port map( C1 => n152, C2 => n341, A => n154, B => n155, ZN 
                           => o(24));
   U174 : OAI211_X1 port map( C1 => n187, C2 => n188, A => n189, B => n190, ZN 
                           => o(18));
   U175 : OAI211_X1 port map( C1 => n182, C2 => n183, A => n184, B => n185, ZN 
                           => o(19));
   U176 : OAI211_X1 port map( C1 => n172, C2 => n334, A => n174, B => n175, ZN 
                           => o(20));
   U177 : OAI211_X1 port map( C1 => n167, C2 => n336, A => n169, B => n170, ZN 
                           => o(21));
   U178 : OAI211_X1 port map( C1 => n162, C2 => n337, A => n164, B => n165, ZN 
                           => o(22));
   U179 : AOI211_X1 port map( C1 => n276, C2 => n247, A => f(0), B => n248, ZN 
                           => n244);
   U180 : NOR2_X1 port map( A1 => n272, A2 => f(0), ZN => n81);
   U181 : NOR2_X1 port map( A1 => n236, A2 => f(0), ZN => n77);
   U182 : OR4_X1 port map( A1 => n247, A2 => f(2), A3 => f(3), A4 => n259, ZN 
                           => n272);
   U183 : INV_X1 port map( A => f(2), ZN => n238);
   U184 : INV_X1 port map( A => a(19), ZN => n183);
   U185 : INV_X1 port map( A => a(17), ZN => n193);
   U186 : INV_X1 port map( A => a(18), ZN => n188);
   U187 : INV_X1 port map( A => a(29), ZN => n128);
   U188 : INV_X1 port map( A => a(30), ZN => n118);
   U189 : INV_X1 port map( A => a(15), ZN => n332);
   U190 : INV_X1 port map( A => a(13), ZN => n328);
   U191 : INV_X1 port map( A => a(3), ZN => n308);
   U192 : INV_X1 port map( A => a(5), ZN => n312);
   U193 : INV_X1 port map( A => a(31), ZN => n345);
   U194 : INV_X1 port map( A => a(23), ZN => n339);
   U195 : INV_X1 port map( A => a(16), ZN => n333);
   U196 : INV_X1 port map( A => a(20), ZN => n334);
   U197 : INV_X1 port map( A => a(22), ZN => n337);
   U198 : INV_X1 port map( A => a(24), ZN => n341);
   U199 : INV_X1 port map( A => a(25), ZN => n342);
   U200 : INV_X1 port map( A => a(26), ZN => n343);
   U201 : INV_X1 port map( A => a(21), ZN => n336);
   U202 : BUF_X4 port map( A => n258, Z => n273);
   U203 : INV_X1 port map( A => n275, ZN => n274);
   U204 : INV_X1 port map( A => a(28), ZN => n275);
   U205 : OAI222_X1 port map( A1 => n266, A2 => n265, B1 => b_new_31_port, B2 
                           => n345, C1 => a(31), C2 => ado_31_port, ZN => n264)
                           ;
   U206 : INV_X1 port map( A => ado_31_port, ZN => n266);
   U207 : XNOR2_X1 port map( A => n273, B => n186, ZN => b_new_19_port);
   U208 : XNOR2_X1 port map( A => n273, B => n191, ZN => b_new_18_port);
   U209 : XNOR2_X1 port map( A => n273, B => n226, ZN => b_new_11_port);
   U210 : CLKBUF_X1 port map( A => c_f, Z => n276);
   U211 : XNOR2_X1 port map( A => n259, B => n211, ZN => b_new_14_port);
   U212 : XNOR2_X1 port map( A => n273, B => n176, ZN => b_new_20_port);
   U213 : XNOR2_X1 port map( A => n259, B => n171, ZN => b_new_21_port);
   U214 : INV_X1 port map( A => n336, ZN => n335);
   U215 : XNOR2_X1 port map( A => n273, B => n221, ZN => b_new_12_port);
   U216 : XNOR2_X1 port map( A => n273, B => n216, ZN => b_new_13_port);
   U217 : XNOR2_X1 port map( A => n273, B => n297, ZN => b_new_1_port);
   U218 : XNOR2_X1 port map( A => n273, B => n300, ZN => b_new_3_port);
   U219 : XNOR2_X1 port map( A => n346, B => n299, ZN => b_new_2_port);
   U220 : NOR2_X1 port map( A1 => f(1), A2 => n246, ZN => n245);
   U221 : AOI211_X1 port map( C1 => n269, C2 => f(1), A => n238, B => n239, ZN 
                           => n76);
   U222 : INV_X1 port map( A => f(1), ZN => n247);
   U223 : NOR4_X1 port map( A1 => ado_3_port, A2 => ado_4_port, A3 => 
                           ado_31_port, A4 => ado_5_port, ZN => n277);
   U224 : OAI211_X1 port map( C1 => n244, C2 => n245, A => n238, B => f(3), ZN 
                           => n243);
   U225 : OR2_X1 port map( A1 => n273, A2 => f(3), ZN => n239);
   U226 : OR3_X1 port map( A1 => f(2), A2 => f(3), A3 => f(1), ZN => n236);
   U227 : INV_X1 port map( A => n270, ZN => n295);
   U228 : XNOR2_X1 port map( A => n346, B => n79, ZN => b_new_9_port);
   U261 : XNOR2_X1 port map( A => n346, B => n301, ZN => b_new_4_port);
   U263 : NAND2_X1 port map( A1 => n255, A2 => n254, ZN => n246);
   U264 : AND2_X1 port map( A1 => n246, A2 => n253, ZN => n252);
   U265 : INV_X1 port map( A => n246, ZN => n248);
   U266 : XNOR2_X1 port map( A => n273, B => n121, ZN => b_new_30_port);
   U267 : XNOR2_X1 port map( A => n273, B => n131, ZN => b_new_29_port);
   U268 : XNOR2_X1 port map( A => n259, B => n136, ZN => b_new_28_port);
   U269 : XNOR2_X1 port map( A => n273, B => n161, ZN => b_new_23_port);
   U270 : XNOR2_X1 port map( A => n273, B => n86, ZN => b_new_8_port);
   U271 : XNOR2_X1 port map( A => n273, B => n96, ZN => b_new_6_port);
   U272 : XNOR2_X1 port map( A => n259, B => n141, ZN => b_new_27_port);
   U273 : XNOR2_X1 port map( A => n259, B => n146, ZN => b_new_26_port);
   U274 : XNOR2_X1 port map( A => n259, B => n151, ZN => b_new_25_port);
   U275 : XNOR2_X1 port map( A => n259, B => n156, ZN => b_new_24_port);
   U276 : XNOR2_X1 port map( A => n346, B => n91, ZN => b_new_7_port);
   U277 : OAI21_X1 port map( B1 => n242, B2 => f(3), A => n243, ZN => n241);
   U278 : AOI22_X1 port map( A1 => n240, A2 => n270, B1 => n241, B2 => n273, ZN
                           => n234);
   U279 : XNOR2_X1 port map( A => n273, B => n101, ZN => b_new_5_port);
   U280 : XNOR2_X1 port map( A => n273, B => n166, ZN => b_new_22_port);
   U281 : AOI22_X1 port map( A1 => n249, A2 => n247, B1 => n250, B2 => f(1), ZN
                           => n242);
   U282 : AOI22_X1 port map( A1 => c_f, A2 => f(2), B1 => n238, B2 => n253, ZN 
                           => n251);
   U283 : OAI211_X1 port map( C1 => n232, C2 => n303, A => n235, B => n234, ZN 
                           => o(0));
   U284 : INV_X1 port map( A => n272, ZN => n286);
   U285 : INV_X2 port map( A => n297, ZN => n296);
   U286 : INV_X1 port map( A => b(3), ZN => n300);
   U287 : INV_X1 port map( A => b(4), ZN => n301);
   U288 : INV_X1 port map( A => n303, ZN => n302);
   U289 : INV_X1 port map( A => a(0), ZN => n303);
   U290 : INV_X1 port map( A => a(1), ZN => n304);
   U291 : INV_X1 port map( A => n306, ZN => n305);
   U292 : INV_X1 port map( A => a(2), ZN => n306);
   U293 : INV_X1 port map( A => n310, ZN => n309);
   U294 : INV_X1 port map( A => a(4), ZN => n310);
   U295 : INV_X1 port map( A => n314, ZN => n313);
   U296 : INV_X1 port map( A => a(6), ZN => n314);
   U297 : INV_X1 port map( A => n316, ZN => n315);
   U298 : INV_X1 port map( A => a(7), ZN => n316);
   U299 : INV_X1 port map( A => n318, ZN => n317);
   U300 : INV_X1 port map( A => a(8), ZN => n318);
   U301 : INV_X1 port map( A => n320, ZN => n319);
   U302 : INV_X1 port map( A => a(9), ZN => n320);
   U303 : INV_X1 port map( A => n322, ZN => n321);
   U304 : INV_X1 port map( A => a(10), ZN => n322);
   U305 : INV_X1 port map( A => n324, ZN => n323);
   U306 : INV_X1 port map( A => a(11), ZN => n324);
   U307 : INV_X1 port map( A => a(12), ZN => n326);
   U308 : INV_X1 port map( A => a(14), ZN => n330);
   U309 : INV_X1 port map( A => a(27), ZN => n344);

end SYN_alu_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE32_3 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0);  
         dout : out std_logic_vector (31 downto 0));

end Mux_DATA_SIZE32_3;

architecture SYN_mux_arch of Mux_DATA_SIZE32_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47,
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66 : std_logic;

begin
   
   U19 : INV_X2 port map( A => n44, ZN => dout(2));
   U1 : INV_X1 port map( A => sel, ZN => n35);
   U2 : INV_X1 port map( A => n55, ZN => dout(1));
   U3 : INV_X1 port map( A => n41, ZN => dout(3));
   U4 : INV_X1 port map( A => n40, ZN => dout(4));
   U5 : INV_X1 port map( A => n38, ZN => dout(6));
   U6 : INV_X1 port map( A => n37, ZN => dout(7));
   U7 : INV_X1 port map( A => n63, ZN => dout(12));
   U8 : INV_X1 port map( A => n62, ZN => dout(13));
   U9 : INV_X1 port map( A => n61, ZN => dout(14));
   U10 : INV_X1 port map( A => n66, ZN => dout(0));
   U11 : AOI22_X1 port map( A1 => din0(7), A2 => n35, B1 => din1(7), B2 => sel,
                           ZN => n37);
   U12 : INV_X1 port map( A => n64, ZN => dout(11));
   U13 : INV_X1 port map( A => n34, ZN => dout(9));
   U14 : AOI22_X1 port map( A1 => din0(9), A2 => n35, B1 => sel, B2 => din1(9),
                           ZN => n34);
   U15 : INV_X1 port map( A => n65, ZN => dout(10));
   U16 : AOI22_X1 port map( A1 => din0(3), A2 => n35, B1 => din1(3), B2 => sel,
                           ZN => n41);
   U17 : AOI22_X1 port map( A1 => din0(4), A2 => n35, B1 => din1(4), B2 => sel,
                           ZN => n40);
   U18 : AOI22_X1 port map( A1 => din0(6), A2 => n35, B1 => din1(6), B2 => sel,
                           ZN => n38);
   U20 : INV_X1 port map( A => n36, ZN => dout(8));
   U21 : AOI22_X1 port map( A1 => din0(8), A2 => n35, B1 => din1(8), B2 => sel,
                           ZN => n36);
   U22 : INV_X1 port map( A => n39, ZN => dout(5));
   U23 : AOI22_X1 port map( A1 => din0(5), A2 => n35, B1 => din1(5), B2 => sel,
                           ZN => n39);
   U24 : AOI22_X1 port map( A1 => din0(2), A2 => n35, B1 => din1(2), B2 => sel,
                           ZN => n44);
   U25 : AOI22_X1 port map( A1 => din0(1), A2 => n35, B1 => din1(1), B2 => sel,
                           ZN => n55);
   U26 : INV_X1 port map( A => n42, ZN => dout(31));
   U27 : AOI22_X1 port map( A1 => din0(31), A2 => n35, B1 => din1(31), B2 => 
                           sel, ZN => n42);
   U28 : INV_X1 port map( A => n58, ZN => dout(17));
   U29 : INV_X1 port map( A => n59, ZN => dout(16));
   U30 : INV_X1 port map( A => n60, ZN => dout(15));
   U31 : INV_X1 port map( A => n51, ZN => dout(23));
   U32 : AOI22_X1 port map( A1 => din0(23), A2 => n35, B1 => din1(23), B2 => 
                           sel, ZN => n51);
   U33 : INV_X1 port map( A => n50, ZN => dout(24));
   U34 : AOI22_X1 port map( A1 => din0(24), A2 => n35, B1 => din1(24), B2 => 
                           sel, ZN => n50);
   U35 : INV_X1 port map( A => n54, ZN => dout(20));
   U36 : AOI22_X1 port map( A1 => din0(20), A2 => n35, B1 => din1(20), B2 => 
                           sel, ZN => n54);
   U37 : INV_X1 port map( A => n49, ZN => dout(25));
   U38 : AOI22_X1 port map( A1 => din0(25), A2 => n35, B1 => din1(25), B2 => 
                           sel, ZN => n49);
   U39 : INV_X1 port map( A => n53, ZN => dout(21));
   U40 : AOI22_X1 port map( A1 => din0(21), A2 => n35, B1 => din1(21), B2 => 
                           sel, ZN => n53);
   U41 : INV_X1 port map( A => n45, ZN => dout(29));
   U42 : AOI22_X1 port map( A1 => din0(29), A2 => n35, B1 => din1(29), B2 => 
                           sel, ZN => n45);
   U43 : INV_X1 port map( A => n46, ZN => dout(28));
   U44 : AOI22_X1 port map( A1 => din0(28), A2 => n35, B1 => din1(28), B2 => 
                           sel, ZN => n46);
   U45 : INV_X1 port map( A => n52, ZN => dout(22));
   U46 : AOI22_X1 port map( A1 => din0(22), A2 => n35, B1 => din1(22), B2 => 
                           sel, ZN => n52);
   U47 : INV_X1 port map( A => n57, ZN => dout(18));
   U48 : INV_X1 port map( A => n56, ZN => dout(19));
   U49 : INV_X1 port map( A => n43, ZN => dout(30));
   U50 : AOI22_X1 port map( A1 => din0(30), A2 => n35, B1 => din1(30), B2 => 
                           sel, ZN => n43);
   U51 : INV_X1 port map( A => n48, ZN => dout(26));
   U52 : AOI22_X1 port map( A1 => din0(26), A2 => n35, B1 => din1(26), B2 => 
                           sel, ZN => n48);
   U53 : INV_X1 port map( A => n47, ZN => dout(27));
   U54 : AOI22_X1 port map( A1 => din0(27), A2 => n35, B1 => din1(27), B2 => 
                           sel, ZN => n47);
   U55 : AOI21_X1 port map( B1 => din1(18), B2 => sel, A => din0(18), ZN => n57
                           );
   U56 : AOI21_X1 port map( B1 => din1(19), B2 => sel, A => din0(19), ZN => n56
                           );
   U57 : AOI21_X1 port map( B1 => din1(17), B2 => sel, A => din0(17), ZN => n58
                           );
   U58 : AOI21_X1 port map( B1 => din1(15), B2 => sel, A => din0(15), ZN => n60
                           );
   U59 : AOI21_X1 port map( B1 => din1(10), B2 => sel, A => din0(10), ZN => n65
                           );
   U60 : AOI21_X1 port map( B1 => din1(11), B2 => sel, A => din0(11), ZN => n64
                           );
   U61 : AOI21_X1 port map( B1 => din1(12), B2 => sel, A => din0(12), ZN => n63
                           );
   U62 : AOI21_X1 port map( B1 => din1(13), B2 => sel, A => din0(13), ZN => n62
                           );
   U63 : AOI21_X1 port map( B1 => din1(14), B2 => sel, A => din0(14), ZN => n61
                           );
   U64 : AOI21_X1 port map( B1 => din1(16), B2 => sel, A => din0(16), ZN => n59
                           );
   U65 : AOI21_X1 port map( B1 => din1(0), B2 => sel, A => din0(0), ZN => n66);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_3 is

   port( reg_c, reg_f, reg_ff : in std_logic_vector (31 downto 0);  addr_c, 
         addr_f, addr_ff : in std_logic_vector (4 downto 0);  valid_f, valid_ff
         , dirty_f, dirty_ff, en : in std_logic;  output : out std_logic_vector
         (31 downto 0);  match_dirty_f, match_dirty_ff : out std_logic);

end FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_3;

architecture SYN_fwd_mux_2_arch of FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
      N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, 
      N106, N107, N108, N109, N110, N111, N112, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
      n72, n73, n74, n75, n76, n77, n78, n79_port, n80_port, n81_port, n82_port
      , n83_port, n84_port, n85_port, n86_port, n87_port, n88_port, n89_port, 
      n90_port, n91_port, n92_port, n93_port, n94_port, n95_port, n96_port, 
      n97_port, n98_port, n99_port, n100_port : std_logic;

begin
   
   match_dirty_ff_reg : DLH_X1 port map( G => en, D => N111, Q => 
                           match_dirty_ff);
   output_reg_31_inst : DLH_X1 port map( G => en, D => N110, Q => output(31));
   output_reg_30_inst : DLH_X1 port map( G => en, D => N109, Q => output(30));
   output_reg_29_inst : DLH_X1 port map( G => en, D => N108, Q => output(29));
   output_reg_28_inst : DLH_X1 port map( G => en, D => N107, Q => output(28));
   output_reg_27_inst : DLH_X1 port map( G => en, D => N106, Q => output(27));
   output_reg_26_inst : DLH_X1 port map( G => en, D => N105, Q => output(26));
   output_reg_25_inst : DLH_X1 port map( G => en, D => N104, Q => output(25));
   output_reg_24_inst : DLH_X1 port map( G => en, D => N103, Q => output(24));
   output_reg_23_inst : DLH_X1 port map( G => en, D => N102, Q => output(23));
   output_reg_22_inst : DLH_X1 port map( G => en, D => N101, Q => output(22));
   output_reg_21_inst : DLH_X1 port map( G => en, D => N100, Q => output(21));
   output_reg_20_inst : DLH_X1 port map( G => en, D => N99, Q => output(20));
   output_reg_19_inst : DLH_X1 port map( G => en, D => N98, Q => output(19));
   output_reg_18_inst : DLH_X1 port map( G => en, D => N97, Q => output(18));
   output_reg_17_inst : DLH_X1 port map( G => en, D => N96, Q => output(17));
   output_reg_16_inst : DLH_X1 port map( G => en, D => N95, Q => output(16));
   match_dirty_f_reg : DLH_X1 port map( G => en, D => N112, Q => match_dirty_f)
                           ;
   U83 : XOR2_X1 port map( A => addr_f(3), B => addr_c(3), Z => n85_port);
   U84 : XOR2_X1 port map( A => addr_f(2), B => addr_c(2), Z => n84_port);
   U85 : XOR2_X1 port map( A => addr_f(4), B => addr_c(4), Z => n83_port);
   U86 : XOR2_X1 port map( A => addr_ff(4), B => addr_c(4), Z => n91_port);
   U87 : XOR2_X1 port map( A => addr_ff(0), B => addr_c(0), Z => n90_port);
   U88 : XOR2_X1 port map( A => addr_ff(1), B => addr_c(1), Z => n89_port);
   U89 : XOR2_X1 port map( A => n76, B => addr_ff(3), Z => n87_port);
   U90 : XOR2_X1 port map( A => n78, B => addr_ff(2), Z => n86_port);
   output_reg_10_inst : DLH_X1 port map( G => en, D => N89, Q => output(10));
   output_reg_9_inst : DLH_X1 port map( G => en, D => N88, Q => output(9));
   output_reg_1_inst : DLH_X1 port map( G => en, D => N80, Q => output(1));
   output_reg_0_inst : DLH_X1 port map( G => en, D => N79, Q => output(0));
   output_reg_4_inst : DLH_X1 port map( G => en, D => N83, Q => output(4));
   output_reg_14_inst : DLH_X1 port map( G => en, D => N93, Q => output(14));
   output_reg_2_inst : DLH_X1 port map( G => en, D => N81, Q => output(2));
   output_reg_12_inst : DLH_X1 port map( G => en, D => N91, Q => output(12));
   output_reg_6_inst : DLH_X1 port map( G => en, D => N85, Q => output(6));
   output_reg_8_inst : DLH_X1 port map( G => en, D => N87, Q => output(8));
   output_reg_7_inst : DLH_X1 port map( G => en, D => N86, Q => output(7));
   output_reg_11_inst : DLH_X1 port map( G => en, D => N90, Q => output(11));
   output_reg_3_inst : DLH_X1 port map( G => en, D => N82, Q => output(3));
   output_reg_5_inst : DLH_X1 port map( G => en, D => N84, Q => output(5));
   output_reg_13_inst : DLH_X1 port map( G => en, D => N92, Q => output(13));
   output_reg_15_inst : DLH_X1 port map( G => en, D => N94, Q => output(15));
   U2 : BUF_X1 port map( A => n39, Z => n95_port);
   U3 : BUF_X1 port map( A => n39, Z => n96_port);
   U4 : BUF_X1 port map( A => n40, Z => n92_port);
   U5 : BUF_X1 port map( A => n40, Z => n93_port);
   U6 : BUF_X1 port map( A => n39, Z => n97_port);
   U7 : BUF_X1 port map( A => n38, Z => n99_port);
   U8 : BUF_X1 port map( A => n38, Z => n98_port);
   U9 : BUF_X1 port map( A => n40, Z => n94_port);
   U10 : BUF_X1 port map( A => n38, Z => n100_port);
   U11 : OAI21_X1 port map( B1 => n75, B2 => n72, A => n73, ZN => n38);
   U12 : AND3_X1 port map( A1 => n73, A2 => n74, A3 => n75, ZN => n39);
   U13 : AND2_X1 port map( A1 => n72, A2 => n73, ZN => n40);
   U14 : INV_X1 port map( A => n74, ZN => n72);
   U15 : NOR3_X1 port map( A1 => n83_port, A2 => n84_port, A3 => n85_port, ZN 
                           => n82_port);
   U16 : NAND4_X1 port map( A1 => n76, A2 => n77, A3 => n78, A4 => n79_port, ZN
                           => n73);
   U17 : INV_X1 port map( A => addr_c(4), ZN => n77);
   U18 : NOR2_X1 port map( A1 => addr_c(1), A2 => addr_c(0), ZN => n79_port);
   U19 : NAND4_X1 port map( A1 => n80_port, A2 => valid_f, A3 => n81_port, A4 
                           => n82_port, ZN => n74);
   U20 : XNOR2_X1 port map( A => addr_c(1), B => addr_f(1), ZN => n80_port);
   U21 : XNOR2_X1 port map( A => addr_c(0), B => addr_f(0), ZN => n81_port);
   U22 : AND4_X1 port map( A1 => n86_port, A2 => valid_ff, A3 => n87_port, A4 
                           => n88_port, ZN => n75);
   U23 : NOR3_X1 port map( A1 => n89_port, A2 => n90_port, A3 => n91_port, ZN 
                           => n88_port);
   U24 : INV_X1 port map( A => addr_c(2), ZN => n78);
   U25 : INV_X1 port map( A => addr_c(3), ZN => n76);
   U26 : INV_X1 port map( A => n51, ZN => N88);
   U27 : AOI222_X1 port map( A1 => reg_c(9), A2 => n99_port, B1 => reg_ff(9), 
                           B2 => n95_port, C1 => reg_f(9), C2 => n92_port, ZN 
                           => n51);
   U28 : INV_X1 port map( A => n59, ZN => N80);
   U29 : AOI222_X1 port map( A1 => reg_c(1), A2 => n99_port, B1 => reg_ff(1), 
                           B2 => n96_port, C1 => reg_f(1), C2 => n93_port, ZN 
                           => n59);
   U30 : INV_X1 port map( A => n60, ZN => N79);
   U31 : AOI222_X1 port map( A1 => reg_c(0), A2 => n98_port, B1 => reg_ff(0), 
                           B2 => n96_port, C1 => reg_f(0), C2 => n93_port, ZN 
                           => n60);
   U32 : INV_X1 port map( A => n58, ZN => N81);
   U33 : AOI222_X1 port map( A1 => reg_c(2), A2 => n99_port, B1 => reg_ff(2), 
                           B2 => n96_port, C1 => reg_f(2), C2 => n93_port, ZN 
                           => n58);
   U34 : INV_X1 port map( A => n55, ZN => N84);
   U35 : AOI222_X1 port map( A1 => reg_c(5), A2 => n99_port, B1 => reg_ff(5), 
                           B2 => n96_port, C1 => reg_f(5), C2 => n93_port, ZN 
                           => n55);
   U36 : INV_X1 port map( A => n52, ZN => N87);
   U37 : AOI222_X1 port map( A1 => reg_c(8), A2 => n99_port, B1 => reg_ff(8), 
                           B2 => n96_port, C1 => reg_f(8), C2 => n93_port, ZN 
                           => n52);
   U38 : INV_X1 port map( A => n50, ZN => N89);
   U39 : AOI222_X1 port map( A1 => reg_c(10), A2 => n99_port, B1 => reg_ff(10),
                           B2 => n95_port, C1 => reg_f(10), C2 => n92_port, ZN 
                           => n50);
   U40 : INV_X1 port map( A => n46, ZN => N93);
   U41 : AOI222_X1 port map( A1 => reg_c(14), A2 => n100_port, B1 => reg_ff(14)
                           , B2 => n95_port, C1 => reg_f(14), C2 => n92_port, 
                           ZN => n46);
   U42 : INV_X1 port map( A => n57, ZN => N82);
   U43 : AOI222_X1 port map( A1 => reg_c(3), A2 => n99_port, B1 => reg_ff(3), 
                           B2 => n96_port, C1 => reg_f(3), C2 => n93_port, ZN 
                           => n57);
   U44 : INV_X1 port map( A => n47, ZN => N92);
   U45 : AOI222_X1 port map( A1 => reg_c(13), A2 => n100_port, B1 => reg_ff(13)
                           , B2 => n95_port, C1 => reg_f(13), C2 => n92_port, 
                           ZN => n47);
   U46 : INV_X1 port map( A => n53, ZN => N86);
   U47 : AOI222_X1 port map( A1 => reg_c(7), A2 => n99_port, B1 => reg_ff(7), 
                           B2 => n96_port, C1 => reg_f(7), C2 => n93_port, ZN 
                           => n53);
   U48 : INV_X1 port map( A => n45, ZN => N94);
   U49 : AOI222_X1 port map( A1 => reg_c(15), A2 => n100_port, B1 => reg_ff(15)
                           , B2 => n95_port, C1 => reg_f(15), C2 => n92_port, 
                           ZN => n45);
   U50 : INV_X1 port map( A => n49, ZN => N90);
   U51 : AOI222_X1 port map( A1 => reg_c(11), A2 => n99_port, B1 => reg_ff(11),
                           B2 => n95_port, C1 => reg_f(11), C2 => n92_port, ZN 
                           => n49);
   U52 : INV_X1 port map( A => n54, ZN => N85);
   U53 : AOI222_X1 port map( A1 => reg_c(6), A2 => n99_port, B1 => reg_ff(6), 
                           B2 => n96_port, C1 => reg_f(6), C2 => n93_port, ZN 
                           => n54);
   U54 : INV_X1 port map( A => n56, ZN => N83);
   U55 : AOI222_X1 port map( A1 => reg_c(4), A2 => n99_port, B1 => reg_ff(4), 
                           B2 => n96_port, C1 => reg_f(4), C2 => n93_port, ZN 
                           => n56);
   U56 : INV_X1 port map( A => n48, ZN => N91);
   U57 : AOI222_X1 port map( A1 => reg_c(12), A2 => n99_port, B1 => reg_ff(12),
                           B2 => n95_port, C1 => reg_f(12), C2 => n92_port, ZN 
                           => n48);
   U58 : INV_X1 port map( A => n70, ZN => N101);
   U59 : AOI222_X1 port map( A1 => reg_c(22), A2 => n98_port, B1 => reg_ff(22),
                           B2 => n97_port, C1 => reg_f(22), C2 => n94_port, ZN 
                           => n70);
   U60 : INV_X1 port map( A => n69, ZN => N102);
   U61 : AOI222_X1 port map( A1 => reg_c(23), A2 => n98_port, B1 => reg_ff(23),
                           B2 => n97_port, C1 => reg_f(23), C2 => n94_port, ZN 
                           => n69);
   U62 : INV_X1 port map( A => n68, ZN => N103);
   U63 : AOI222_X1 port map( A1 => reg_c(24), A2 => n98_port, B1 => reg_ff(24),
                           B2 => n97_port, C1 => reg_f(24), C2 => n94_port, ZN 
                           => n68);
   U64 : INV_X1 port map( A => n67, ZN => N104);
   U65 : AOI222_X1 port map( A1 => reg_c(25), A2 => n98_port, B1 => reg_ff(25),
                           B2 => n97_port, C1 => reg_f(25), C2 => n94_port, ZN 
                           => n67);
   U66 : INV_X1 port map( A => n66, ZN => N105);
   U67 : AOI222_X1 port map( A1 => reg_c(26), A2 => n98_port, B1 => reg_ff(26),
                           B2 => n97_port, C1 => reg_f(26), C2 => n94_port, ZN 
                           => n66);
   U68 : INV_X1 port map( A => n65, ZN => N106);
   U69 : AOI222_X1 port map( A1 => reg_c(27), A2 => n98_port, B1 => reg_ff(27),
                           B2 => n97_port, C1 => reg_f(27), C2 => n94_port, ZN 
                           => n65);
   U70 : INV_X1 port map( A => n64, ZN => N107);
   U71 : AOI222_X1 port map( A1 => reg_c(28), A2 => n98_port, B1 => reg_ff(28),
                           B2 => n97_port, C1 => reg_f(28), C2 => n94_port, ZN 
                           => n64);
   U72 : INV_X1 port map( A => n63, ZN => N108);
   U73 : AOI222_X1 port map( A1 => reg_c(29), A2 => n98_port, B1 => reg_ff(29),
                           B2 => n97_port, C1 => reg_f(29), C2 => n94_port, ZN 
                           => n63);
   U74 : INV_X1 port map( A => n44, ZN => N95);
   U75 : AOI222_X1 port map( A1 => reg_c(16), A2 => n100_port, B1 => reg_ff(16)
                           , B2 => n95_port, C1 => reg_f(16), C2 => n92_port, 
                           ZN => n44);
   U76 : INV_X1 port map( A => n43, ZN => N96);
   U77 : AOI222_X1 port map( A1 => reg_c(17), A2 => n100_port, B1 => reg_ff(17)
                           , B2 => n95_port, C1 => reg_f(17), C2 => n92_port, 
                           ZN => n43);
   U78 : INV_X1 port map( A => n42, ZN => N97);
   U79 : AOI222_X1 port map( A1 => reg_c(18), A2 => n100_port, B1 => reg_ff(18)
                           , B2 => n95_port, C1 => reg_f(18), C2 => n92_port, 
                           ZN => n42);
   U80 : INV_X1 port map( A => n41, ZN => N98);
   U81 : AOI222_X1 port map( A1 => reg_c(19), A2 => n100_port, B1 => reg_ff(19)
                           , B2 => n95_port, C1 => reg_f(19), C2 => n92_port, 
                           ZN => n41);
   U82 : INV_X1 port map( A => n37, ZN => N99);
   U91 : AOI222_X1 port map( A1 => reg_c(20), A2 => n100_port, B1 => reg_ff(20)
                           , B2 => n96_port, C1 => reg_f(20), C2 => n93_port, 
                           ZN => n37);
   U92 : INV_X1 port map( A => n71, ZN => N100);
   U93 : AOI222_X1 port map( A1 => reg_c(21), A2 => n98_port, B1 => reg_ff(21),
                           B2 => n95_port, C1 => reg_f(21), C2 => n92_port, ZN 
                           => n71);
   U94 : INV_X1 port map( A => n62, ZN => N109);
   U95 : AOI222_X1 port map( A1 => reg_c(30), A2 => n98_port, B1 => reg_ff(30),
                           B2 => n96_port, C1 => reg_f(30), C2 => n93_port, ZN 
                           => n62);
   U96 : INV_X1 port map( A => n61, ZN => N110);
   U97 : AOI222_X1 port map( A1 => reg_c(31), A2 => n98_port, B1 => reg_ff(31),
                           B2 => n96_port, C1 => reg_f(31), C2 => n93_port, ZN 
                           => n61);
   U98 : AND2_X1 port map( A1 => dirty_ff, A2 => n97_port, ZN => N111);
   U99 : AND2_X1 port map( A1 => dirty_f, A2 => n94_port, ZN => N112);

end SYN_fwd_mux_2_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE5_6 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 0); 
         dout : out std_logic_vector (4 downto 0));

end Reg_DATA_SIZE5_6;

architecture SYN_reg_arch of Reg_DATA_SIZE5_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, net109193, net109194, net109195, net109196, 
      net109197, n6, n7, n8, n9, n10 : std_logic;

begin
   
   dout_reg_4_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           dout(4), QN => net109197);
   dout_reg_3_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           dout(3), QN => net109196);
   dout_reg_2_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           dout(2), QN => net109195);
   dout_reg_1_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           dout(1), QN => net109194);
   dout_reg_0_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           dout(0), QN => net109193);
   U2 : OAI21_X1 port map( B1 => net109193, B2 => en, A => n6, ZN => n5);
   U3 : NAND2_X1 port map( A1 => en, A2 => din(0), ZN => n6);
   U4 : OAI21_X1 port map( B1 => net109194, B2 => en, A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => din(1), A2 => en, ZN => n7);
   U6 : OAI21_X1 port map( B1 => net109195, B2 => en, A => n8, ZN => n3);
   U7 : NAND2_X1 port map( A1 => din(2), A2 => en, ZN => n8);
   U8 : OAI21_X1 port map( B1 => net109196, B2 => en, A => n9, ZN => n2);
   U9 : NAND2_X1 port map( A1 => din(3), A2 => en, ZN => n9);
   U10 : OAI21_X1 port map( B1 => net109197, B2 => en, A => n10, ZN => n1);
   U11 : NAND2_X1 port map( A1 => din(4), A2 => en, ZN => n10);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE5_0 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 0); 
         dout : out std_logic_vector (4 downto 0));

end Reg_DATA_SIZE5_0;

architecture SYN_reg_arch of Reg_DATA_SIZE5_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n11, n12, n13, n14, n15, net108611, net108612, net108613, net108614, 
      net108615, n1, n2, n3, n4, n5 : std_logic;

begin
   
   dout_reg_4_inst : DFFR_X1 port map( D => n15, CK => clk, RN => rst, Q => 
                           dout(4), QN => net108615);
   dout_reg_3_inst : DFFR_X1 port map( D => n14, CK => clk, RN => rst, Q => 
                           dout(3), QN => net108614);
   dout_reg_2_inst : DFFR_X1 port map( D => n13, CK => clk, RN => rst, Q => 
                           dout(2), QN => net108613);
   dout_reg_1_inst : DFFR_X1 port map( D => n12, CK => clk, RN => rst, Q => 
                           dout(1), QN => net108612);
   dout_reg_0_inst : DFFR_X1 port map( D => n11, CK => clk, RN => rst, Q => 
                           dout(0), QN => net108611);
   U2 : OAI21_X1 port map( B1 => net108611, B2 => en, A => n5, ZN => n11);
   U3 : NAND2_X1 port map( A1 => din(0), A2 => en, ZN => n5);
   U4 : OAI21_X1 port map( B1 => net108612, B2 => en, A => n4, ZN => n12);
   U5 : NAND2_X1 port map( A1 => din(1), A2 => en, ZN => n4);
   U6 : OAI21_X1 port map( B1 => net108613, B2 => en, A => n3, ZN => n13);
   U7 : NAND2_X1 port map( A1 => din(2), A2 => en, ZN => n3);
   U8 : OAI21_X1 port map( B1 => net108614, B2 => en, A => n2, ZN => n14);
   U9 : NAND2_X1 port map( A1 => din(3), A2 => en, ZN => n2);
   U10 : OAI21_X1 port map( B1 => net108615, B2 => en, A => n1, ZN => n15);
   U11 : NAND2_X1 port map( A1 => en, A2 => din(4), ZN => n1);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_4 is

   port( reg_c, reg_f, reg_ff : in std_logic_vector (31 downto 0);  addr_c, 
         addr_f, addr_ff : in std_logic_vector (4 downto 0);  valid_f, valid_ff
         , dirty_f, dirty_ff, en : in std_logic;  output : out std_logic_vector
         (31 downto 0);  match_dirty_f, match_dirty_ff : out std_logic);

end FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_4;

architecture SYN_fwd_mux_2_arch of FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_4 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
      N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, 
      N106, N107, N108, N109, N110, N111, N112, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
      n72, n73, n74, n75, n76, n77, n78, n79_port, n80_port, n81_port, n82_port
      , n83_port, n84_port, n85_port, n86_port, n87_port, n88_port, n89_port, 
      n90_port, n91_port, n92_port, n93_port, n94_port, n95_port, n96_port, 
      n97_port, n98_port, n99_port, n100_port : std_logic;

begin
   
   match_dirty_ff_reg : DLH_X1 port map( G => en, D => N111, Q => 
                           match_dirty_ff);
   output_reg_31_inst : DLH_X1 port map( G => en, D => N110, Q => output(31));
   output_reg_30_inst : DLH_X1 port map( G => en, D => N109, Q => output(30));
   output_reg_29_inst : DLH_X1 port map( G => en, D => N108, Q => output(29));
   output_reg_28_inst : DLH_X1 port map( G => en, D => N107, Q => output(28));
   output_reg_27_inst : DLH_X1 port map( G => en, D => N106, Q => output(27));
   output_reg_26_inst : DLH_X1 port map( G => en, D => N105, Q => output(26));
   output_reg_25_inst : DLH_X1 port map( G => en, D => N104, Q => output(25));
   output_reg_24_inst : DLH_X1 port map( G => en, D => N103, Q => output(24));
   output_reg_23_inst : DLH_X1 port map( G => en, D => N102, Q => output(23));
   output_reg_22_inst : DLH_X1 port map( G => en, D => N101, Q => output(22));
   output_reg_21_inst : DLH_X1 port map( G => en, D => N100, Q => output(21));
   output_reg_20_inst : DLH_X1 port map( G => en, D => N99, Q => output(20));
   output_reg_19_inst : DLH_X1 port map( G => en, D => N98, Q => output(19));
   output_reg_18_inst : DLH_X1 port map( G => en, D => N97, Q => output(18));
   output_reg_17_inst : DLH_X1 port map( G => en, D => N96, Q => output(17));
   output_reg_16_inst : DLH_X1 port map( G => en, D => N95, Q => output(16));
   output_reg_15_inst : DLH_X1 port map( G => en, D => N94, Q => output(15));
   output_reg_14_inst : DLH_X1 port map( G => en, D => N93, Q => output(14));
   output_reg_13_inst : DLH_X1 port map( G => en, D => N92, Q => output(13));
   output_reg_12_inst : DLH_X1 port map( G => en, D => N91, Q => output(12));
   output_reg_11_inst : DLH_X1 port map( G => en, D => N90, Q => output(11));
   output_reg_10_inst : DLH_X1 port map( G => en, D => N89, Q => output(10));
   output_reg_9_inst : DLH_X1 port map( G => en, D => N88, Q => output(9));
   output_reg_8_inst : DLH_X1 port map( G => en, D => N87, Q => output(8));
   output_reg_7_inst : DLH_X1 port map( G => en, D => N86, Q => output(7));
   output_reg_6_inst : DLH_X1 port map( G => en, D => N85, Q => output(6));
   output_reg_5_inst : DLH_X1 port map( G => en, D => N84, Q => output(5));
   output_reg_4_inst : DLH_X1 port map( G => en, D => N83, Q => output(4));
   output_reg_3_inst : DLH_X1 port map( G => en, D => N82, Q => output(3));
   output_reg_2_inst : DLH_X1 port map( G => en, D => N81, Q => output(2));
   output_reg_1_inst : DLH_X1 port map( G => en, D => N80, Q => output(1));
   output_reg_0_inst : DLH_X1 port map( G => en, D => N79, Q => output(0));
   match_dirty_f_reg : DLH_X1 port map( G => en, D => N112, Q => match_dirty_f)
                           ;
   U83 : XOR2_X1 port map( A => addr_f(3), B => addr_c(3), Z => n85_port);
   U84 : XOR2_X1 port map( A => addr_f(2), B => addr_c(2), Z => n84_port);
   U85 : XOR2_X1 port map( A => addr_f(4), B => addr_c(4), Z => n83_port);
   U86 : XOR2_X1 port map( A => addr_ff(4), B => addr_c(4), Z => n91_port);
   U87 : XOR2_X1 port map( A => addr_ff(0), B => addr_c(0), Z => n90_port);
   U88 : XOR2_X1 port map( A => addr_ff(1), B => addr_c(1), Z => n89_port);
   U89 : XOR2_X1 port map( A => n76, B => addr_ff(3), Z => n87_port);
   U90 : XOR2_X1 port map( A => n78, B => addr_ff(2), Z => n86_port);
   U2 : BUF_X1 port map( A => n39, Z => n95_port);
   U3 : BUF_X1 port map( A => n40, Z => n92_port);
   U4 : BUF_X1 port map( A => n39, Z => n97_port);
   U5 : BUF_X1 port map( A => n39, Z => n96_port);
   U6 : BUF_X1 port map( A => n38, Z => n99_port);
   U7 : BUF_X1 port map( A => n40, Z => n94_port);
   U8 : BUF_X1 port map( A => n40, Z => n93_port);
   U9 : BUF_X1 port map( A => n38, Z => n98_port);
   U10 : BUF_X1 port map( A => n38, Z => n100_port);
   U11 : OAI21_X1 port map( B1 => n75, B2 => n72, A => n73, ZN => n38);
   U12 : AND3_X1 port map( A1 => n73, A2 => n74, A3 => n75, ZN => n39);
   U13 : AND2_X1 port map( A1 => n72, A2 => n73, ZN => n40);
   U14 : INV_X1 port map( A => n74, ZN => n72);
   U15 : NOR3_X1 port map( A1 => n83_port, A2 => n84_port, A3 => n85_port, ZN 
                           => n82_port);
   U16 : NAND4_X1 port map( A1 => n76, A2 => n77, A3 => n78, A4 => n79_port, ZN
                           => n73);
   U17 : INV_X1 port map( A => addr_c(4), ZN => n77);
   U18 : NOR2_X1 port map( A1 => addr_c(1), A2 => addr_c(0), ZN => n79_port);
   U19 : NAND4_X1 port map( A1 => n80_port, A2 => valid_f, A3 => n81_port, A4 
                           => n82_port, ZN => n74);
   U20 : XNOR2_X1 port map( A => addr_c(1), B => addr_f(1), ZN => n80_port);
   U21 : XNOR2_X1 port map( A => addr_c(0), B => addr_f(0), ZN => n81_port);
   U22 : INV_X1 port map( A => n60, ZN => N79);
   U23 : AND4_X1 port map( A1 => n86_port, A2 => valid_ff, A3 => n87_port, A4 
                           => n88_port, ZN => n75);
   U24 : NOR3_X1 port map( A1 => n89_port, A2 => n90_port, A3 => n91_port, ZN 
                           => n88_port);
   U25 : INV_X1 port map( A => addr_c(2), ZN => n78);
   U26 : INV_X1 port map( A => n70, ZN => N101);
   U27 : AOI222_X1 port map( A1 => reg_c(22), A2 => n98_port, B1 => reg_ff(22),
                           B2 => n97_port, C1 => reg_f(22), C2 => n94_port, ZN 
                           => n70);
   U28 : INV_X1 port map( A => n69, ZN => N102);
   U29 : AOI222_X1 port map( A1 => reg_c(23), A2 => n98_port, B1 => reg_ff(23),
                           B2 => n97_port, C1 => reg_f(23), C2 => n94_port, ZN 
                           => n69);
   U30 : INV_X1 port map( A => n68, ZN => N103);
   U31 : AOI222_X1 port map( A1 => reg_c(24), A2 => n98_port, B1 => reg_ff(24),
                           B2 => n97_port, C1 => reg_f(24), C2 => n94_port, ZN 
                           => n68);
   U32 : INV_X1 port map( A => n67, ZN => N104);
   U33 : AOI222_X1 port map( A1 => reg_c(25), A2 => n98_port, B1 => reg_ff(25),
                           B2 => n97_port, C1 => reg_f(25), C2 => n94_port, ZN 
                           => n67);
   U34 : INV_X1 port map( A => n66, ZN => N105);
   U35 : AOI222_X1 port map( A1 => reg_c(26), A2 => n98_port, B1 => reg_ff(26),
                           B2 => n97_port, C1 => reg_f(26), C2 => n94_port, ZN 
                           => n66);
   U36 : INV_X1 port map( A => n65, ZN => N106);
   U37 : AOI222_X1 port map( A1 => reg_c(27), A2 => n98_port, B1 => reg_ff(27),
                           B2 => n97_port, C1 => reg_f(27), C2 => n94_port, ZN 
                           => n65);
   U38 : INV_X1 port map( A => n64, ZN => N107);
   U39 : AOI222_X1 port map( A1 => reg_c(28), A2 => n98_port, B1 => reg_ff(28),
                           B2 => n97_port, C1 => reg_f(28), C2 => n94_port, ZN 
                           => n64);
   U40 : INV_X1 port map( A => n63, ZN => N108);
   U41 : AOI222_X1 port map( A1 => reg_c(29), A2 => n98_port, B1 => reg_ff(29),
                           B2 => n97_port, C1 => reg_f(29), C2 => n94_port, ZN 
                           => n63);
   U42 : INV_X1 port map( A => n59, ZN => N80);
   U43 : AOI222_X1 port map( A1 => reg_c(1), A2 => n99_port, B1 => reg_ff(1), 
                           B2 => n96_port, C1 => reg_f(1), C2 => n93_port, ZN 
                           => n59);
   U44 : INV_X1 port map( A => n58, ZN => N81);
   U45 : AOI222_X1 port map( A1 => reg_c(2), A2 => n99_port, B1 => reg_ff(2), 
                           B2 => n96_port, C1 => reg_f(2), C2 => n93_port, ZN 
                           => n58);
   U46 : INV_X1 port map( A => n57, ZN => N82);
   U47 : AOI222_X1 port map( A1 => reg_c(3), A2 => n99_port, B1 => reg_ff(3), 
                           B2 => n96_port, C1 => reg_f(3), C2 => n93_port, ZN 
                           => n57);
   U48 : INV_X1 port map( A => n56, ZN => N83);
   U49 : AOI222_X1 port map( A1 => reg_c(4), A2 => n99_port, B1 => reg_ff(4), 
                           B2 => n96_port, C1 => reg_f(4), C2 => n93_port, ZN 
                           => n56);
   U50 : INV_X1 port map( A => n55, ZN => N84);
   U51 : AOI222_X1 port map( A1 => reg_c(5), A2 => n99_port, B1 => reg_ff(5), 
                           B2 => n96_port, C1 => reg_f(5), C2 => n93_port, ZN 
                           => n55);
   U52 : INV_X1 port map( A => n54, ZN => N85);
   U53 : AOI222_X1 port map( A1 => reg_c(6), A2 => n99_port, B1 => reg_ff(6), 
                           B2 => n96_port, C1 => reg_f(6), C2 => n93_port, ZN 
                           => n54);
   U54 : INV_X1 port map( A => n53, ZN => N86);
   U55 : AOI222_X1 port map( A1 => reg_c(7), A2 => n99_port, B1 => reg_ff(7), 
                           B2 => n96_port, C1 => reg_f(7), C2 => n93_port, ZN 
                           => n53);
   U56 : INV_X1 port map( A => n52, ZN => N87);
   U57 : AOI222_X1 port map( A1 => reg_c(8), A2 => n99_port, B1 => reg_ff(8), 
                           B2 => n96_port, C1 => reg_f(8), C2 => n93_port, ZN 
                           => n52);
   U58 : INV_X1 port map( A => n51, ZN => N88);
   U59 : AOI222_X1 port map( A1 => reg_c(9), A2 => n99_port, B1 => reg_ff(9), 
                           B2 => n95_port, C1 => reg_f(9), C2 => n92_port, ZN 
                           => n51);
   U60 : INV_X1 port map( A => n50, ZN => N89);
   U61 : AOI222_X1 port map( A1 => reg_c(10), A2 => n99_port, B1 => reg_ff(10),
                           B2 => n95_port, C1 => reg_f(10), C2 => n92_port, ZN 
                           => n50);
   U62 : INV_X1 port map( A => n49, ZN => N90);
   U63 : AOI222_X1 port map( A1 => reg_c(11), A2 => n99_port, B1 => reg_ff(11),
                           B2 => n95_port, C1 => reg_f(11), C2 => n92_port, ZN 
                           => n49);
   U64 : INV_X1 port map( A => n48, ZN => N91);
   U65 : AOI222_X1 port map( A1 => reg_c(12), A2 => n99_port, B1 => reg_ff(12),
                           B2 => n95_port, C1 => reg_f(12), C2 => n92_port, ZN 
                           => n48);
   U66 : INV_X1 port map( A => n47, ZN => N92);
   U67 : AOI222_X1 port map( A1 => reg_c(13), A2 => n100_port, B1 => reg_ff(13)
                           , B2 => n95_port, C1 => reg_f(13), C2 => n92_port, 
                           ZN => n47);
   U68 : INV_X1 port map( A => n46, ZN => N93);
   U69 : AOI222_X1 port map( A1 => reg_c(14), A2 => n100_port, B1 => reg_ff(14)
                           , B2 => n95_port, C1 => reg_f(14), C2 => n92_port, 
                           ZN => n46);
   U70 : INV_X1 port map( A => n45, ZN => N94);
   U71 : AOI222_X1 port map( A1 => reg_c(15), A2 => n100_port, B1 => reg_ff(15)
                           , B2 => n95_port, C1 => reg_f(15), C2 => n92_port, 
                           ZN => n45);
   U72 : INV_X1 port map( A => n44, ZN => N95);
   U73 : AOI222_X1 port map( A1 => reg_c(16), A2 => n100_port, B1 => reg_ff(16)
                           , B2 => n95_port, C1 => reg_f(16), C2 => n92_port, 
                           ZN => n44);
   U74 : INV_X1 port map( A => n43, ZN => N96);
   U75 : AOI222_X1 port map( A1 => reg_c(17), A2 => n100_port, B1 => reg_ff(17)
                           , B2 => n95_port, C1 => reg_f(17), C2 => n92_port, 
                           ZN => n43);
   U76 : INV_X1 port map( A => n42, ZN => N97);
   U77 : AOI222_X1 port map( A1 => reg_c(18), A2 => n100_port, B1 => reg_ff(18)
                           , B2 => n95_port, C1 => reg_f(18), C2 => n92_port, 
                           ZN => n42);
   U78 : INV_X1 port map( A => n41, ZN => N98);
   U79 : AOI222_X1 port map( A1 => reg_c(19), A2 => n100_port, B1 => reg_ff(19)
                           , B2 => n95_port, C1 => reg_f(19), C2 => n92_port, 
                           ZN => n41);
   U80 : INV_X1 port map( A => n37, ZN => N99);
   U81 : AOI222_X1 port map( A1 => reg_c(20), A2 => n100_port, B1 => reg_ff(20)
                           , B2 => n96_port, C1 => reg_f(20), C2 => n93_port, 
                           ZN => n37);
   U82 : INV_X1 port map( A => n71, ZN => N100);
   U91 : AOI222_X1 port map( A1 => reg_c(21), A2 => n98_port, B1 => reg_ff(21),
                           B2 => n95_port, C1 => reg_f(21), C2 => n92_port, ZN 
                           => n71);
   U92 : INV_X1 port map( A => n62, ZN => N109);
   U93 : AOI222_X1 port map( A1 => reg_c(30), A2 => n98_port, B1 => reg_ff(30),
                           B2 => n96_port, C1 => reg_f(30), C2 => n93_port, ZN 
                           => n62);
   U94 : INV_X1 port map( A => n61, ZN => N110);
   U95 : AOI222_X1 port map( A1 => reg_c(31), A2 => n98_port, B1 => reg_ff(31),
                           B2 => n96_port, C1 => reg_f(31), C2 => n93_port, ZN 
                           => n61);
   U96 : INV_X1 port map( A => addr_c(3), ZN => n76);
   U97 : AND2_X1 port map( A1 => dirty_ff, A2 => n97_port, ZN => N111);
   U98 : AND2_X1 port map( A1 => dirty_f, A2 => n94_port, ZN => N112);
   U99 : AOI222_X1 port map( A1 => reg_c(0), A2 => n98_port, B1 => reg_ff(0), 
                           B2 => n96_port, C1 => reg_f(0), C2 => n93_port, ZN 
                           => n60);

end SYN_fwd_mux_2_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_0 is

   port( reg_c, reg_f, reg_ff : in std_logic_vector (31 downto 0);  addr_c, 
         addr_f, addr_ff : in std_logic_vector (4 downto 0);  valid_f, valid_ff
         , dirty_f, dirty_ff, en : in std_logic;  output : out std_logic_vector
         (31 downto 0);  match_dirty_f, match_dirty_ff : out std_logic);

end FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_0;

architecture SYN_fwd_mux_2_arch of FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_0 is

   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
      N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, 
      N106, N107, N108, N109, N110, N111, N112, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
      n72, n73, n74, n75, n76, n77, n78, n79_port, n80_port, n81_port, n82_port
      , n83_port, n84_port, n85_port, n86_port, n87_port, n88_port, n89_port, 
      n90_port, n91_port, n92_port, n93_port, n94_port, n95_port, n96_port, 
      n97_port, n98_port, n99_port, n100_port : std_logic;

begin
   
   match_dirty_ff_reg : DLH_X1 port map( G => en, D => N111, Q => 
                           match_dirty_ff);
   output_reg_31_inst : DLH_X1 port map( G => en, D => N110, Q => output(31));
   output_reg_30_inst : DLH_X1 port map( G => en, D => N109, Q => output(30));
   output_reg_29_inst : DLH_X1 port map( G => en, D => N108, Q => output(29));
   output_reg_28_inst : DLH_X1 port map( G => en, D => N107, Q => output(28));
   output_reg_27_inst : DLH_X1 port map( G => en, D => N106, Q => output(27));
   output_reg_26_inst : DLH_X1 port map( G => en, D => N105, Q => output(26));
   output_reg_25_inst : DLH_X1 port map( G => en, D => N104, Q => output(25));
   output_reg_24_inst : DLH_X1 port map( G => en, D => N103, Q => output(24));
   output_reg_23_inst : DLH_X1 port map( G => en, D => N102, Q => output(23));
   output_reg_22_inst : DLH_X1 port map( G => en, D => N101, Q => output(22));
   output_reg_21_inst : DLH_X1 port map( G => en, D => N100, Q => output(21));
   output_reg_20_inst : DLH_X1 port map( G => en, D => N99, Q => output(20));
   output_reg_19_inst : DLH_X1 port map( G => en, D => N98, Q => output(19));
   output_reg_18_inst : DLH_X1 port map( G => en, D => N97, Q => output(18));
   output_reg_17_inst : DLH_X1 port map( G => en, D => N96, Q => output(17));
   output_reg_16_inst : DLH_X1 port map( G => en, D => N95, Q => output(16));
   output_reg_15_inst : DLH_X1 port map( G => en, D => N94, Q => output(15));
   output_reg_14_inst : DLH_X1 port map( G => en, D => N93, Q => output(14));
   output_reg_13_inst : DLH_X1 port map( G => en, D => N92, Q => output(13));
   output_reg_12_inst : DLH_X1 port map( G => en, D => N91, Q => output(12));
   output_reg_11_inst : DLH_X1 port map( G => en, D => N90, Q => output(11));
   output_reg_10_inst : DLH_X1 port map( G => en, D => N89, Q => output(10));
   output_reg_9_inst : DLH_X1 port map( G => en, D => N88, Q => output(9));
   output_reg_8_inst : DLH_X1 port map( G => en, D => N87, Q => output(8));
   output_reg_7_inst : DLH_X1 port map( G => en, D => N86, Q => output(7));
   output_reg_6_inst : DLH_X1 port map( G => en, D => N85, Q => output(6));
   output_reg_5_inst : DLH_X1 port map( G => en, D => N84, Q => output(5));
   output_reg_4_inst : DLH_X1 port map( G => en, D => N83, Q => output(4));
   output_reg_3_inst : DLH_X1 port map( G => en, D => N82, Q => output(3));
   output_reg_2_inst : DLH_X1 port map( G => en, D => N81, Q => output(2));
   output_reg_1_inst : DLH_X1 port map( G => en, D => N80, Q => output(1));
   output_reg_0_inst : DLH_X1 port map( G => en, D => N79, Q => output(0));
   U83 : XOR2_X1 port map( A => addr_f(3), B => addr_c(3), Z => n85_port);
   U84 : XOR2_X1 port map( A => addr_f(2), B => addr_c(2), Z => n84_port);
   U85 : XOR2_X1 port map( A => addr_f(4), B => addr_c(4), Z => n83_port);
   U86 : XOR2_X1 port map( A => addr_ff(4), B => addr_c(4), Z => n91_port);
   U87 : XOR2_X1 port map( A => addr_ff(0), B => addr_c(0), Z => n90_port);
   U88 : XOR2_X1 port map( A => addr_ff(1), B => addr_c(1), Z => n89_port);
   U89 : XOR2_X1 port map( A => n76, B => addr_ff(3), Z => n87_port);
   U90 : XOR2_X1 port map( A => n78, B => addr_ff(2), Z => n86_port);
   match_dirty_f_reg : DLH_X1 port map( G => en, D => N112, Q => match_dirty_f)
                           ;
   U2 : BUF_X1 port map( A => n39, Z => n95_port);
   U3 : BUF_X1 port map( A => n40, Z => n92_port);
   U4 : BUF_X1 port map( A => n39, Z => n97_port);
   U5 : BUF_X1 port map( A => n39, Z => n96_port);
   U6 : BUF_X1 port map( A => n38, Z => n99_port);
   U7 : BUF_X1 port map( A => n40, Z => n94_port);
   U8 : BUF_X1 port map( A => n40, Z => n93_port);
   U9 : BUF_X1 port map( A => n38, Z => n98_port);
   U10 : BUF_X1 port map( A => n38, Z => n100_port);
   U11 : OAI21_X1 port map( B1 => n75, B2 => n72, A => n73, ZN => n38);
   U12 : AND3_X1 port map( A1 => n73, A2 => n74, A3 => n75, ZN => n39);
   U13 : AND2_X1 port map( A1 => n72, A2 => n73, ZN => n40);
   U14 : INV_X1 port map( A => n74, ZN => n72);
   U15 : NOR3_X1 port map( A1 => n83_port, A2 => n84_port, A3 => n85_port, ZN 
                           => n82_port);
   U16 : NAND4_X1 port map( A1 => n76, A2 => n77, A3 => n78, A4 => n79_port, ZN
                           => n73);
   U17 : INV_X1 port map( A => addr_c(4), ZN => n77);
   U18 : NOR2_X1 port map( A1 => addr_c(1), A2 => addr_c(0), ZN => n79_port);
   U19 : NAND4_X1 port map( A1 => n80_port, A2 => valid_f, A3 => n81_port, A4 
                           => n82_port, ZN => n74);
   U20 : XNOR2_X1 port map( A => addr_c(1), B => addr_f(1), ZN => n80_port);
   U21 : XNOR2_X1 port map( A => addr_c(0), B => addr_f(0), ZN => n81_port);
   U22 : INV_X1 port map( A => n60, ZN => N79);
   U23 : AND4_X1 port map( A1 => n86_port, A2 => valid_ff, A3 => n87_port, A4 
                           => n88_port, ZN => n75);
   U24 : NOR3_X1 port map( A1 => n89_port, A2 => n90_port, A3 => n91_port, ZN 
                           => n88_port);
   U25 : INV_X1 port map( A => addr_c(2), ZN => n78);
   U26 : INV_X1 port map( A => n70, ZN => N101);
   U27 : AOI222_X1 port map( A1 => reg_c(22), A2 => n98_port, B1 => reg_ff(22),
                           B2 => n97_port, C1 => reg_f(22), C2 => n94_port, ZN 
                           => n70);
   U28 : INV_X1 port map( A => n69, ZN => N102);
   U29 : AOI222_X1 port map( A1 => reg_c(23), A2 => n98_port, B1 => reg_ff(23),
                           B2 => n97_port, C1 => reg_f(23), C2 => n94_port, ZN 
                           => n69);
   U30 : INV_X1 port map( A => n68, ZN => N103);
   U31 : AOI222_X1 port map( A1 => reg_c(24), A2 => n98_port, B1 => reg_ff(24),
                           B2 => n97_port, C1 => reg_f(24), C2 => n94_port, ZN 
                           => n68);
   U32 : INV_X1 port map( A => n67, ZN => N104);
   U33 : AOI222_X1 port map( A1 => reg_c(25), A2 => n98_port, B1 => reg_ff(25),
                           B2 => n97_port, C1 => reg_f(25), C2 => n94_port, ZN 
                           => n67);
   U34 : INV_X1 port map( A => n66, ZN => N105);
   U35 : AOI222_X1 port map( A1 => reg_c(26), A2 => n98_port, B1 => reg_ff(26),
                           B2 => n97_port, C1 => reg_f(26), C2 => n94_port, ZN 
                           => n66);
   U36 : INV_X1 port map( A => n65, ZN => N106);
   U37 : AOI222_X1 port map( A1 => reg_c(27), A2 => n98_port, B1 => reg_ff(27),
                           B2 => n97_port, C1 => reg_f(27), C2 => n94_port, ZN 
                           => n65);
   U38 : INV_X1 port map( A => n64, ZN => N107);
   U39 : AOI222_X1 port map( A1 => reg_c(28), A2 => n98_port, B1 => reg_ff(28),
                           B2 => n97_port, C1 => reg_f(28), C2 => n94_port, ZN 
                           => n64);
   U40 : INV_X1 port map( A => n63, ZN => N108);
   U41 : AOI222_X1 port map( A1 => reg_c(29), A2 => n98_port, B1 => reg_ff(29),
                           B2 => n97_port, C1 => reg_f(29), C2 => n94_port, ZN 
                           => n63);
   U42 : INV_X1 port map( A => n59, ZN => N80);
   U43 : AOI222_X1 port map( A1 => reg_c(1), A2 => n99_port, B1 => reg_ff(1), 
                           B2 => n96_port, C1 => reg_f(1), C2 => n93_port, ZN 
                           => n59);
   U44 : INV_X1 port map( A => n58, ZN => N81);
   U45 : AOI222_X1 port map( A1 => reg_c(2), A2 => n99_port, B1 => reg_ff(2), 
                           B2 => n96_port, C1 => reg_f(2), C2 => n93_port, ZN 
                           => n58);
   U46 : INV_X1 port map( A => n57, ZN => N82);
   U47 : AOI222_X1 port map( A1 => reg_c(3), A2 => n99_port, B1 => reg_ff(3), 
                           B2 => n96_port, C1 => reg_f(3), C2 => n93_port, ZN 
                           => n57);
   U48 : INV_X1 port map( A => n56, ZN => N83);
   U49 : AOI222_X1 port map( A1 => reg_c(4), A2 => n99_port, B1 => reg_ff(4), 
                           B2 => n96_port, C1 => reg_f(4), C2 => n93_port, ZN 
                           => n56);
   U50 : INV_X1 port map( A => n55, ZN => N84);
   U51 : AOI222_X1 port map( A1 => reg_c(5), A2 => n99_port, B1 => reg_ff(5), 
                           B2 => n96_port, C1 => reg_f(5), C2 => n93_port, ZN 
                           => n55);
   U52 : INV_X1 port map( A => n54, ZN => N85);
   U53 : AOI222_X1 port map( A1 => reg_c(6), A2 => n99_port, B1 => reg_ff(6), 
                           B2 => n96_port, C1 => reg_f(6), C2 => n93_port, ZN 
                           => n54);
   U54 : INV_X1 port map( A => n53, ZN => N86);
   U55 : AOI222_X1 port map( A1 => reg_c(7), A2 => n99_port, B1 => reg_ff(7), 
                           B2 => n96_port, C1 => reg_f(7), C2 => n93_port, ZN 
                           => n53);
   U56 : INV_X1 port map( A => n52, ZN => N87);
   U57 : AOI222_X1 port map( A1 => reg_c(8), A2 => n99_port, B1 => reg_ff(8), 
                           B2 => n96_port, C1 => reg_f(8), C2 => n93_port, ZN 
                           => n52);
   U58 : INV_X1 port map( A => n51, ZN => N88);
   U59 : AOI222_X1 port map( A1 => reg_c(9), A2 => n99_port, B1 => reg_ff(9), 
                           B2 => n95_port, C1 => reg_f(9), C2 => n92_port, ZN 
                           => n51);
   U60 : INV_X1 port map( A => n50, ZN => N89);
   U61 : AOI222_X1 port map( A1 => reg_c(10), A2 => n99_port, B1 => reg_ff(10),
                           B2 => n95_port, C1 => reg_f(10), C2 => n92_port, ZN 
                           => n50);
   U62 : INV_X1 port map( A => n49, ZN => N90);
   U63 : AOI222_X1 port map( A1 => reg_c(11), A2 => n99_port, B1 => reg_ff(11),
                           B2 => n95_port, C1 => reg_f(11), C2 => n92_port, ZN 
                           => n49);
   U64 : INV_X1 port map( A => n48, ZN => N91);
   U65 : AOI222_X1 port map( A1 => reg_c(12), A2 => n99_port, B1 => reg_ff(12),
                           B2 => n95_port, C1 => reg_f(12), C2 => n92_port, ZN 
                           => n48);
   U66 : INV_X1 port map( A => n47, ZN => N92);
   U67 : AOI222_X1 port map( A1 => reg_c(13), A2 => n100_port, B1 => reg_ff(13)
                           , B2 => n95_port, C1 => reg_f(13), C2 => n92_port, 
                           ZN => n47);
   U68 : INV_X1 port map( A => n46, ZN => N93);
   U69 : AOI222_X1 port map( A1 => reg_c(14), A2 => n100_port, B1 => reg_ff(14)
                           , B2 => n95_port, C1 => reg_f(14), C2 => n92_port, 
                           ZN => n46);
   U70 : INV_X1 port map( A => n45, ZN => N94);
   U71 : AOI222_X1 port map( A1 => reg_c(15), A2 => n100_port, B1 => reg_ff(15)
                           , B2 => n95_port, C1 => reg_f(15), C2 => n92_port, 
                           ZN => n45);
   U72 : INV_X1 port map( A => n44, ZN => N95);
   U73 : AOI222_X1 port map( A1 => reg_c(16), A2 => n100_port, B1 => reg_ff(16)
                           , B2 => n95_port, C1 => reg_f(16), C2 => n92_port, 
                           ZN => n44);
   U74 : INV_X1 port map( A => n43, ZN => N96);
   U75 : AOI222_X1 port map( A1 => reg_c(17), A2 => n100_port, B1 => reg_ff(17)
                           , B2 => n95_port, C1 => reg_f(17), C2 => n92_port, 
                           ZN => n43);
   U76 : INV_X1 port map( A => n42, ZN => N97);
   U77 : AOI222_X1 port map( A1 => reg_c(18), A2 => n100_port, B1 => reg_ff(18)
                           , B2 => n95_port, C1 => reg_f(18), C2 => n92_port, 
                           ZN => n42);
   U78 : INV_X1 port map( A => n41, ZN => N98);
   U79 : AOI222_X1 port map( A1 => reg_c(19), A2 => n100_port, B1 => reg_ff(19)
                           , B2 => n95_port, C1 => reg_f(19), C2 => n92_port, 
                           ZN => n41);
   U80 : INV_X1 port map( A => n37, ZN => N99);
   U81 : AOI222_X1 port map( A1 => reg_c(20), A2 => n100_port, B1 => reg_ff(20)
                           , B2 => n96_port, C1 => reg_f(20), C2 => n93_port, 
                           ZN => n37);
   U82 : INV_X1 port map( A => n71, ZN => N100);
   U91 : AOI222_X1 port map( A1 => reg_c(21), A2 => n98_port, B1 => reg_ff(21),
                           B2 => n95_port, C1 => reg_f(21), C2 => n92_port, ZN 
                           => n71);
   U92 : INV_X1 port map( A => n62, ZN => N109);
   U93 : AOI222_X1 port map( A1 => reg_c(30), A2 => n98_port, B1 => reg_ff(30),
                           B2 => n96_port, C1 => reg_f(30), C2 => n93_port, ZN 
                           => n62);
   U94 : INV_X1 port map( A => n61, ZN => N110);
   U95 : AOI222_X1 port map( A1 => reg_c(31), A2 => n98_port, B1 => reg_ff(31),
                           B2 => n96_port, C1 => reg_f(31), C2 => n93_port, ZN 
                           => n61);
   U96 : INV_X1 port map( A => addr_c(3), ZN => n76);
   U97 : AND2_X1 port map( A1 => dirty_f, A2 => n94_port, ZN => N112);
   U98 : AND2_X1 port map( A1 => dirty_ff, A2 => n97_port, ZN => N111);
   U99 : AOI222_X1 port map( A1 => reg_c(0), A2 => n98_port, B1 => reg_ff(0), 
                           B2 => n96_port, C1 => reg_f(0), C2 => n93_port, ZN 
                           => n60);

end SYN_fwd_mux_2_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity RegisterFile_DATA_SIZE32_REG_NUM32 is

   port( clk, rst, en, rd1_en, rd2_en, wr_en, link_en : in std_logic;  rd1_addr
         , rd2_addr, wr_addr : in std_logic_vector (4 downto 0);  d_out1, 
         d_out2 : out std_logic_vector (31 downto 0);  d_in, d_link : in 
         std_logic_vector (31 downto 0));

end RegisterFile_DATA_SIZE32_REG_NUM32;

architecture SYN_register_file_arch of RegisterFile_DATA_SIZE32_REG_NUM32 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal d_out2_31_port, d_out2_30_port, d_out2_29_port, d_out2_28_port, 
      d_out2_27_port, d_out2_26_port, d_out2_25_port, d_out2_24_port, 
      d_out2_23_port, d_out2_22_port, d_out2_21_port, d_out2_20_port, 
      d_out2_19_port, d_out2_18_port, d_out2_17_port, d_out2_16_port, 
      d_out2_15_port, d_out2_14_port, d_out2_13_port, d_out2_12_port, 
      d_out2_11_port, d_out2_10_port, d_out2_9_port, d_out2_8_port, 
      d_out2_7_port, d_out2_6_port, d_out2_5_port, d_out2_4_port, d_out2_3_port
      , d_out2_2_port, d_out2_1_port, d_out2_0_port, registers_2_31_port, 
      registers_2_30_port, registers_2_29_port, registers_2_28_port, 
      registers_2_27_port, registers_2_26_port, registers_2_25_port, 
      registers_2_24_port, registers_2_23_port, registers_2_22_port, 
      registers_2_21_port, registers_2_20_port, registers_2_19_port, 
      registers_2_18_port, registers_2_17_port, registers_2_16_port, 
      registers_2_15_port, registers_2_14_port, registers_2_13_port, 
      registers_2_12_port, registers_2_11_port, registers_2_10_port, 
      registers_2_9_port, registers_2_8_port, registers_2_7_port, 
      registers_2_6_port, registers_2_5_port, registers_2_4_port, 
      registers_2_3_port, registers_2_2_port, registers_2_1_port, 
      registers_2_0_port, registers_3_31_port, registers_3_30_port, 
      registers_3_29_port, registers_3_28_port, registers_3_27_port, 
      registers_3_26_port, registers_3_25_port, registers_3_24_port, 
      registers_3_23_port, registers_3_22_port, registers_3_21_port, 
      registers_3_20_port, registers_3_19_port, registers_3_18_port, 
      registers_3_17_port, registers_3_16_port, registers_3_15_port, 
      registers_3_14_port, registers_3_13_port, registers_3_12_port, 
      registers_3_11_port, registers_3_10_port, registers_3_9_port, 
      registers_3_8_port, registers_3_7_port, registers_3_6_port, 
      registers_3_5_port, registers_3_4_port, registers_3_3_port, 
      registers_3_2_port, registers_3_1_port, registers_3_0_port, 
      registers_5_31_port, registers_5_30_port, registers_5_29_port, 
      registers_5_28_port, registers_5_27_port, registers_5_26_port, 
      registers_5_25_port, registers_5_24_port, registers_5_23_port, 
      registers_5_22_port, registers_5_21_port, registers_5_20_port, 
      registers_5_19_port, registers_5_18_port, registers_5_17_port, 
      registers_5_16_port, registers_5_15_port, registers_5_14_port, 
      registers_5_13_port, registers_5_12_port, registers_5_11_port, 
      registers_5_10_port, registers_5_9_port, registers_5_8_port, 
      registers_5_7_port, registers_5_6_port, registers_5_5_port, 
      registers_5_4_port, registers_5_3_port, registers_5_2_port, 
      registers_5_1_port, registers_5_0_port, registers_7_31_port, 
      registers_7_30_port, registers_7_29_port, registers_7_28_port, 
      registers_7_27_port, registers_7_26_port, registers_7_25_port, 
      registers_7_24_port, registers_7_23_port, registers_7_22_port, 
      registers_7_21_port, registers_7_20_port, registers_7_19_port, 
      registers_7_18_port, registers_7_17_port, registers_7_16_port, 
      registers_7_15_port, registers_7_14_port, registers_7_13_port, 
      registers_7_12_port, registers_7_11_port, registers_7_10_port, 
      registers_7_9_port, registers_7_8_port, registers_7_7_port, 
      registers_7_6_port, registers_7_5_port, registers_7_4_port, 
      registers_7_3_port, registers_7_2_port, registers_7_1_port, 
      registers_7_0_port, registers_8_31_port, registers_8_30_port, 
      registers_8_29_port, registers_8_28_port, registers_8_27_port, 
      registers_8_26_port, registers_8_25_port, registers_8_24_port, 
      registers_8_23_port, registers_8_22_port, registers_8_21_port, 
      registers_8_20_port, registers_8_19_port, registers_8_18_port, 
      registers_8_17_port, registers_8_16_port, registers_8_15_port, 
      registers_8_14_port, registers_8_13_port, registers_8_12_port, 
      registers_8_11_port, registers_8_10_port, registers_8_9_port, 
      registers_8_8_port, registers_8_7_port, registers_8_6_port, 
      registers_8_5_port, registers_8_4_port, registers_8_3_port, 
      registers_8_2_port, registers_8_1_port, registers_8_0_port, 
      registers_9_31_port, registers_9_30_port, registers_9_29_port, 
      registers_9_28_port, registers_9_27_port, registers_9_26_port, 
      registers_9_25_port, registers_9_24_port, registers_9_23_port, 
      registers_9_22_port, registers_9_21_port, registers_9_20_port, 
      registers_9_19_port, registers_9_18_port, registers_9_17_port, 
      registers_9_16_port, registers_9_15_port, registers_9_14_port, 
      registers_9_13_port, registers_9_12_port, registers_9_11_port, 
      registers_9_10_port, registers_9_9_port, registers_9_8_port, 
      registers_9_7_port, registers_9_6_port, registers_9_5_port, 
      registers_9_4_port, registers_9_3_port, registers_9_2_port, 
      registers_9_1_port, registers_9_0_port, registers_11_31_port, 
      registers_11_30_port, registers_11_29_port, registers_11_28_port, 
      registers_11_27_port, registers_11_26_port, registers_11_25_port, 
      registers_11_24_port, registers_11_23_port, registers_11_22_port, 
      registers_11_21_port, registers_11_20_port, registers_11_19_port, 
      registers_11_18_port, registers_11_17_port, registers_11_16_port, 
      registers_11_15_port, registers_11_14_port, registers_11_13_port, 
      registers_11_12_port, registers_11_11_port, registers_11_10_port, 
      registers_11_9_port, registers_11_8_port, registers_11_7_port, 
      registers_11_6_port, registers_11_5_port, registers_11_4_port, 
      registers_11_3_port, registers_11_2_port, registers_11_1_port, 
      registers_11_0_port, registers_12_0_port, registers_13_31_port, 
      registers_13_30_port, registers_13_29_port, registers_13_28_port, 
      registers_13_27_port, registers_13_26_port, registers_13_25_port, 
      registers_13_24_port, registers_13_23_port, registers_13_22_port, 
      registers_13_21_port, registers_13_20_port, registers_13_19_port, 
      registers_13_18_port, registers_13_17_port, registers_13_16_port, 
      registers_13_15_port, registers_13_14_port, registers_13_13_port, 
      registers_13_12_port, registers_13_11_port, registers_13_10_port, 
      registers_13_9_port, registers_13_8_port, registers_13_7_port, 
      registers_13_6_port, registers_13_5_port, registers_13_4_port, 
      registers_13_3_port, registers_13_2_port, registers_13_1_port, 
      registers_13_0_port, registers_14_31_port, registers_14_30_port, 
      registers_14_29_port, registers_14_28_port, registers_14_27_port, 
      registers_14_26_port, registers_14_25_port, registers_14_24_port, 
      registers_14_23_port, registers_14_22_port, registers_14_21_port, 
      registers_14_20_port, registers_14_19_port, registers_14_18_port, 
      registers_14_17_port, registers_14_16_port, registers_14_15_port, 
      registers_14_14_port, registers_14_13_port, registers_14_12_port, 
      registers_14_11_port, registers_14_10_port, registers_14_9_port, 
      registers_14_8_port, registers_14_7_port, registers_14_6_port, 
      registers_14_5_port, registers_14_4_port, registers_14_3_port, 
      registers_14_2_port, registers_14_1_port, registers_14_0_port, 
      registers_15_31_port, registers_15_30_port, registers_15_29_port, 
      registers_15_28_port, registers_15_27_port, registers_15_26_port, 
      registers_15_25_port, registers_15_24_port, registers_15_23_port, 
      registers_15_22_port, registers_15_21_port, registers_15_20_port, 
      registers_15_19_port, registers_15_18_port, registers_15_17_port, 
      registers_15_16_port, registers_15_15_port, registers_15_14_port, 
      registers_15_13_port, registers_15_12_port, registers_15_11_port, 
      registers_15_10_port, registers_15_9_port, registers_15_8_port, 
      registers_15_7_port, registers_15_6_port, registers_15_5_port, 
      registers_15_4_port, registers_15_3_port, registers_15_2_port, 
      registers_15_1_port, registers_15_0_port, registers_16_31_port, 
      registers_16_30_port, registers_16_29_port, registers_16_28_port, 
      registers_16_27_port, registers_16_26_port, registers_16_25_port, 
      registers_16_24_port, registers_16_23_port, registers_16_22_port, 
      registers_16_21_port, registers_16_20_port, registers_16_19_port, 
      registers_16_18_port, registers_16_17_port, registers_16_16_port, 
      registers_16_15_port, registers_16_14_port, registers_16_13_port, 
      registers_16_12_port, registers_16_11_port, registers_16_10_port, 
      registers_16_9_port, registers_16_8_port, registers_16_7_port, 
      registers_16_6_port, registers_16_5_port, registers_16_4_port, 
      registers_16_3_port, registers_16_2_port, registers_16_1_port, 
      registers_16_0_port, registers_17_31_port, registers_17_30_port, 
      registers_17_29_port, registers_17_28_port, registers_17_27_port, 
      registers_17_26_port, registers_17_25_port, registers_17_24_port, 
      registers_17_23_port, registers_17_22_port, registers_17_21_port, 
      registers_17_20_port, registers_17_19_port, registers_17_18_port, 
      registers_17_17_port, registers_17_16_port, registers_17_15_port, 
      registers_17_14_port, registers_17_13_port, registers_17_12_port, 
      registers_17_11_port, registers_17_10_port, registers_17_9_port, 
      registers_17_8_port, registers_17_7_port, registers_17_6_port, 
      registers_17_5_port, registers_17_4_port, registers_17_3_port, 
      registers_17_2_port, registers_17_1_port, registers_17_0_port, 
      registers_19_31_port, registers_19_30_port, registers_19_29_port, 
      registers_19_28_port, registers_19_27_port, registers_19_26_port, 
      registers_19_25_port, registers_19_24_port, registers_19_23_port, 
      registers_19_22_port, registers_19_21_port, registers_19_20_port, 
      registers_19_19_port, registers_19_18_port, registers_19_17_port, 
      registers_19_16_port, registers_19_15_port, registers_19_14_port, 
      registers_19_13_port, registers_19_12_port, registers_19_11_port, 
      registers_19_10_port, registers_19_9_port, registers_19_8_port, 
      registers_19_7_port, registers_19_6_port, registers_19_5_port, 
      registers_19_4_port, registers_19_3_port, registers_19_2_port, 
      registers_19_1_port, registers_19_0_port, registers_20_31_port, 
      registers_20_30_port, registers_20_29_port, registers_20_28_port, 
      registers_20_27_port, registers_20_26_port, registers_20_25_port, 
      registers_20_24_port, registers_20_23_port, registers_20_22_port, 
      registers_20_21_port, registers_20_20_port, registers_20_19_port, 
      registers_20_18_port, registers_20_17_port, registers_20_16_port, 
      registers_20_15_port, registers_20_14_port, registers_20_13_port, 
      registers_20_12_port, registers_20_11_port, registers_20_10_port, 
      registers_20_9_port, registers_20_8_port, registers_20_7_port, 
      registers_20_6_port, registers_20_5_port, registers_20_4_port, 
      registers_20_3_port, registers_20_2_port, registers_20_1_port, 
      registers_21_31_port, registers_21_30_port, registers_21_29_port, 
      registers_21_28_port, registers_21_27_port, registers_21_26_port, 
      registers_21_25_port, registers_21_24_port, registers_21_23_port, 
      registers_21_22_port, registers_21_21_port, registers_21_20_port, 
      registers_21_19_port, registers_21_18_port, registers_21_17_port, 
      registers_21_16_port, registers_21_15_port, registers_21_14_port, 
      registers_21_13_port, registers_21_12_port, registers_21_11_port, 
      registers_21_10_port, registers_21_9_port, registers_21_8_port, 
      registers_21_7_port, registers_21_6_port, registers_21_5_port, 
      registers_21_4_port, registers_21_3_port, registers_21_2_port, 
      registers_21_1_port, registers_21_0_port, registers_22_31_port, 
      registers_22_30_port, registers_22_29_port, registers_22_28_port, 
      registers_22_27_port, registers_22_26_port, registers_22_25_port, 
      registers_22_24_port, registers_22_23_port, registers_22_22_port, 
      registers_22_21_port, registers_22_20_port, registers_22_19_port, 
      registers_22_18_port, registers_22_17_port, registers_22_16_port, 
      registers_22_15_port, registers_22_14_port, registers_22_13_port, 
      registers_22_12_port, registers_22_11_port, registers_22_10_port, 
      registers_22_9_port, registers_22_8_port, registers_22_7_port, 
      registers_22_6_port, registers_22_5_port, registers_22_4_port, 
      registers_22_3_port, registers_22_2_port, registers_22_1_port, 
      registers_22_0_port, registers_25_31_port, registers_25_30_port, 
      registers_25_29_port, registers_25_28_port, registers_25_27_port, 
      registers_25_26_port, registers_25_25_port, registers_25_24_port, 
      registers_25_23_port, registers_25_22_port, registers_25_21_port, 
      registers_25_20_port, registers_25_19_port, registers_25_18_port, 
      registers_25_17_port, registers_25_16_port, registers_25_15_port, 
      registers_25_14_port, registers_25_13_port, registers_25_12_port, 
      registers_25_11_port, registers_25_10_port, registers_25_9_port, 
      registers_25_8_port, registers_25_7_port, registers_25_6_port, 
      registers_25_5_port, registers_25_4_port, registers_25_3_port, 
      registers_25_2_port, registers_25_1_port, registers_25_0_port, 
      registers_26_31_port, registers_26_30_port, registers_26_29_port, 
      registers_26_28_port, registers_26_27_port, registers_26_26_port, 
      registers_26_25_port, registers_26_24_port, registers_26_23_port, 
      registers_26_22_port, registers_26_21_port, registers_26_20_port, 
      registers_26_19_port, registers_26_18_port, registers_26_17_port, 
      registers_26_16_port, registers_26_15_port, registers_26_14_port, 
      registers_26_13_port, registers_26_12_port, registers_26_11_port, 
      registers_26_10_port, registers_26_9_port, registers_26_8_port, 
      registers_26_7_port, registers_26_6_port, registers_26_5_port, 
      registers_26_4_port, registers_26_3_port, registers_26_2_port, 
      registers_26_1_port, registers_26_0_port, registers_27_31_port, 
      registers_27_30_port, registers_27_29_port, registers_27_28_port, 
      registers_27_27_port, registers_27_26_port, registers_27_25_port, 
      registers_27_24_port, registers_27_23_port, registers_27_22_port, 
      registers_27_21_port, registers_27_20_port, registers_27_19_port, 
      registers_27_18_port, registers_27_17_port, registers_27_16_port, 
      registers_27_15_port, registers_27_14_port, registers_27_13_port, 
      registers_27_12_port, registers_27_11_port, registers_27_10_port, 
      registers_27_9_port, registers_27_8_port, registers_27_7_port, 
      registers_27_6_port, registers_27_5_port, registers_27_4_port, 
      registers_27_3_port, registers_27_2_port, registers_27_1_port, 
      registers_28_31_port, registers_28_30_port, registers_28_29_port, 
      registers_28_28_port, registers_28_27_port, registers_28_26_port, 
      registers_28_25_port, registers_28_24_port, registers_28_23_port, 
      registers_28_22_port, registers_28_21_port, registers_28_20_port, 
      registers_28_19_port, registers_28_18_port, registers_28_17_port, 
      registers_28_16_port, registers_28_15_port, registers_28_14_port, 
      registers_28_13_port, registers_28_12_port, registers_28_11_port, 
      registers_28_10_port, registers_28_9_port, registers_28_8_port, 
      registers_28_7_port, registers_28_6_port, registers_28_5_port, 
      registers_28_4_port, registers_28_3_port, registers_28_2_port, 
      registers_28_1_port, registers_28_0_port, registers_29_31_port, 
      registers_29_30_port, registers_29_29_port, registers_29_28_port, 
      registers_29_27_port, registers_29_26_port, registers_29_25_port, 
      registers_29_24_port, registers_29_23_port, registers_29_22_port, 
      registers_29_21_port, registers_29_20_port, registers_29_19_port, 
      registers_29_18_port, registers_29_17_port, registers_29_16_port, 
      registers_29_15_port, registers_29_14_port, registers_29_13_port, 
      registers_29_12_port, registers_29_11_port, registers_29_10_port, 
      registers_29_9_port, registers_29_8_port, registers_29_7_port, 
      registers_29_6_port, registers_29_5_port, registers_29_4_port, 
      registers_29_3_port, registers_29_2_port, registers_29_1_port, 
      registers_29_0_port, registers_30_31_port, registers_30_30_port, 
      registers_30_29_port, registers_30_28_port, registers_30_27_port, 
      registers_30_26_port, registers_30_25_port, registers_30_24_port, 
      registers_30_23_port, registers_30_22_port, registers_30_21_port, 
      registers_30_20_port, registers_30_19_port, registers_30_18_port, 
      registers_30_17_port, registers_30_16_port, registers_30_15_port, 
      registers_30_14_port, registers_30_13_port, registers_30_12_port, 
      registers_30_11_port, registers_30_10_port, registers_30_9_port, 
      registers_30_8_port, registers_30_7_port, registers_30_6_port, 
      registers_30_5_port, registers_30_4_port, registers_30_3_port, 
      registers_30_2_port, registers_30_1_port, registers_30_0_port, 
      registers_31_30_port, registers_31_29_port, registers_31_28_port, 
      registers_31_27_port, registers_31_26_port, registers_31_25_port, 
      registers_31_24_port, registers_31_23_port, registers_31_22_port, 
      registers_31_21_port, registers_31_20_port, registers_31_19_port, 
      registers_31_18_port, registers_31_17_port, registers_31_16_port, 
      registers_31_15_port, registers_31_14_port, registers_31_13_port, 
      registers_31_12_port, registers_31_11_port, registers_31_10_port, 
      registers_31_9_port, registers_31_8_port, registers_31_7_port, 
      registers_31_6_port, registers_31_5_port, registers_31_4_port, 
      registers_31_3_port, registers_31_2_port, registers_31_1_port, 
      registers_31_0_port, n2951, n2952, n2953, n2954, n2955, n2956, n2957, 
      n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, 
      n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, 
      n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, 
      n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, 
      n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, 
      n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, 
      n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, 
      n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, 
      n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, 
      n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, 
      n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, 
      n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, 
      n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, 
      n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, 
      n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, 
      n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, 
      n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, 
      n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, 
      n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, 
      n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, 
      n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, 
      n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, 
      n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, 
      n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, 
      n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, 
      n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, 
      n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, 
      n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, 
      n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, 
      n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, 
      n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, 
      n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, 
      n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, 
      n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, 
      n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, 
      n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, 
      n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, 
      n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, 
      n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, 
      n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, 
      n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, 
      n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, 
      n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, 
      n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, 
      n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, 
      n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, 
      n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, 
      n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, 
      n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, 
      n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, 
      n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, 
      n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, 
      n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, 
      n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, 
      n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, 
      n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, 
      n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, 
      n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, 
      n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, 
      n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, 
      n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, 
      n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, 
      n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, 
      n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, 
      n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, 
      n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, 
      n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, 
      n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, 
      n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, 
      n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, 
      n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, 
      n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, 
      n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, 
      n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, 
      n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, 
      n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, 
      n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, 
      n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, 
      n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, 
      n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, 
      n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, 
      n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, 
      n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, 
      n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, 
      n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, 
      n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, 
      n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, 
      n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, 
      n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, 
      n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, 
      n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, 
      n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, 
      n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, 
      n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, 
      n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, 
      n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, 
      n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, 
      n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, 
      n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, 
      n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, 
      n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, 
      n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, 
      n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, 
      n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, 
      n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n640, 
      net108129, net108130, net108131, net108132, net108133, net108134, 
      net108135, net108136, net108137, net108138, net108139, net108140, 
      net108141, net108142, net108143, net108144, net108145, net108146, 
      net108147, net108148, net108149, net108150, net108151, net108152, 
      net108153, net108154, net108155, net108156, net108157, net108158, 
      net108159, net108160, net108161, net108162, net108355, n1628, n1629, 
      n1632, n1634, n1636, n1638, n1640, n1642, n1644, n1646, n1648, n1650, 
      n1652, n1654, n1656, n1658, n1660, n1662, n1664, n1666, n1668, n1670, 
      n1672, n1674, n1676, n1678, n1680, n1682, n1684, n1686, n1688, n1690, 
      n1692, n1694, n1695, n1696, n1698, n1699, n1700, n1701, n1702, n1703, 
      n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, 
      n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, 
      n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1765, n1766, n1767, 
      n1768, n1769, n1803, n1804, n1805, n1838, n1839, n1873, n1907, n1909, 
      n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, 
      n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, 
      n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, 
      n1940, n1941, n1942, n1976, n2010, n2044, n2078, n2079, n2081, n2082, 
      n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, 
      n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, 
      n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2113, 
      n2147, n2180, n2181, n2182, n2183, n2217, n2218, n2252, n2286, n2320, 
      n2321, n2355, n2356, n2390, n2424, n2458, n2492, n2493, n2527, n2561, 
      n2595, n2629, n2630, n2664, n2665, n2699, n2700, n2702, n2703, n2704, 
      n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, 
      n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, 
      n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, 
      n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, 
      n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, 
      n2755, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, 
      n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2776, 
      n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, 
      n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2795, n2796, n2797, 
      n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, 
      n2808, n2809, n2810, n2811, n2812, n2814, n2815, n2816, n2817, n2818, 
      n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, 
      n2829, n2830, n2831, n2833, n2834, n2835, n2836, n2837, n2838, n2839, 
      n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, 
      n2850, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, 
      n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2871, 
      n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, 
      n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2890, n2891, n2892, 
      n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, 
      n2903, n2904, n2905, n2906, n2907, n2909, n2910, n2911, n2912, n2913, 
      n2914, n2915, n2916, n2917, n2918, n2950, n4007, n4008, n4009, n4010, 
      n4011, n4012, n4013, n4015, n4016, n4017, n4018, n4019, n4020, n4021, 
      n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, 
      n4032, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, 
      n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4053, 
      n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, 
      n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4072, n4073, n4074, 
      n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, 
      n4085, n4086, n4087, n4088, n4089, n4091, n4092, n4093, n4094, n4095, 
      n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, 
      n4106, n4107, n4108, n4110, n4111, n4112, n4113, n4114, n4115, n4116, 
      n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, 
      n4127, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, 
      n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4148, 
      n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, 
      n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4167, n4168, n4169, 
      n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, 
      n4180, n4181, n4182, n4183, n4184, n4186, n4187, n4188, n4189, n4190, 
      n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, 
      n4201, n4202, n4203, n4205, n4206, n4207, n4208, n4209, n4210, n4211, 
      n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, 
      n4222, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, 
      n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4243, 
      n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, 
      n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4262, n4263, n4264, 
      n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, 
      n4275, n4276, n4277, n4278, n4279, n4281, n4282, n4283, n4284, n4285, 
      n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, 
      n4296, n4297, n4298, n4300, n4301, n4302, n4303, n4304, n4305, n4306, 
      n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, 
      n4317, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, 
      n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4338, 
      n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, 
      n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4357, n4358, n4359, 
      n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, 
      n4370, n4371, n4372, n4373, n4374, n4376, n4377, n4378, n4379, n4380, 
      n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, 
      n4391, n4392, n4393, n4395, n4396, n4397, n4398, n4399, n4400, n4401, 
      n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, 
      n4412, n4413, n4414, n4415, n4417, n4418, n4419, n4420, n4421, n4422, 
      n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4432, n4433, 
      n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, 
      n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, 
      n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, 
      n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, 
      n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, 
      n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, 
      n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, 
      n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, 
      n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, 
      n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, 
      n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, 
      n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, 
      n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, 
      n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, 
      n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, 
      n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, 
      n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, 
      n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, 
      n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, 
      n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, 
      n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, 
      n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, 
      n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, 
      n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, 
      n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, 
      n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, 
      n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, 
      n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, 
      n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, 
      n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, 
      n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, 
      n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, 
      n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, 
      n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, 
      n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, 
      n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, 
      n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, 
      n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, 
      n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, 
      n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, 
      n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, 
      n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, 
      n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, 
      n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, 
      n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, 
      n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, 
      n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, 
      n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, 
      n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, 
      n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, 
      n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, 
      n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, 
      n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, 
      n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, 
      n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, 
      n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, 
      n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, 
      n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, 
      n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, 
      n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, 
      n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, 
      n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, 
      n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, 
      n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, 
      n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, 
      n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, 
      n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n2050, 
      n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, 
      n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, 
      n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2080, n2112, n2114, 
      n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, 
      n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, 
      n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, 
      n2145, n2146, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, 
      n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, 
      n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, 
      n2176, n2177, n2178, n2179, n2184, n2185, n2186, n2187, n2188, n2189, 
      n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, 
      n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, 
      n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2219, n2220, n2221, 
      n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, 
      n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, 
      n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, 
      n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, 
      n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, 
      n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, 
      n2283, n2284, n2285, n2287, n2288, n2289, n2290, n2291, n2292, n2293, 
      n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, 
      n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, 
      n2314, n2315, n2316, n2317, n2318, n2319, n2322, n2323, n2324, n2325, 
      n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, 
      n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, 
      n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2357, 
      n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, 
      n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, 
      n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, 
      n2388, n2389, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, 
      n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, 
      n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, 
      n2419, n2420, n2421, n2422, n2423, n2425, n2426, n2427, n2428, n2429, 
      n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, 
      n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, 
      n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2459, n2460, 
      n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, 
      n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, 
      n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, 
      n2491, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, 
      n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, 
      n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, 
      n2523, n2524, n2525, n2526, n2528, n2529, n2530, n2531, n2532, n2533, 
      n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, 
      n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, 
      n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2562, n2563, n2564, 
      n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, 
      n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584, 
      n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594, 
      n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, 
      n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, 
      n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, 
      n2626, n2627, n2628, n2631, n2632, n2633, n2634, n2635, n2636, n2637, 
      n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, 
      n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, 
      n2658, n2659, n2660, n2661, n2662, n2663, n2666, n2667, n2668, n2669, 
      n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, 
      n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, 
      n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2701, 
      n2756, n2775, n2794, n2813, n2832, n2851, n2870, n2889, n2908, n2919, 
      n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, 
      n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, 
      n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, 
      n4014, n4033, n4052, n4071, n4090, n4109, n4128, n4147, n4166, n4185, 
      n4204, n4223, n4242, n4261, n4280, n4299, n4318, n4337, n4356, n4375, 
      n4394, n4416, n4431, n5103, n5104, n5105, n5106, n5107, n5108, n5109, 
      n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, 
      n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, 
      n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, 
      n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, 
      n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, 
      n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, 
      n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, 
      n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, 
      n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, 
      n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, 
      n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, 
      n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, 
      n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, 
      n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, 
      n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, 
      n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, 
      n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, 
      n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, 
      n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, 
      n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, 
      n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, 
      n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, 
      n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, 
      n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, 
      n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, 
      n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, 
      n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, 
      n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, 
      n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, 
      n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, 
      n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, 
      n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, 
      n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, 
      n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, 
      n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, 
      n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, 
      n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, 
      n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, 
      n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, 
      n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, 
      n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, 
      n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, 
      n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, 
      n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, 
      n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, 
      n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, 
      n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, 
      n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, 
      n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, 
      n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, 
      n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, 
      n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, 
      n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, 
      n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, 
      n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, 
      n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, 
      n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, 
      n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, 
      n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, 
      n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, 
      n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, 
      n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, 
      n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, 
      n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, 
      n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, 
      n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, 
      n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, 
      n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, 
      n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, 
      n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, 
      n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, 
      n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, 
      n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, 
      n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, 
      n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, 
      n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, 
      n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, 
      n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, 
      n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, 
      n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, 
      n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, 
      n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, 
      n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, 
      n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, 
      n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, 
      n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, 
      n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, 
      n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, 
      n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, 
      n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, 
      n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, 
      n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, 
      n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, 
      n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, 
      n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, 
      n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, 
      n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, 
      n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, 
      n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, 
      n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, 
      n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, 
      n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, 
      n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, 
      n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, 
      n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, 
      n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, 
      n6170, net163747, net163748, net163749, net163750, net163751, net163752, 
      net163753, net163754, net163755, net163756, net163757, net163758, 
      net163759, net163760, net163761, net163762, net163763, net163764, 
      net163765, net163766, net163767, net163768, net163769, net163770, 
      net163771, net163772, net163773, net163774, net163775, net163776, 
      net163777, net163778, net163779, net163780, net163781, net163782, 
      net163783, net163784, net163785, net163786, net163787, net163788, 
      net163789, net163790, net163791, net163792, net163793, net163794, 
      net163795, net163796, net163797, net163798, net163799, net163800, 
      net163801, net163802, net163803, net163804, net163805, net163806, 
      net163807, net163808, net163809, net163810, net163811, net163812, 
      net163813, net163814, net163815, net163816, net163817, net163818, 
      net163819, net163820, net163821, net163822, net163823, net163824, 
      net163825, net163826, net163827, net163828, net163829, net163830, 
      net163831, net163832, net163833, net163834, net163835, net163836, 
      net163837, net163838, net163839, net163840, net163841, net163842, 
      net163843, net163844, net163845, net163846, net163847, net163848, 
      net163849, net163850, net163851, net163852, net163853, net163854, 
      net163855, net163856, net163857, net163858, net163859, net163860, 
      net163861, net163862, net163863, net163864, net163865, net163866, 
      net163867, net163868, net163869, net163870, net163871, net163872, 
      net163873, net163874, net163875, net163876, net163877, net163878, 
      net163879, net163880, net163881, net163882, net163883, net163884, 
      net163885, net163886, net163887, net163888, net163889, net163890, 
      net163891, net163892, net163893, net163894, net163895, net163896, 
      net163897, net163898, net163899, net163900, net163901, net163902, 
      net163903, net163904, net163905, net163906, net163907, net163908, 
      net163909, net163910, net163911, net163912, net163913, net163914, 
      net163915, net163916, net163917, net163918, net163919, net163920, 
      net163921, net163922, net163923, net163924, net163925, net163926, 
      net163927, net163928, net163929, net163930, net163931, net163932, 
      net163933, net163934, net163935, net163936, net163937, net163938, 
      net163939, net163940, net163941, net163942, net163943, net163944, 
      net163945, net163946, net163947, net163948, net163949, net163950, 
      net163951, net163952, net163953, net163954, net163955, net163956, 
      net163957, net163958, net163959, net163960, net163961, net163962, 
      net163963, net163964, net163965, net163966, net163967, net163968, 
      net163969, net163970, net163971, net163972, net163973, net163974, 
      net163975, net163976, net163977, net163978, net163979, net163980, 
      net163981, net163982, net163983, net163984, net163985, net163986, 
      net163987, net163988, net163989, net163990, net163991, net163992, 
      net163993, net163994, net163995, net163996, net163997, net163998, 
      net163999, net164000, net164001, net164002, net164003, net164004, 
      net164005, net164006, net164007, net164008, net164009, net164010, 
      net164011, net164012, net164013, net164014, net164015, net164016, 
      net164017, net164018, net164019, net164020, net164021, net164022, 
      net164023, net164024, net164025, net164026, net164027, net164028, 
      net164029, net164030, net164031, net164032, net164033, net164034, 
      net164035, net164036, net164037, net164038, net164039, net164040, 
      net164041, net164042, net164043, net164044, net164045, net164046, 
      net164047, net164048, net164049, net164050, net164051, net164052, 
      net164053, net164054, net164055, net164056, net164057, net164058, 
      net164059, net164060, net164061, net164062, net164063, net164064, 
      net164065, net164066, net164067, net164068, net164069, net164070, 
      net164071, net164072, net164073, net164074, net164075, net164076, 
      net164077, net164078, net164079, net164080, net164081, net164082, 
      net164083, net164084, net164085, net164086, net164087, net164088, 
      net164089, net164090, net164091, net164092, net164093, net164094, 
      net164095, net164096, net164097, net164098, net164099, net164100, 
      net164101, net164102, net164103, net164104, net164105, net164106, 
      net164107, net164108, net164109, net164110, net164111, net164112, 
      net164113, net164114, net164115, net164116, net164117, net164118, 
      net164119, net164120, net164121, net164122, net164123, net164124, 
      net164125, net164126, net164127, net164128, net164129, net164130 : 
      std_logic;

begin
   d_out2 <= ( d_out2_31_port, d_out2_30_port, d_out2_29_port, d_out2_28_port, 
      d_out2_27_port, d_out2_26_port, d_out2_25_port, d_out2_24_port, 
      d_out2_23_port, d_out2_22_port, d_out2_21_port, d_out2_20_port, 
      d_out2_19_port, d_out2_18_port, d_out2_17_port, d_out2_16_port, 
      d_out2_15_port, d_out2_14_port, d_out2_13_port, d_out2_12_port, 
      d_out2_11_port, d_out2_10_port, d_out2_9_port, d_out2_8_port, 
      d_out2_7_port, d_out2_6_port, d_out2_5_port, d_out2_4_port, d_out2_3_port
      , d_out2_2_port, d_out2_1_port, d_out2_0_port );
   
   registers_reg_1_31_inst : DFFR_X1 port map( D => n4006, CK => n640, RN => 
                           n6084, Q => net164130, QN => n2115);
   registers_reg_1_30_inst : DFFR_X1 port map( D => n4005, CK => n640, RN => 
                           n6081, Q => net164129, QN => n2114);
   registers_reg_1_29_inst : DFFR_X1 port map( D => n4004, CK => n640, RN => 
                           n6079, Q => net164128, QN => n2112);
   registers_reg_1_28_inst : DFFR_X1 port map( D => n4003, CK => n640, RN => 
                           n6076, Q => net164127, QN => n2080);
   registers_reg_1_27_inst : DFFR_X1 port map( D => n4002, CK => n640, RN => 
                           n6091, Q => net164126, QN => n2077);
   registers_reg_1_26_inst : DFFR_X1 port map( D => n4001, CK => n640, RN => 
                           n6101, Q => net164125, QN => n2076);
   registers_reg_1_25_inst : DFFR_X1 port map( D => n4000, CK => n640, RN => 
                           n6109, Q => net164124, QN => n2075);
   registers_reg_1_24_inst : DFFR_X1 port map( D => n3999, CK => n640, RN => 
                           n6089, Q => net164123, QN => n2074);
   registers_reg_1_23_inst : DFFR_X1 port map( D => n3998, CK => n640, RN => 
                           n6099, Q => net164122, QN => n2073);
   registers_reg_1_22_inst : DFFR_X1 port map( D => n3997, CK => n640, RN => 
                           n6106, Q => net164121, QN => n2072);
   registers_reg_1_21_inst : DFFR_X1 port map( D => n3996, CK => n640, RN => 
                           n6119, Q => net164120, QN => n2071);
   registers_reg_1_20_inst : DFFR_X1 port map( D => n3995, CK => n640, RN => 
                           n6096, Q => net164119, QN => n2070);
   registers_reg_1_19_inst : DFFR_X1 port map( D => n3994, CK => n640, RN => 
                           n6124, Q => net164118, QN => n2069);
   registers_reg_1_18_inst : DFFR_X1 port map( D => n3993, CK => n640, RN => 
                           n6116, Q => net164117, QN => n2068);
   registers_reg_1_17_inst : DFFR_X1 port map( D => n3992, CK => n640, RN => 
                           n6131, Q => net164116, QN => n2067);
   registers_reg_1_16_inst : DFFR_X1 port map( D => n3991, CK => n640, RN => 
                           n6129, Q => net164115, QN => n2066);
   registers_reg_1_15_inst : DFFR_X1 port map( D => n3990, CK => n640, RN => 
                           n6114, Q => net164114, QN => n2065);
   registers_reg_1_14_inst : DFFR_X1 port map( D => n3989, CK => n640, RN => 
                           n6139, Q => net164113, QN => n2064);
   registers_reg_1_13_inst : DFFR_X1 port map( D => n3988, CK => n640, RN => 
                           n6136, Q => net164112, QN => n2063);
   registers_reg_1_12_inst : DFFR_X1 port map( D => n3987, CK => n640, RN => 
                           n6134, Q => net164111, QN => n2062);
   registers_reg_1_11_inst : DFFR_X1 port map( D => n3986, CK => n640, RN => 
                           n6144, Q => net164110, QN => n2061);
   registers_reg_1_10_inst : DFFR_X1 port map( D => n3985, CK => n640, RN => 
                           n6149, Q => net164109, QN => n2060);
   registers_reg_1_9_inst : DFFR_X1 port map( D => n3984, CK => n640, RN => 
                           n6086, Q => net164108, QN => n2059);
   registers_reg_1_8_inst : DFFR_X1 port map( D => n3983, CK => n640, RN => 
                           n6111, Q => net164107, QN => n2058);
   registers_reg_1_7_inst : DFFR_X1 port map( D => n3982, CK => n640, RN => 
                           n6104, Q => net164106, QN => n2057);
   registers_reg_1_6_inst : DFFR_X1 port map( D => n3981, CK => n640, RN => 
                           n6141, Q => net164105, QN => n2056);
   registers_reg_1_5_inst : DFFR_X1 port map( D => n3980, CK => n640, RN => 
                           n6094, Q => net164104, QN => n2055);
   registers_reg_1_4_inst : DFFR_X1 port map( D => n3979, CK => n640, RN => 
                           n6121, Q => net164103, QN => n2054);
   registers_reg_1_3_inst : DFFR_X1 port map( D => n3978, CK => n640, RN => 
                           n6146, Q => net164102, QN => n2053);
   registers_reg_1_2_inst : DFFR_X1 port map( D => n3977, CK => n640, RN => 
                           n6151, Q => net164101, QN => n2052);
   registers_reg_1_1_inst : DFFR_X1 port map( D => n3976, CK => n640, RN => 
                           n6126, Q => net164100, QN => n2051);
   registers_reg_1_0_inst : DFFR_X1 port map( D => n3975, CK => n640, RN => 
                           n6074, Q => net164099, QN => n2153);
   registers_reg_2_31_inst : DFFR_X1 port map( D => n3974, CK => n640, RN => 
                           n6084, Q => registers_2_31_port, QN => net164098);
   registers_reg_2_30_inst : DFFR_X1 port map( D => n3973, CK => n640, RN => 
                           n6081, Q => registers_2_30_port, QN => net164097);
   registers_reg_2_29_inst : DFFR_X1 port map( D => n3972, CK => n640, RN => 
                           n6079, Q => registers_2_29_port, QN => net164096);
   registers_reg_2_28_inst : DFFR_X1 port map( D => n3971, CK => n640, RN => 
                           n6076, Q => registers_2_28_port, QN => net164095);
   registers_reg_2_27_inst : DFFR_X1 port map( D => n3970, CK => n640, RN => 
                           n6091, Q => registers_2_27_port, QN => net164094);
   registers_reg_2_26_inst : DFFR_X1 port map( D => n3969, CK => n640, RN => 
                           n6101, Q => registers_2_26_port, QN => net164093);
   registers_reg_2_25_inst : DFFR_X1 port map( D => n3968, CK => n640, RN => 
                           n6109, Q => registers_2_25_port, QN => net164092);
   registers_reg_2_24_inst : DFFR_X1 port map( D => n3967, CK => n640, RN => 
                           n6089, Q => registers_2_24_port, QN => net164091);
   registers_reg_2_23_inst : DFFR_X1 port map( D => n3966, CK => n640, RN => 
                           n6099, Q => registers_2_23_port, QN => net164090);
   registers_reg_2_22_inst : DFFR_X1 port map( D => n3965, CK => n640, RN => 
                           n6106, Q => registers_2_22_port, QN => net164089);
   registers_reg_2_21_inst : DFFR_X1 port map( D => n3964, CK => n640, RN => 
                           n6119, Q => registers_2_21_port, QN => net164088);
   registers_reg_2_20_inst : DFFR_X1 port map( D => n3963, CK => n640, RN => 
                           n6096, Q => registers_2_20_port, QN => net164087);
   registers_reg_2_19_inst : DFFR_X1 port map( D => n3962, CK => n640, RN => 
                           n6124, Q => registers_2_19_port, QN => net164086);
   registers_reg_2_18_inst : DFFR_X1 port map( D => n3961, CK => n640, RN => 
                           n6116, Q => registers_2_18_port, QN => net164085);
   registers_reg_2_17_inst : DFFR_X1 port map( D => n3960, CK => n640, RN => 
                           n6131, Q => registers_2_17_port, QN => net164084);
   registers_reg_2_16_inst : DFFR_X1 port map( D => n3959, CK => n640, RN => 
                           n6129, Q => registers_2_16_port, QN => net164083);
   registers_reg_2_15_inst : DFFR_X1 port map( D => n3958, CK => n640, RN => 
                           n6114, Q => registers_2_15_port, QN => net164082);
   registers_reg_2_14_inst : DFFR_X1 port map( D => n3957, CK => n640, RN => 
                           n6139, Q => registers_2_14_port, QN => net164081);
   registers_reg_2_13_inst : DFFR_X1 port map( D => n3956, CK => n640, RN => 
                           n6136, Q => registers_2_13_port, QN => net164080);
   registers_reg_2_12_inst : DFFR_X1 port map( D => n3955, CK => n640, RN => 
                           n6134, Q => registers_2_12_port, QN => net164079);
   registers_reg_2_11_inst : DFFR_X1 port map( D => n3954, CK => n640, RN => 
                           n6144, Q => registers_2_11_port, QN => net164078);
   registers_reg_2_10_inst : DFFR_X1 port map( D => n3953, CK => n640, RN => 
                           n6149, Q => registers_2_10_port, QN => net164077);
   registers_reg_2_9_inst : DFFR_X1 port map( D => n3952, CK => n640, RN => 
                           n6086, Q => registers_2_9_port, QN => net164076);
   registers_reg_2_8_inst : DFFR_X1 port map( D => n3951, CK => n640, RN => 
                           n6111, Q => registers_2_8_port, QN => net164075);
   registers_reg_2_7_inst : DFFR_X1 port map( D => n3950, CK => n640, RN => 
                           n6104, Q => registers_2_7_port, QN => net164074);
   registers_reg_2_6_inst : DFFR_X1 port map( D => n3949, CK => n640, RN => 
                           n6141, Q => registers_2_6_port, QN => net164073);
   registers_reg_2_5_inst : DFFR_X1 port map( D => n3948, CK => n640, RN => 
                           n6094, Q => registers_2_5_port, QN => net164072);
   registers_reg_2_4_inst : DFFR_X1 port map( D => n3947, CK => n640, RN => 
                           n6121, Q => registers_2_4_port, QN => net164071);
   registers_reg_2_3_inst : DFFR_X1 port map( D => n3946, CK => n640, RN => 
                           n6146, Q => registers_2_3_port, QN => net164070);
   registers_reg_2_2_inst : DFFR_X1 port map( D => n3945, CK => n640, RN => 
                           n6151, Q => registers_2_2_port, QN => net164069);
   registers_reg_2_1_inst : DFFR_X1 port map( D => n3944, CK => n640, RN => 
                           n6126, Q => registers_2_1_port, QN => net164068);
   registers_reg_2_0_inst : DFFR_X1 port map( D => n3943, CK => n640, RN => 
                           n6074, Q => registers_2_0_port, QN => net164067);
   registers_reg_3_31_inst : DFFR_X1 port map( D => n3942, CK => n640, RN => 
                           n6084, Q => registers_3_31_port, QN => n5183);
   registers_reg_3_30_inst : DFFR_X1 port map( D => n3941, CK => n640, RN => 
                           n6081, Q => registers_3_30_port, QN => n5182);
   registers_reg_3_29_inst : DFFR_X1 port map( D => n3940, CK => n640, RN => 
                           n6079, Q => registers_3_29_port, QN => n5181);
   registers_reg_3_28_inst : DFFR_X1 port map( D => n3939, CK => n640, RN => 
                           n6076, Q => registers_3_28_port, QN => n5180);
   registers_reg_3_27_inst : DFFR_X1 port map( D => n3938, CK => n640, RN => 
                           n6091, Q => registers_3_27_port, QN => n2388);
   registers_reg_3_26_inst : DFFR_X1 port map( D => n3937, CK => n640, RN => 
                           n6101, Q => registers_3_26_port, QN => n5179);
   registers_reg_3_25_inst : DFFR_X1 port map( D => n3936, CK => n640, RN => 
                           n6109, Q => registers_3_25_port, QN => n5178);
   registers_reg_3_24_inst : DFFR_X1 port map( D => n3935, CK => n640, RN => 
                           n6089, Q => registers_3_24_port, QN => n5177);
   registers_reg_3_23_inst : DFFR_X1 port map( D => n3934, CK => n640, RN => 
                           n6099, Q => registers_3_23_port, QN => n5176);
   registers_reg_3_22_inst : DFFR_X1 port map( D => n3933, CK => n640, RN => 
                           n6106, Q => registers_3_22_port, QN => n5175);
   registers_reg_3_21_inst : DFFR_X1 port map( D => n3932, CK => n640, RN => 
                           n6119, Q => registers_3_21_port, QN => n5174);
   registers_reg_3_20_inst : DFFR_X1 port map( D => n3931, CK => n640, RN => 
                           n6096, Q => registers_3_20_port, QN => n5173);
   registers_reg_3_19_inst : DFFR_X1 port map( D => n3930, CK => n640, RN => 
                           n6124, Q => registers_3_19_port, QN => n5172);
   registers_reg_3_18_inst : DFFR_X1 port map( D => n3929, CK => n640, RN => 
                           n6116, Q => registers_3_18_port, QN => n5171);
   registers_reg_3_17_inst : DFFR_X1 port map( D => n3928, CK => n640, RN => 
                           n6131, Q => registers_3_17_port, QN => n5170);
   registers_reg_3_16_inst : DFFR_X1 port map( D => n3927, CK => n640, RN => 
                           n6129, Q => registers_3_16_port, QN => n5169);
   registers_reg_3_15_inst : DFFR_X1 port map( D => n3926, CK => n640, RN => 
                           n6114, Q => registers_3_15_port, QN => n5168);
   registers_reg_3_14_inst : DFFR_X1 port map( D => n3925, CK => n640, RN => 
                           n6139, Q => registers_3_14_port, QN => n5167);
   registers_reg_3_13_inst : DFFR_X1 port map( D => n3924, CK => n640, RN => 
                           n6136, Q => registers_3_13_port, QN => n5166);
   registers_reg_3_12_inst : DFFR_X1 port map( D => n3923, CK => n640, RN => 
                           n6134, Q => registers_3_12_port, QN => n5165);
   registers_reg_3_11_inst : DFFR_X1 port map( D => n3922, CK => n640, RN => 
                           n6144, Q => registers_3_11_port, QN => n5164);
   registers_reg_3_10_inst : DFFR_X1 port map( D => n3921, CK => n640, RN => 
                           n6149, Q => registers_3_10_port, QN => n5163);
   registers_reg_3_9_inst : DFFR_X1 port map( D => n3920, CK => n640, RN => 
                           n6086, Q => registers_3_9_port, QN => n5162);
   registers_reg_3_8_inst : DFFR_X1 port map( D => n3919, CK => n640, RN => 
                           n6111, Q => registers_3_8_port, QN => n5161);
   registers_reg_3_7_inst : DFFR_X1 port map( D => n3918, CK => n640, RN => 
                           n6104, Q => registers_3_7_port, QN => n5160);
   registers_reg_3_6_inst : DFFR_X1 port map( D => n3917, CK => n640, RN => 
                           n6141, Q => registers_3_6_port, QN => n5159);
   registers_reg_3_5_inst : DFFR_X1 port map( D => n3916, CK => n640, RN => 
                           n6094, Q => registers_3_5_port, QN => n5158);
   registers_reg_3_4_inst : DFFR_X1 port map( D => n3915, CK => n640, RN => 
                           n6121, Q => registers_3_4_port, QN => n5157);
   registers_reg_3_3_inst : DFFR_X1 port map( D => n3914, CK => n640, RN => 
                           n6146, Q => registers_3_3_port, QN => n5156);
   registers_reg_3_2_inst : DFFR_X1 port map( D => n3913, CK => n640, RN => 
                           n6151, Q => registers_3_2_port, QN => n5155);
   registers_reg_3_1_inst : DFFR_X1 port map( D => n3912, CK => n640, RN => 
                           n6126, Q => registers_3_1_port, QN => n5154);
   registers_reg_3_0_inst : DFFR_X1 port map( D => n3911, CK => n640, RN => 
                           n6074, Q => registers_3_0_port, QN => n5123);
   registers_reg_4_31_inst : DFFR_X1 port map( D => n3910, CK => n640, RN => 
                           n6084, Q => net164066, QN => n2139);
   registers_reg_4_30_inst : DFFR_X1 port map( D => n3909, CK => n640, RN => 
                           n6081, Q => net164065, QN => n2138);
   registers_reg_4_29_inst : DFFR_X1 port map( D => n3908, CK => n640, RN => 
                           n6079, Q => net164064, QN => n2152);
   registers_reg_4_28_inst : DFFR_X1 port map( D => n3907, CK => n640, RN => 
                           n6076, Q => net164063, QN => n2149);
   registers_reg_4_27_inst : DFFR_X1 port map( D => n3906, CK => n640, RN => 
                           n6091, Q => net164062, QN => n2148);
   registers_reg_4_26_inst : DFFR_X1 port map( D => n3905, CK => n640, RN => 
                           n6101, Q => net164061, QN => n2151);
   registers_reg_4_25_inst : DFFR_X1 port map( D => n3904, CK => n640, RN => 
                           n6109, Q => net164060, QN => n2146);
   registers_reg_4_24_inst : DFFR_X1 port map( D => n3903, CK => n640, RN => 
                           n6089, Q => net164059, QN => n2145);
   registers_reg_4_23_inst : DFFR_X1 port map( D => n3902, CK => n640, RN => 
                           n6099, Q => net164058, QN => n2144);
   registers_reg_4_22_inst : DFFR_X1 port map( D => n3901, CK => n640, RN => 
                           n6106, Q => net164057, QN => n2143);
   registers_reg_4_21_inst : DFFR_X1 port map( D => n3900, CK => n640, RN => 
                           n6119, Q => net164056, QN => n2142);
   registers_reg_4_20_inst : DFFR_X1 port map( D => n3899, CK => n640, RN => 
                           n6096, Q => net164055, QN => n2141);
   registers_reg_4_19_inst : DFFR_X1 port map( D => n3898, CK => n640, RN => 
                           n6124, Q => net164054, QN => n2137);
   registers_reg_4_18_inst : DFFR_X1 port map( D => n3897, CK => n640, RN => 
                           n6116, Q => net164053, QN => n2136);
   registers_reg_4_17_inst : DFFR_X1 port map( D => n3896, CK => n640, RN => 
                           n6132, Q => net164052, QN => n2150);
   registers_reg_4_16_inst : DFFR_X1 port map( D => n3895, CK => n640, RN => 
                           n6129, Q => net164051, QN => n2135);
   registers_reg_4_15_inst : DFFR_X1 port map( D => n3894, CK => n640, RN => 
                           n6114, Q => net164050, QN => n2134);
   registers_reg_4_14_inst : DFFR_X1 port map( D => n3893, CK => n640, RN => 
                           n6139, Q => net164049, QN => n2133);
   registers_reg_4_13_inst : DFFR_X1 port map( D => n3892, CK => n640, RN => 
                           n6137, Q => net164048, QN => n2132);
   registers_reg_4_12_inst : DFFR_X1 port map( D => n3891, CK => n640, RN => 
                           n6134, Q => net164047, QN => n2131);
   registers_reg_4_11_inst : DFFR_X1 port map( D => n3890, CK => n640, RN => 
                           n6144, Q => net164046, QN => n2130);
   registers_reg_4_10_inst : DFFR_X1 port map( D => n3889, CK => n640, RN => 
                           n6149, Q => net164045, QN => n2129);
   registers_reg_4_9_inst : DFFR_X1 port map( D => n3888, CK => n640, RN => 
                           n6086, Q => net164044, QN => n2128);
   registers_reg_4_8_inst : DFFR_X1 port map( D => n3887, CK => n640, RN => 
                           n6111, Q => net164043, QN => n2140);
   registers_reg_4_7_inst : DFFR_X1 port map( D => n3886, CK => n640, RN => 
                           n6104, Q => net164042, QN => n2127);
   registers_reg_4_6_inst : DFFR_X1 port map( D => n3885, CK => n640, RN => 
                           n6142, Q => net164041, QN => n2126);
   registers_reg_4_5_inst : DFFR_X1 port map( D => n3884, CK => n640, RN => 
                           n6094, Q => net164040, QN => n2125);
   registers_reg_4_4_inst : DFFR_X1 port map( D => n3883, CK => n640, RN => 
                           n6121, Q => net164039, QN => n2124);
   registers_reg_4_3_inst : DFFR_X1 port map( D => n3882, CK => n640, RN => 
                           n6147, Q => net164038, QN => n2123);
   registers_reg_4_2_inst : DFFR_X1 port map( D => n3881, CK => n640, RN => 
                           n6152, Q => net164037, QN => n2122);
   registers_reg_4_1_inst : DFFR_X1 port map( D => n3880, CK => n640, RN => 
                           n6126, Q => net164036, QN => n2121);
   registers_reg_4_0_inst : DFFR_X1 port map( D => n3879, CK => n640, RN => 
                           n6074, Q => net164035, QN => n2511);
   registers_reg_5_31_inst : DFFR_X1 port map( D => n3878, CK => n640, RN => 
                           n6084, Q => registers_5_31_port, QN => n2546);
   registers_reg_5_30_inst : DFFR_X1 port map( D => n3877, CK => n640, RN => 
                           n6082, Q => registers_5_30_port, QN => n2545);
   registers_reg_5_29_inst : DFFR_X1 port map( D => n3876, CK => n640, RN => 
                           n6079, Q => registers_5_29_port, QN => n2554);
   registers_reg_5_28_inst : DFFR_X1 port map( D => n3875, CK => n640, RN => 
                           n6077, Q => registers_5_28_port, QN => n2553);
   registers_reg_5_27_inst : DFFR_X1 port map( D => n3874, CK => n640, RN => 
                           n6092, Q => registers_5_27_port, QN => n2552);
   registers_reg_5_26_inst : DFFR_X1 port map( D => n3873, CK => n640, RN => 
                           n6102, Q => registers_5_26_port, QN => n2551);
   registers_reg_5_25_inst : DFFR_X1 port map( D => n3872, CK => n640, RN => 
                           n6109, Q => registers_5_25_port, QN => n2550);
   registers_reg_5_24_inst : DFFR_X1 port map( D => n3871, CK => n640, RN => 
                           n6089, Q => registers_5_24_port, QN => n2549);
   registers_reg_5_23_inst : DFFR_X1 port map( D => n3870, CK => n640, RN => 
                           n6099, Q => registers_5_23_port, QN => n2548);
   registers_reg_5_22_inst : DFFR_X1 port map( D => n3869, CK => n640, RN => 
                           n6107, Q => registers_5_22_port, QN => n2547);
   registers_reg_5_21_inst : DFFR_X1 port map( D => n3868, CK => n640, RN => 
                           n6119, Q => registers_5_21_port, QN => n2544);
   registers_reg_5_20_inst : DFFR_X1 port map( D => n3867, CK => n640, RN => 
                           n6097, Q => registers_5_20_port, QN => n2543);
   registers_reg_5_19_inst : DFFR_X1 port map( D => n3866, CK => n640, RN => 
                           n6124, Q => registers_5_19_port, QN => n2542);
   registers_reg_5_18_inst : DFFR_X1 port map( D => n3865, CK => n640, RN => 
                           n6117, Q => registers_5_18_port, QN => n2541);
   registers_reg_5_17_inst : DFFR_X1 port map( D => n3864, CK => n640, RN => 
                           n6132, Q => registers_5_17_port, QN => n2540);
   registers_reg_5_16_inst : DFFR_X1 port map( D => n3863, CK => n640, RN => 
                           n6129, Q => registers_5_16_port, QN => n2539);
   registers_reg_5_15_inst : DFFR_X1 port map( D => n3862, CK => n640, RN => 
                           n6114, Q => registers_5_15_port, QN => n2538);
   registers_reg_5_14_inst : DFFR_X1 port map( D => n3861, CK => n640, RN => 
                           n6139, Q => registers_5_14_port, QN => n2537);
   registers_reg_5_13_inst : DFFR_X1 port map( D => n3860, CK => n640, RN => 
                           n6137, Q => registers_5_13_port, QN => n2536);
   registers_reg_5_12_inst : DFFR_X1 port map( D => n3859, CK => n640, RN => 
                           n6134, Q => registers_5_12_port, QN => n2535);
   registers_reg_5_11_inst : DFFR_X1 port map( D => n3858, CK => n640, RN => 
                           n6144, Q => registers_5_11_port, QN => n2534);
   registers_reg_5_10_inst : DFFR_X1 port map( D => n3857, CK => n640, RN => 
                           n6149, Q => registers_5_10_port, QN => n2533);
   registers_reg_5_9_inst : DFFR_X1 port map( D => n3856, CK => n640, RN => 
                           n6087, Q => registers_5_9_port, QN => n2532);
   registers_reg_5_8_inst : DFFR_X1 port map( D => n3855, CK => n640, RN => 
                           n6112, Q => registers_5_8_port, QN => n2531);
   registers_reg_5_7_inst : DFFR_X1 port map( D => n3854, CK => n640, RN => 
                           n6104, Q => registers_5_7_port, QN => n2530);
   registers_reg_5_6_inst : DFFR_X1 port map( D => n3853, CK => n640, RN => 
                           n6142, Q => registers_5_6_port, QN => n2529);
   registers_reg_5_5_inst : DFFR_X1 port map( D => n3852, CK => n640, RN => 
                           n6094, Q => registers_5_5_port, QN => n2528);
   registers_reg_5_4_inst : DFFR_X1 port map( D => n3851, CK => n640, RN => 
                           n6122, Q => registers_5_4_port, QN => n2526);
   registers_reg_5_3_inst : DFFR_X1 port map( D => n3850, CK => n640, RN => 
                           n6147, Q => registers_5_3_port, QN => n2525);
   registers_reg_5_2_inst : DFFR_X1 port map( D => n3849, CK => n640, RN => 
                           n6152, Q => registers_5_2_port, QN => n2524);
   registers_reg_5_1_inst : DFFR_X1 port map( D => n3848, CK => n640, RN => 
                           n6127, Q => registers_5_1_port, QN => n2523);
   registers_reg_5_0_inst : DFFR_X1 port map( D => n3847, CK => n640, RN => 
                           n6074, Q => registers_5_0_port, QN => net164034);
   registers_reg_6_31_inst : DFFR_X1 port map( D => n3846, CK => n640, RN => 
                           n6084, Q => net164033, QN => n2287);
   registers_reg_6_30_inst : DFFR_X1 port map( D => n3845, CK => n640, RN => 
                           n6082, Q => net164032, QN => n2285);
   registers_reg_6_29_inst : DFFR_X1 port map( D => n3844, CK => n640, RN => 
                           n6079, Q => net164031, QN => n2284);
   registers_reg_6_28_inst : DFFR_X1 port map( D => n3843, CK => n640, RN => 
                           n6077, Q => net164030, QN => n2283);
   registers_reg_6_27_inst : DFFR_X1 port map( D => n3842, CK => n640, RN => 
                           n6092, Q => net164029, QN => n2120);
   registers_reg_6_26_inst : DFFR_X1 port map( D => n3841, CK => n640, RN => 
                           n6102, Q => net164028, QN => n2119);
   registers_reg_6_25_inst : DFFR_X1 port map( D => n3840, CK => n640, RN => 
                           n6109, Q => net164027, QN => n2282);
   registers_reg_6_24_inst : DFFR_X1 port map( D => n3839, CK => n640, RN => 
                           n6089, Q => net164026, QN => n2281);
   registers_reg_6_23_inst : DFFR_X1 port map( D => n3838, CK => n640, RN => 
                           n6099, Q => net164025, QN => n2280);
   registers_reg_6_22_inst : DFFR_X1 port map( D => n3837, CK => n640, RN => 
                           n6107, Q => net164024, QN => n2279);
   registers_reg_6_21_inst : DFFR_X1 port map( D => n3836, CK => n640, RN => 
                           n6119, Q => net164023, QN => n2278);
   registers_reg_6_20_inst : DFFR_X1 port map( D => n3835, CK => n640, RN => 
                           n6097, Q => net164022, QN => n2277);
   registers_reg_6_19_inst : DFFR_X1 port map( D => n3834, CK => n640, RN => 
                           n6124, Q => net164021, QN => n2276);
   registers_reg_6_18_inst : DFFR_X1 port map( D => n3833, CK => n640, RN => 
                           n6117, Q => net164020, QN => n2275);
   registers_reg_6_17_inst : DFFR_X1 port map( D => n3832, CK => n640, RN => 
                           n6132, Q => net164019, QN => n2274);
   registers_reg_6_16_inst : DFFR_X1 port map( D => n3831, CK => n640, RN => 
                           n6129, Q => net164018, QN => n2273);
   registers_reg_6_15_inst : DFFR_X1 port map( D => n3830, CK => n640, RN => 
                           n6114, Q => net164017, QN => n2272);
   registers_reg_6_14_inst : DFFR_X1 port map( D => n3829, CK => n640, RN => 
                           n6139, Q => net164016, QN => n2271);
   registers_reg_6_13_inst : DFFR_X1 port map( D => n3828, CK => n640, RN => 
                           n6137, Q => net164015, QN => n2270);
   registers_reg_6_12_inst : DFFR_X1 port map( D => n3827, CK => n640, RN => 
                           n6134, Q => net164014, QN => n2269);
   registers_reg_6_11_inst : DFFR_X1 port map( D => n3826, CK => n640, RN => 
                           n6144, Q => net164013, QN => n2268);
   registers_reg_6_10_inst : DFFR_X1 port map( D => n3825, CK => n640, RN => 
                           n6149, Q => net164012, QN => n2267);
   registers_reg_6_9_inst : DFFR_X1 port map( D => n3824, CK => n640, RN => 
                           n6087, Q => net164011, QN => n2266);
   registers_reg_6_8_inst : DFFR_X1 port map( D => n3823, CK => n640, RN => 
                           n6112, Q => net164010, QN => n2265);
   registers_reg_6_7_inst : DFFR_X1 port map( D => n3822, CK => n640, RN => 
                           n6104, Q => net164009, QN => n2264);
   registers_reg_6_6_inst : DFFR_X1 port map( D => n3821, CK => n640, RN => 
                           n6142, Q => net164008, QN => n2263);
   registers_reg_6_5_inst : DFFR_X1 port map( D => n3820, CK => n640, RN => 
                           n6094, Q => net164007, QN => n2262);
   registers_reg_6_4_inst : DFFR_X1 port map( D => n3819, CK => n640, RN => 
                           n6122, Q => net164006, QN => n2261);
   registers_reg_6_3_inst : DFFR_X1 port map( D => n3818, CK => n640, RN => 
                           n6147, Q => net164005, QN => n2260);
   registers_reg_6_2_inst : DFFR_X1 port map( D => n3817, CK => n640, RN => 
                           n6152, Q => net164004, QN => n2259);
   registers_reg_6_1_inst : DFFR_X1 port map( D => n3816, CK => n640, RN => 
                           n6127, Q => net164003, QN => n2258);
   registers_reg_6_0_inst : DFFR_X1 port map( D => n3815, CK => n640, RN => 
                           n6074, Q => net164002, QN => n2227);
   registers_reg_7_31_inst : DFFR_X1 port map( D => n3814, CK => n640, RN => 
                           n6084, Q => registers_7_31_port, QN => n5144);
   registers_reg_7_30_inst : DFFR_X1 port map( D => n3813, CK => n640, RN => 
                           n6082, Q => registers_7_30_port, QN => n5143);
   registers_reg_7_29_inst : DFFR_X1 port map( D => n3812, CK => n640, RN => 
                           n6079, Q => registers_7_29_port, QN => n5153);
   registers_reg_7_28_inst : DFFR_X1 port map( D => n3811, CK => n640, RN => 
                           n6077, Q => registers_7_28_port, QN => n5142);
   registers_reg_7_27_inst : DFFR_X1 port map( D => n3810, CK => n640, RN => 
                           n6092, Q => registers_7_27_port, QN => n5141);
   registers_reg_7_26_inst : DFFR_X1 port map( D => n3809, CK => n640, RN => 
                           n6102, Q => registers_7_26_port, QN => n2386);
   registers_reg_7_25_inst : DFFR_X1 port map( D => n3808, CK => n640, RN => 
                           n6109, Q => registers_7_25_port, QN => n5140);
   registers_reg_7_24_inst : DFFR_X1 port map( D => n3807, CK => n640, RN => 
                           n6089, Q => registers_7_24_port, QN => n5139);
   registers_reg_7_23_inst : DFFR_X1 port map( D => n3806, CK => n640, RN => 
                           n6099, Q => registers_7_23_port, QN => n5152);
   registers_reg_7_22_inst : DFFR_X1 port map( D => n3805, CK => n640, RN => 
                           n6107, Q => registers_7_22_port, QN => n5138);
   registers_reg_7_21_inst : DFFR_X1 port map( D => n3804, CK => n640, RN => 
                           n6119, Q => registers_7_21_port, QN => n5137);
   registers_reg_7_20_inst : DFFR_X1 port map( D => n3803, CK => n640, RN => 
                           n6097, Q => registers_7_20_port, QN => n5151);
   registers_reg_7_19_inst : DFFR_X1 port map( D => n3802, CK => n640, RN => 
                           n6124, Q => registers_7_19_port, QN => n5136);
   registers_reg_7_18_inst : DFFR_X1 port map( D => n3801, CK => n640, RN => 
                           n6117, Q => registers_7_18_port, QN => n5135);
   registers_reg_7_17_inst : DFFR_X1 port map( D => n3800, CK => n640, RN => 
                           n6132, Q => registers_7_17_port, QN => n5150);
   registers_reg_7_16_inst : DFFR_X1 port map( D => n3799, CK => n640, RN => 
                           n6129, Q => registers_7_16_port, QN => n5134);
   registers_reg_7_15_inst : DFFR_X1 port map( D => n3798, CK => n640, RN => 
                           n6114, Q => registers_7_15_port, QN => n5133);
   registers_reg_7_14_inst : DFFR_X1 port map( D => n3797, CK => n640, RN => 
                           n6139, Q => registers_7_14_port, QN => n5149);
   registers_reg_7_13_inst : DFFR_X1 port map( D => n3796, CK => n640, RN => 
                           n6137, Q => registers_7_13_port, QN => n5132);
   registers_reg_7_12_inst : DFFR_X1 port map( D => n3795, CK => n640, RN => 
                           n6134, Q => registers_7_12_port, QN => n5131);
   registers_reg_7_11_inst : DFFR_X1 port map( D => n3794, CK => n640, RN => 
                           n6144, Q => registers_7_11_port, QN => n5148);
   registers_reg_7_10_inst : DFFR_X1 port map( D => n3793, CK => n640, RN => 
                           n6149, Q => registers_7_10_port, QN => n5130);
   registers_reg_7_9_inst : DFFR_X1 port map( D => n3792, CK => n640, RN => 
                           n6087, Q => registers_7_9_port, QN => n5129);
   registers_reg_7_8_inst : DFFR_X1 port map( D => n3791, CK => n640, RN => 
                           n6112, Q => registers_7_8_port, QN => n5147);
   registers_reg_7_7_inst : DFFR_X1 port map( D => n3790, CK => n640, RN => 
                           n6104, Q => registers_7_7_port, QN => n5128);
   registers_reg_7_6_inst : DFFR_X1 port map( D => n3789, CK => n640, RN => 
                           n6142, Q => registers_7_6_port, QN => n5127);
   registers_reg_7_5_inst : DFFR_X1 port map( D => n3788, CK => n640, RN => 
                           n6094, Q => registers_7_5_port, QN => n5146);
   registers_reg_7_4_inst : DFFR_X1 port map( D => n3787, CK => n640, RN => 
                           n6122, Q => registers_7_4_port, QN => n5126);
   registers_reg_7_3_inst : DFFR_X1 port map( D => n3786, CK => n640, RN => 
                           n6147, Q => registers_7_3_port, QN => n5125);
   registers_reg_7_2_inst : DFFR_X1 port map( D => n3785, CK => n640, RN => 
                           n6152, Q => registers_7_2_port, QN => n5145);
   registers_reg_7_1_inst : DFFR_X1 port map( D => n3784, CK => n640, RN => 
                           n6127, Q => registers_7_1_port, QN => n5124);
   registers_reg_7_0_inst : DFFR_X1 port map( D => n3783, CK => n640, RN => 
                           n6074, Q => registers_7_0_port, QN => n5122);
   registers_reg_8_31_inst : DFFR_X1 port map( D => n3782, CK => n640, RN => 
                           n6084, Q => registers_8_31_port, QN => net164001);
   registers_reg_8_30_inst : DFFR_X1 port map( D => n3781, CK => n640, RN => 
                           n6082, Q => registers_8_30_port, QN => net164000);
   registers_reg_8_29_inst : DFFR_X1 port map( D => n3780, CK => n640, RN => 
                           n6079, Q => registers_8_29_port, QN => net163999);
   registers_reg_8_28_inst : DFFR_X1 port map( D => n3779, CK => n640, RN => 
                           n6077, Q => registers_8_28_port, QN => net163998);
   registers_reg_8_27_inst : DFFR_X1 port map( D => n3778, CK => n640, RN => 
                           n6092, Q => registers_8_27_port, QN => net163997);
   registers_reg_8_26_inst : DFFR_X1 port map( D => n3777, CK => n640, RN => 
                           n6102, Q => registers_8_26_port, QN => net163996);
   registers_reg_8_25_inst : DFFR_X1 port map( D => n3776, CK => n640, RN => 
                           n6109, Q => registers_8_25_port, QN => net163995);
   registers_reg_8_24_inst : DFFR_X1 port map( D => n3775, CK => n640, RN => 
                           n6089, Q => registers_8_24_port, QN => net163994);
   registers_reg_8_23_inst : DFFR_X1 port map( D => n3774, CK => n640, RN => 
                           n6099, Q => registers_8_23_port, QN => net163993);
   registers_reg_8_22_inst : DFFR_X1 port map( D => n3773, CK => n640, RN => 
                           n6107, Q => registers_8_22_port, QN => net163992);
   registers_reg_8_21_inst : DFFR_X1 port map( D => n3772, CK => n640, RN => 
                           n6119, Q => registers_8_21_port, QN => net163991);
   registers_reg_8_20_inst : DFFR_X1 port map( D => n3771, CK => n640, RN => 
                           n6097, Q => registers_8_20_port, QN => net163990);
   registers_reg_8_19_inst : DFFR_X1 port map( D => n3770, CK => n640, RN => 
                           n6124, Q => registers_8_19_port, QN => net163989);
   registers_reg_8_18_inst : DFFR_X1 port map( D => n3769, CK => n640, RN => 
                           n6117, Q => registers_8_18_port, QN => net163988);
   registers_reg_8_17_inst : DFFR_X1 port map( D => n3768, CK => n640, RN => 
                           n6132, Q => registers_8_17_port, QN => net163987);
   registers_reg_8_16_inst : DFFR_X1 port map( D => n3767, CK => n640, RN => 
                           n6129, Q => registers_8_16_port, QN => net163986);
   registers_reg_8_15_inst : DFFR_X1 port map( D => n3766, CK => n640, RN => 
                           n6114, Q => registers_8_15_port, QN => net163985);
   registers_reg_8_14_inst : DFFR_X1 port map( D => n3765, CK => n640, RN => 
                           n6139, Q => registers_8_14_port, QN => net163984);
   registers_reg_8_13_inst : DFFR_X1 port map( D => n3764, CK => n640, RN => 
                           n6137, Q => registers_8_13_port, QN => net163983);
   registers_reg_8_12_inst : DFFR_X1 port map( D => n3763, CK => n640, RN => 
                           n6134, Q => registers_8_12_port, QN => net163982);
   registers_reg_8_11_inst : DFFR_X1 port map( D => n3762, CK => n640, RN => 
                           n6144, Q => registers_8_11_port, QN => net163981);
   registers_reg_8_10_inst : DFFR_X1 port map( D => n3761, CK => n640, RN => 
                           n6149, Q => registers_8_10_port, QN => net163980);
   registers_reg_8_9_inst : DFFR_X1 port map( D => n3760, CK => n640, RN => 
                           n6087, Q => registers_8_9_port, QN => net163979);
   registers_reg_8_8_inst : DFFR_X1 port map( D => n3759, CK => n640, RN => 
                           n6112, Q => registers_8_8_port, QN => net163978);
   registers_reg_8_7_inst : DFFR_X1 port map( D => n3758, CK => n640, RN => 
                           n6104, Q => registers_8_7_port, QN => net163977);
   registers_reg_8_6_inst : DFFR_X1 port map( D => n3757, CK => n640, RN => 
                           n6142, Q => registers_8_6_port, QN => net163976);
   registers_reg_8_5_inst : DFFR_X1 port map( D => n3756, CK => n640, RN => 
                           n6094, Q => registers_8_5_port, QN => net163975);
   registers_reg_8_4_inst : DFFR_X1 port map( D => n3755, CK => n640, RN => 
                           n6122, Q => registers_8_4_port, QN => net163974);
   registers_reg_8_3_inst : DFFR_X1 port map( D => n3754, CK => n640, RN => 
                           n6147, Q => registers_8_3_port, QN => net163973);
   registers_reg_8_2_inst : DFFR_X1 port map( D => n3753, CK => n640, RN => 
                           n6152, Q => registers_8_2_port, QN => net163972);
   registers_reg_8_1_inst : DFFR_X1 port map( D => n3752, CK => n640, RN => 
                           n6127, Q => registers_8_1_port, QN => net163971);
   registers_reg_8_0_inst : DFFR_X1 port map( D => n3751, CK => n640, RN => 
                           n6074, Q => registers_8_0_port, QN => net163970);
   registers_reg_9_31_inst : DFFR_X1 port map( D => n3750, CK => n640, RN => 
                           n6084, Q => registers_9_31_port, QN => n5121);
   registers_reg_9_30_inst : DFFR_X1 port map( D => n3749, CK => n640, RN => 
                           n6082, Q => registers_9_30_port, QN => n5120);
   registers_reg_9_29_inst : DFFR_X1 port map( D => n3748, CK => n640, RN => 
                           n6079, Q => registers_9_29_port, QN => n5119);
   registers_reg_9_28_inst : DFFR_X1 port map( D => n3747, CK => n640, RN => 
                           n6077, Q => registers_9_28_port, QN => n5118);
   registers_reg_9_27_inst : DFFR_X1 port map( D => n3746, CK => n640, RN => 
                           n6092, Q => registers_9_27_port, QN => n5117);
   registers_reg_9_26_inst : DFFR_X1 port map( D => n3745, CK => n640, RN => 
                           n6102, Q => registers_9_26_port, QN => n5116);
   registers_reg_9_25_inst : DFFR_X1 port map( D => n3744, CK => n640, RN => 
                           n6109, Q => registers_9_25_port, QN => n5115);
   registers_reg_9_24_inst : DFFR_X1 port map( D => n3743, CK => n640, RN => 
                           n6089, Q => registers_9_24_port, QN => n5114);
   registers_reg_9_23_inst : DFFR_X1 port map( D => n3742, CK => n640, RN => 
                           n6099, Q => registers_9_23_port, QN => n5113);
   registers_reg_9_22_inst : DFFR_X1 port map( D => n3741, CK => n640, RN => 
                           n6107, Q => registers_9_22_port, QN => n5112);
   registers_reg_9_21_inst : DFFR_X1 port map( D => n3740, CK => n640, RN => 
                           n6119, Q => registers_9_21_port, QN => n5111);
   registers_reg_9_20_inst : DFFR_X1 port map( D => n3739, CK => n640, RN => 
                           n6097, Q => registers_9_20_port, QN => n5110);
   registers_reg_9_19_inst : DFFR_X1 port map( D => n3738, CK => n640, RN => 
                           n6124, Q => registers_9_19_port, QN => n5109);
   registers_reg_9_18_inst : DFFR_X1 port map( D => n3737, CK => n640, RN => 
                           n6117, Q => registers_9_18_port, QN => n5108);
   registers_reg_9_17_inst : DFFR_X1 port map( D => n3736, CK => n640, RN => 
                           n6132, Q => registers_9_17_port, QN => n5107);
   registers_reg_9_16_inst : DFFR_X1 port map( D => n3735, CK => n640, RN => 
                           n6129, Q => registers_9_16_port, QN => n5106);
   registers_reg_9_15_inst : DFFR_X1 port map( D => n3734, CK => n640, RN => 
                           n6114, Q => registers_9_15_port, QN => n5105);
   registers_reg_9_14_inst : DFFR_X1 port map( D => n3733, CK => n640, RN => 
                           n6139, Q => registers_9_14_port, QN => n5104);
   registers_reg_9_13_inst : DFFR_X1 port map( D => n3732, CK => n640, RN => 
                           n6137, Q => registers_9_13_port, QN => n5103);
   registers_reg_9_12_inst : DFFR_X1 port map( D => n3731, CK => n640, RN => 
                           n6134, Q => registers_9_12_port, QN => n4431);
   registers_reg_9_11_inst : DFFR_X1 port map( D => n3730, CK => n640, RN => 
                           n6144, Q => registers_9_11_port, QN => n4416);
   registers_reg_9_10_inst : DFFR_X1 port map( D => n3729, CK => n640, RN => 
                           n6149, Q => registers_9_10_port, QN => n4394);
   registers_reg_9_9_inst : DFFR_X1 port map( D => n3728, CK => n640, RN => 
                           n6087, Q => registers_9_9_port, QN => n4375);
   registers_reg_9_8_inst : DFFR_X1 port map( D => n3727, CK => n640, RN => 
                           n6112, Q => registers_9_8_port, QN => n4356);
   registers_reg_9_7_inst : DFFR_X1 port map( D => n3726, CK => n640, RN => 
                           n6104, Q => registers_9_7_port, QN => n4337);
   registers_reg_9_6_inst : DFFR_X1 port map( D => n3725, CK => n640, RN => 
                           n6142, Q => registers_9_6_port, QN => n4318);
   registers_reg_9_5_inst : DFFR_X1 port map( D => n3724, CK => n640, RN => 
                           n6094, Q => registers_9_5_port, QN => n4299);
   registers_reg_9_4_inst : DFFR_X1 port map( D => n3723, CK => n640, RN => 
                           n6122, Q => registers_9_4_port, QN => n4280);
   registers_reg_9_3_inst : DFFR_X1 port map( D => n3722, CK => n640, RN => 
                           n6147, Q => registers_9_3_port, QN => n4261);
   registers_reg_9_2_inst : DFFR_X1 port map( D => n3721, CK => n640, RN => 
                           n6152, Q => registers_9_2_port, QN => n4242);
   registers_reg_9_1_inst : DFFR_X1 port map( D => n3720, CK => n640, RN => 
                           n6127, Q => registers_9_1_port, QN => n4223);
   registers_reg_9_0_inst : DFFR_X1 port map( D => n3719, CK => n640, RN => 
                           n6074, Q => registers_9_0_port, QN => n2387);
   registers_reg_10_31_inst : DFFR_X1 port map( D => n3718, CK => n640, RN => 
                           n6084, Q => net163969, QN => n2247);
   registers_reg_10_30_inst : DFFR_X1 port map( D => n3717, CK => n640, RN => 
                           n6082, Q => net163968, QN => n2246);
   registers_reg_10_29_inst : DFFR_X1 port map( D => n3716, CK => n640, RN => 
                           n6079, Q => net163967, QN => n2257);
   registers_reg_10_28_inst : DFFR_X1 port map( D => n3715, CK => n640, RN => 
                           n6077, Q => net163966, QN => n2245);
   registers_reg_10_27_inst : DFFR_X1 port map( D => n3714, CK => n640, RN => 
                           n6092, Q => net163965, QN => n2117);
   registers_reg_10_26_inst : DFFR_X1 port map( D => n3713, CK => n640, RN => 
                           n6102, Q => net163964, QN => n2118);
   registers_reg_10_25_inst : DFFR_X1 port map( D => n3712, CK => n640, RN => 
                           n6109, Q => net163963, QN => n2244);
   registers_reg_10_24_inst : DFFR_X1 port map( D => n3711, CK => n640, RN => 
                           n6089, Q => net163962, QN => n2243);
   registers_reg_10_23_inst : DFFR_X1 port map( D => n3710, CK => n640, RN => 
                           n6099, Q => net163961, QN => n2256);
   registers_reg_10_22_inst : DFFR_X1 port map( D => n3709, CK => n640, RN => 
                           n6107, Q => net163960, QN => n2242);
   registers_reg_10_21_inst : DFFR_X1 port map( D => n3708, CK => n640, RN => 
                           n6119, Q => net163959, QN => n2241);
   registers_reg_10_20_inst : DFFR_X1 port map( D => n3707, CK => n640, RN => 
                           n6097, Q => net163958, QN => n2255);
   registers_reg_10_19_inst : DFFR_X1 port map( D => n3706, CK => n640, RN => 
                           n6124, Q => net163957, QN => n2240);
   registers_reg_10_18_inst : DFFR_X1 port map( D => n3705, CK => n640, RN => 
                           n6117, Q => net163956, QN => n2239);
   registers_reg_10_17_inst : DFFR_X1 port map( D => n3704, CK => n640, RN => 
                           n6132, Q => net163955, QN => n2254);
   registers_reg_10_16_inst : DFFR_X1 port map( D => n3703, CK => n640, RN => 
                           n6130, Q => net163954, QN => n2238);
   registers_reg_10_15_inst : DFFR_X1 port map( D => n3702, CK => n640, RN => 
                           n6114, Q => net163953, QN => n2237);
   registers_reg_10_14_inst : DFFR_X1 port map( D => n3701, CK => n640, RN => 
                           n6140, Q => net163952, QN => n2253);
   registers_reg_10_13_inst : DFFR_X1 port map( D => n3700, CK => n640, RN => 
                           n6137, Q => net163951, QN => n2236);
   registers_reg_10_12_inst : DFFR_X1 port map( D => n3699, CK => n640, RN => 
                           n6135, Q => net163950, QN => n2235);
   registers_reg_10_11_inst : DFFR_X1 port map( D => n3698, CK => n640, RN => 
                           n6145, Q => net163949, QN => n2251);
   registers_reg_10_10_inst : DFFR_X1 port map( D => n3697, CK => n640, RN => 
                           n6150, Q => net163948, QN => n2234);
   registers_reg_10_9_inst : DFFR_X1 port map( D => n3696, CK => n640, RN => 
                           n6087, Q => net163947, QN => n2233);
   registers_reg_10_8_inst : DFFR_X1 port map( D => n3695, CK => n640, RN => 
                           n6112, Q => net163946, QN => n2250);
   registers_reg_10_7_inst : DFFR_X1 port map( D => n3694, CK => n640, RN => 
                           n6104, Q => net163945, QN => n2232);
   registers_reg_10_6_inst : DFFR_X1 port map( D => n3693, CK => n640, RN => 
                           n6142, Q => net163944, QN => n2231);
   registers_reg_10_5_inst : DFFR_X1 port map( D => n3692, CK => n640, RN => 
                           n6094, Q => net163943, QN => n2249);
   registers_reg_10_4_inst : DFFR_X1 port map( D => n3691, CK => n640, RN => 
                           n6122, Q => net163942, QN => n2230);
   registers_reg_10_3_inst : DFFR_X1 port map( D => n3690, CK => n640, RN => 
                           n6147, Q => net163941, QN => n2229);
   registers_reg_10_2_inst : DFFR_X1 port map( D => n3689, CK => n640, RN => 
                           n6152, Q => net163940, QN => n2248);
   registers_reg_10_1_inst : DFFR_X1 port map( D => n3688, CK => n640, RN => 
                           n6127, Q => net163939, QN => n2228);
   registers_reg_10_0_inst : DFFR_X1 port map( D => n3687, CK => n640, RN => 
                           n6074, Q => net163938, QN => n2226);
   registers_reg_11_31_inst : DFFR_X1 port map( D => n3686, CK => n640, RN => 
                           n6085, Q => registers_11_31_port, QN => n2929);
   registers_reg_11_30_inst : DFFR_X1 port map( D => n3685, CK => n640, RN => 
                           n6082, Q => registers_11_30_port, QN => n2928);
   registers_reg_11_29_inst : DFFR_X1 port map( D => n3684, CK => n640, RN => 
                           n6080, Q => registers_11_29_port, QN => n2927);
   registers_reg_11_28_inst : DFFR_X1 port map( D => n3683, CK => n640, RN => 
                           n6077, Q => registers_11_28_port, QN => n2926);
   registers_reg_11_27_inst : DFFR_X1 port map( D => n3682, CK => n640, RN => 
                           n6092, Q => registers_11_27_port, QN => n2925);
   registers_reg_11_26_inst : DFFR_X1 port map( D => n3681, CK => n640, RN => 
                           n6102, Q => registers_11_26_port, QN => n2924);
   registers_reg_11_25_inst : DFFR_X1 port map( D => n3680, CK => n640, RN => 
                           n6110, Q => registers_11_25_port, QN => n2923);
   registers_reg_11_24_inst : DFFR_X1 port map( D => n3679, CK => n640, RN => 
                           n6090, Q => registers_11_24_port, QN => n2922);
   registers_reg_11_23_inst : DFFR_X1 port map( D => n3678, CK => n640, RN => 
                           n6100, Q => registers_11_23_port, QN => n2813);
   registers_reg_11_22_inst : DFFR_X1 port map( D => n3677, CK => n640, RN => 
                           n6107, Q => registers_11_22_port, QN => n2794);
   registers_reg_11_21_inst : DFFR_X1 port map( D => n3676, CK => n640, RN => 
                           n6120, Q => registers_11_21_port, QN => n2775);
   registers_reg_11_20_inst : DFFR_X1 port map( D => n3675, CK => n640, RN => 
                           n6097, Q => registers_11_20_port, QN => n2756);
   registers_reg_11_19_inst : DFFR_X1 port map( D => n3674, CK => n640, RN => 
                           n6125, Q => registers_11_19_port, QN => n2701);
   registers_reg_11_18_inst : DFFR_X1 port map( D => n3673, CK => n640, RN => 
                           n6117, Q => registers_11_18_port, QN => n2698);
   registers_reg_11_17_inst : DFFR_X1 port map( D => n3672, CK => n640, RN => 
                           n6132, Q => registers_11_17_port, QN => n2697);
   registers_reg_11_16_inst : DFFR_X1 port map( D => n3671, CK => n640, RN => 
                           n6130, Q => registers_11_16_port, QN => n2696);
   registers_reg_11_15_inst : DFFR_X1 port map( D => n3670, CK => n640, RN => 
                           n6115, Q => registers_11_15_port, QN => n2695);
   registers_reg_11_14_inst : DFFR_X1 port map( D => n3669, CK => n640, RN => 
                           n6140, Q => registers_11_14_port, QN => n2694);
   registers_reg_11_13_inst : DFFR_X1 port map( D => n3668, CK => n640, RN => 
                           n6137, Q => registers_11_13_port, QN => n2693);
   registers_reg_11_12_inst : DFFR_X1 port map( D => n3667, CK => n640, RN => 
                           n6135, Q => registers_11_12_port, QN => n2692);
   registers_reg_11_11_inst : DFFR_X1 port map( D => n3666, CK => n640, RN => 
                           n6145, Q => registers_11_11_port, QN => n2691);
   registers_reg_11_10_inst : DFFR_X1 port map( D => n3665, CK => n640, RN => 
                           n6150, Q => registers_11_10_port, QN => n2690);
   registers_reg_11_9_inst : DFFR_X1 port map( D => n3664, CK => n640, RN => 
                           n6087, Q => registers_11_9_port, QN => n2689);
   registers_reg_11_8_inst : DFFR_X1 port map( D => n3663, CK => n640, RN => 
                           n6112, Q => registers_11_8_port, QN => n2688);
   registers_reg_11_7_inst : DFFR_X1 port map( D => n3662, CK => n640, RN => 
                           n6105, Q => registers_11_7_port, QN => n2687);
   registers_reg_11_6_inst : DFFR_X1 port map( D => n3661, CK => n640, RN => 
                           n6142, Q => registers_11_6_port, QN => n2686);
   registers_reg_11_5_inst : DFFR_X1 port map( D => n3660, CK => n640, RN => 
                           n6095, Q => registers_11_5_port, QN => n2685);
   registers_reg_11_4_inst : DFFR_X1 port map( D => n3659, CK => n640, RN => 
                           n6122, Q => registers_11_4_port, QN => n2684);
   registers_reg_11_3_inst : DFFR_X1 port map( D => n3658, CK => n640, RN => 
                           n6147, Q => registers_11_3_port, QN => n2683);
   registers_reg_11_2_inst : DFFR_X1 port map( D => n3657, CK => n640, RN => 
                           n6152, Q => registers_11_2_port, QN => n2682);
   registers_reg_11_1_inst : DFFR_X1 port map( D => n3656, CK => n640, RN => 
                           n6127, Q => registers_11_1_port, QN => n2681);
   registers_reg_11_0_inst : DFFR_X1 port map( D => n3655, CK => n640, RN => 
                           n6074, Q => registers_11_0_port, QN => n2680);
   registers_reg_12_31_inst : DFFR_X1 port map( D => n3654, CK => n640, RN => 
                           n6085, Q => net163937, QN => n2318);
   registers_reg_12_30_inst : DFFR_X1 port map( D => n3653, CK => n640, RN => 
                           n6082, Q => net163936, QN => n2317);
   registers_reg_12_29_inst : DFFR_X1 port map( D => n3652, CK => n640, RN => 
                           n6080, Q => net163935, QN => n2316);
   registers_reg_12_28_inst : DFFR_X1 port map( D => n3651, CK => n640, RN => 
                           n6077, Q => net163934, QN => n2315);
   registers_reg_12_27_inst : DFFR_X1 port map( D => n3650, CK => n640, RN => 
                           n6092, Q => net163933, QN => n2314);
   registers_reg_12_26_inst : DFFR_X1 port map( D => n3649, CK => n640, RN => 
                           n6102, Q => net163932, QN => n2313);
   registers_reg_12_25_inst : DFFR_X1 port map( D => n3648, CK => n640, RN => 
                           n6110, Q => net163931, QN => n2312);
   registers_reg_12_24_inst : DFFR_X1 port map( D => n3647, CK => n640, RN => 
                           n6090, Q => net163930, QN => n2311);
   registers_reg_12_23_inst : DFFR_X1 port map( D => n3646, CK => n640, RN => 
                           n6100, Q => net163929, QN => n2310);
   registers_reg_12_22_inst : DFFR_X1 port map( D => n3645, CK => n640, RN => 
                           n6107, Q => net163928, QN => n2309);
   registers_reg_12_21_inst : DFFR_X1 port map( D => n3644, CK => n640, RN => 
                           n6120, Q => net163927, QN => n2308);
   registers_reg_12_20_inst : DFFR_X1 port map( D => n3643, CK => n640, RN => 
                           n6097, Q => net163926, QN => n2307);
   registers_reg_12_19_inst : DFFR_X1 port map( D => n3642, CK => n640, RN => 
                           n6125, Q => net163925, QN => n2306);
   registers_reg_12_18_inst : DFFR_X1 port map( D => n3641, CK => n640, RN => 
                           n6117, Q => net163924, QN => n2305);
   registers_reg_12_17_inst : DFFR_X1 port map( D => n3640, CK => n640, RN => 
                           n6132, Q => net163923, QN => n2304);
   registers_reg_12_16_inst : DFFR_X1 port map( D => n3639, CK => n640, RN => 
                           n6130, Q => net163922, QN => n2303);
   registers_reg_12_15_inst : DFFR_X1 port map( D => n3638, CK => n640, RN => 
                           n6115, Q => net163921, QN => n2302);
   registers_reg_12_14_inst : DFFR_X1 port map( D => n3637, CK => n640, RN => 
                           n6140, Q => net163920, QN => n2301);
   registers_reg_12_13_inst : DFFR_X1 port map( D => n3636, CK => n640, RN => 
                           n6137, Q => net163919, QN => n2300);
   registers_reg_12_12_inst : DFFR_X1 port map( D => n3635, CK => n640, RN => 
                           n6135, Q => net163918, QN => n2299);
   registers_reg_12_11_inst : DFFR_X1 port map( D => n3634, CK => n640, RN => 
                           n6145, Q => net163917, QN => n2298);
   registers_reg_12_10_inst : DFFR_X1 port map( D => n3633, CK => n640, RN => 
                           n6150, Q => net163916, QN => n2297);
   registers_reg_12_9_inst : DFFR_X1 port map( D => n3632, CK => n640, RN => 
                           n6087, Q => net163915, QN => n2296);
   registers_reg_12_8_inst : DFFR_X1 port map( D => n3631, CK => n640, RN => 
                           n6112, Q => net163914, QN => n2295);
   registers_reg_12_7_inst : DFFR_X1 port map( D => n3630, CK => n640, RN => 
                           n6105, Q => net163913, QN => n2294);
   registers_reg_12_6_inst : DFFR_X1 port map( D => n3629, CK => n640, RN => 
                           n6142, Q => net163912, QN => n2293);
   registers_reg_12_5_inst : DFFR_X1 port map( D => n3628, CK => n640, RN => 
                           n6095, Q => net163911, QN => n2292);
   registers_reg_12_4_inst : DFFR_X1 port map( D => n3627, CK => n640, RN => 
                           n6122, Q => net163910, QN => n2291);
   registers_reg_12_3_inst : DFFR_X1 port map( D => n3626, CK => n640, RN => 
                           n6147, Q => net163909, QN => n2290);
   registers_reg_12_2_inst : DFFR_X1 port map( D => n3625, CK => n640, RN => 
                           n6152, Q => net163908, QN => n2289);
   registers_reg_12_1_inst : DFFR_X1 port map( D => n3624, CK => n640, RN => 
                           n6127, Q => net163907, QN => n2288);
   registers_reg_12_0_inst : DFFR_X1 port map( D => n3623, CK => n640, RN => 
                           n6074, Q => registers_12_0_port, QN => n5311);
   registers_reg_13_31_inst : DFFR_X1 port map( D => n3622, CK => n640, RN => 
                           n6085, Q => registers_13_31_port, QN => net163906);
   registers_reg_13_30_inst : DFFR_X1 port map( D => n3621, CK => n640, RN => 
                           n6082, Q => registers_13_30_port, QN => net163905);
   registers_reg_13_29_inst : DFFR_X1 port map( D => n3620, CK => n640, RN => 
                           n6080, Q => registers_13_29_port, QN => net163904);
   registers_reg_13_28_inst : DFFR_X1 port map( D => n3619, CK => n640, RN => 
                           n6077, Q => registers_13_28_port, QN => net163903);
   registers_reg_13_27_inst : DFFR_X1 port map( D => n3618, CK => n640, RN => 
                           n6092, Q => registers_13_27_port, QN => net163902);
   registers_reg_13_26_inst : DFFR_X1 port map( D => n3617, CK => n640, RN => 
                           n6102, Q => registers_13_26_port, QN => net163901);
   registers_reg_13_25_inst : DFFR_X1 port map( D => n3616, CK => n640, RN => 
                           n6110, Q => registers_13_25_port, QN => net163900);
   registers_reg_13_24_inst : DFFR_X1 port map( D => n3615, CK => n640, RN => 
                           n6090, Q => registers_13_24_port, QN => net163899);
   registers_reg_13_23_inst : DFFR_X1 port map( D => n3614, CK => n640, RN => 
                           n6100, Q => registers_13_23_port, QN => net163898);
   registers_reg_13_22_inst : DFFR_X1 port map( D => n3613, CK => n640, RN => 
                           n6107, Q => registers_13_22_port, QN => net163897);
   registers_reg_13_21_inst : DFFR_X1 port map( D => n3612, CK => n640, RN => 
                           n6120, Q => registers_13_21_port, QN => net163896);
   registers_reg_13_20_inst : DFFR_X1 port map( D => n3611, CK => n640, RN => 
                           n6097, Q => registers_13_20_port, QN => net163895);
   registers_reg_13_19_inst : DFFR_X1 port map( D => n3610, CK => n640, RN => 
                           n6125, Q => registers_13_19_port, QN => net163894);
   registers_reg_13_18_inst : DFFR_X1 port map( D => n3609, CK => n640, RN => 
                           n6117, Q => registers_13_18_port, QN => net163893);
   registers_reg_13_17_inst : DFFR_X1 port map( D => n3608, CK => n640, RN => 
                           n6132, Q => registers_13_17_port, QN => net163892);
   registers_reg_13_16_inst : DFFR_X1 port map( D => n3607, CK => n640, RN => 
                           n6130, Q => registers_13_16_port, QN => net163891);
   registers_reg_13_15_inst : DFFR_X1 port map( D => n3606, CK => n640, RN => 
                           n6115, Q => registers_13_15_port, QN => net163890);
   registers_reg_13_14_inst : DFFR_X1 port map( D => n3605, CK => n640, RN => 
                           n6140, Q => registers_13_14_port, QN => net163889);
   registers_reg_13_13_inst : DFFR_X1 port map( D => n3604, CK => n640, RN => 
                           n6137, Q => registers_13_13_port, QN => net163888);
   registers_reg_13_12_inst : DFFR_X1 port map( D => n3603, CK => n640, RN => 
                           n6135, Q => registers_13_12_port, QN => net163887);
   registers_reg_13_11_inst : DFFR_X1 port map( D => n3602, CK => n640, RN => 
                           n6145, Q => registers_13_11_port, QN => net163886);
   registers_reg_13_10_inst : DFFR_X1 port map( D => n3601, CK => n640, RN => 
                           n6150, Q => registers_13_10_port, QN => net163885);
   registers_reg_13_9_inst : DFFR_X1 port map( D => n3600, CK => n640, RN => 
                           n6087, Q => registers_13_9_port, QN => net163884);
   registers_reg_13_8_inst : DFFR_X1 port map( D => n3599, CK => n640, RN => 
                           n6112, Q => registers_13_8_port, QN => net163883);
   registers_reg_13_7_inst : DFFR_X1 port map( D => n3598, CK => n640, RN => 
                           n6105, Q => registers_13_7_port, QN => net163882);
   registers_reg_13_6_inst : DFFR_X1 port map( D => n3597, CK => n640, RN => 
                           n6142, Q => registers_13_6_port, QN => net163881);
   registers_reg_13_5_inst : DFFR_X1 port map( D => n3596, CK => n640, RN => 
                           n6095, Q => registers_13_5_port, QN => net163880);
   registers_reg_13_4_inst : DFFR_X1 port map( D => n3595, CK => n640, RN => 
                           n6122, Q => registers_13_4_port, QN => net163879);
   registers_reg_13_3_inst : DFFR_X1 port map( D => n3594, CK => n640, RN => 
                           n6147, Q => registers_13_3_port, QN => net163878);
   registers_reg_13_2_inst : DFFR_X1 port map( D => n3593, CK => n640, RN => 
                           n6152, Q => registers_13_2_port, QN => net163877);
   registers_reg_13_1_inst : DFFR_X1 port map( D => n3592, CK => n640, RN => 
                           n6127, Q => registers_13_1_port, QN => net163876);
   registers_reg_13_0_inst : DFFR_X1 port map( D => n3591, CK => n640, RN => 
                           n6075, Q => registers_13_0_port, QN => n2479);
   registers_reg_14_31_inst : DFFR_X1 port map( D => n3590, CK => n640, RN => 
                           n6085, Q => registers_14_31_port, QN => n2352);
   registers_reg_14_30_inst : DFFR_X1 port map( D => n3589, CK => n640, RN => 
                           n6082, Q => registers_14_30_port, QN => n2351);
   registers_reg_14_29_inst : DFFR_X1 port map( D => n3588, CK => n640, RN => 
                           n6080, Q => registers_14_29_port, QN => n2350);
   registers_reg_14_28_inst : DFFR_X1 port map( D => n3587, CK => n640, RN => 
                           n6077, Q => registers_14_28_port, QN => n2349);
   registers_reg_14_27_inst : DFFR_X1 port map( D => n3586, CK => n640, RN => 
                           n6092, Q => registers_14_27_port, QN => n2348);
   registers_reg_14_26_inst : DFFR_X1 port map( D => n3585, CK => n640, RN => 
                           n6102, Q => registers_14_26_port, QN => n2347);
   registers_reg_14_25_inst : DFFR_X1 port map( D => n3584, CK => n640, RN => 
                           n6110, Q => registers_14_25_port, QN => n2346);
   registers_reg_14_24_inst : DFFR_X1 port map( D => n3583, CK => n640, RN => 
                           n6090, Q => registers_14_24_port, QN => n2345);
   registers_reg_14_23_inst : DFFR_X1 port map( D => n3582, CK => n640, RN => 
                           n6100, Q => registers_14_23_port, QN => n2344);
   registers_reg_14_22_inst : DFFR_X1 port map( D => n3581, CK => n640, RN => 
                           n6107, Q => registers_14_22_port, QN => n2343);
   registers_reg_14_21_inst : DFFR_X1 port map( D => n3580, CK => n640, RN => 
                           n6120, Q => registers_14_21_port, QN => n2342);
   registers_reg_14_20_inst : DFFR_X1 port map( D => n3579, CK => n640, RN => 
                           n6097, Q => registers_14_20_port, QN => n2341);
   registers_reg_14_19_inst : DFFR_X1 port map( D => n3578, CK => n640, RN => 
                           n6125, Q => registers_14_19_port, QN => n2340);
   registers_reg_14_18_inst : DFFR_X1 port map( D => n3577, CK => n640, RN => 
                           n6117, Q => registers_14_18_port, QN => n2339);
   registers_reg_14_17_inst : DFFR_X1 port map( D => n3576, CK => n640, RN => 
                           n6132, Q => registers_14_17_port, QN => n2338);
   registers_reg_14_16_inst : DFFR_X1 port map( D => n3575, CK => n640, RN => 
                           n6130, Q => registers_14_16_port, QN => n2337);
   registers_reg_14_15_inst : DFFR_X1 port map( D => n3574, CK => n640, RN => 
                           n6115, Q => registers_14_15_port, QN => n2336);
   registers_reg_14_14_inst : DFFR_X1 port map( D => n3573, CK => n640, RN => 
                           n6140, Q => registers_14_14_port, QN => n2335);
   registers_reg_14_13_inst : DFFR_X1 port map( D => n3572, CK => n640, RN => 
                           n6137, Q => registers_14_13_port, QN => n2334);
   registers_reg_14_12_inst : DFFR_X1 port map( D => n3571, CK => n640, RN => 
                           n6135, Q => registers_14_12_port, QN => n2333);
   registers_reg_14_11_inst : DFFR_X1 port map( D => n3570, CK => n640, RN => 
                           n6145, Q => registers_14_11_port, QN => n2332);
   registers_reg_14_10_inst : DFFR_X1 port map( D => n3569, CK => n640, RN => 
                           n6150, Q => registers_14_10_port, QN => n2331);
   registers_reg_14_9_inst : DFFR_X1 port map( D => n3568, CK => n640, RN => 
                           n6087, Q => registers_14_9_port, QN => n2330);
   registers_reg_14_8_inst : DFFR_X1 port map( D => n3567, CK => n640, RN => 
                           n6112, Q => registers_14_8_port, QN => n2329);
   registers_reg_14_7_inst : DFFR_X1 port map( D => n3566, CK => n640, RN => 
                           n6105, Q => registers_14_7_port, QN => n2328);
   registers_reg_14_6_inst : DFFR_X1 port map( D => n3565, CK => n640, RN => 
                           n6142, Q => registers_14_6_port, QN => n2327);
   registers_reg_14_5_inst : DFFR_X1 port map( D => n3564, CK => n640, RN => 
                           n6095, Q => registers_14_5_port, QN => n2326);
   registers_reg_14_4_inst : DFFR_X1 port map( D => n3563, CK => n640, RN => 
                           n6122, Q => registers_14_4_port, QN => n2325);
   registers_reg_14_3_inst : DFFR_X1 port map( D => n3562, CK => n640, RN => 
                           n6147, Q => registers_14_3_port, QN => n2324);
   registers_reg_14_2_inst : DFFR_X1 port map( D => n3561, CK => n640, RN => 
                           n6152, Q => registers_14_2_port, QN => n2323);
   registers_reg_14_1_inst : DFFR_X1 port map( D => n3560, CK => n640, RN => 
                           n6127, Q => registers_14_1_port, QN => n2322);
   registers_reg_14_0_inst : DFFR_X1 port map( D => n3559, CK => n640, RN => 
                           n6075, Q => registers_14_0_port, QN => n2319);
   registers_reg_15_31_inst : DFFR_X1 port map( D => n3558, CK => n640, RN => 
                           n6085, Q => registers_15_31_port, QN => n2653);
   registers_reg_15_30_inst : DFFR_X1 port map( D => n3557, CK => n640, RN => 
                           n6082, Q => registers_15_30_port, QN => n2652);
   registers_reg_15_29_inst : DFFR_X1 port map( D => n3556, CK => n640, RN => 
                           n6080, Q => registers_15_29_port, QN => n2651);
   registers_reg_15_28_inst : DFFR_X1 port map( D => n3555, CK => n640, RN => 
                           n6077, Q => registers_15_28_port, QN => n2650);
   registers_reg_15_27_inst : DFFR_X1 port map( D => n3554, CK => n640, RN => 
                           n6092, Q => registers_15_27_port, QN => n2649);
   registers_reg_15_26_inst : DFFR_X1 port map( D => n3553, CK => n640, RN => 
                           n6102, Q => registers_15_26_port, QN => n2648);
   registers_reg_15_25_inst : DFFR_X1 port map( D => n3552, CK => n640, RN => 
                           n6110, Q => registers_15_25_port, QN => n2613);
   registers_reg_15_24_inst : DFFR_X1 port map( D => n3551, CK => n640, RN => 
                           n6090, Q => registers_15_24_port, QN => n2612);
   registers_reg_15_23_inst : DFFR_X1 port map( D => n3550, CK => n640, RN => 
                           n6100, Q => registers_15_23_port, QN => n2611);
   registers_reg_15_22_inst : DFFR_X1 port map( D => n3549, CK => n640, RN => 
                           n6107, Q => registers_15_22_port, QN => n2610);
   registers_reg_15_21_inst : DFFR_X1 port map( D => n3548, CK => n640, RN => 
                           n6120, Q => registers_15_21_port, QN => n2609);
   registers_reg_15_20_inst : DFFR_X1 port map( D => n3547, CK => n640, RN => 
                           n6097, Q => registers_15_20_port, QN => n2608);
   registers_reg_15_19_inst : DFFR_X1 port map( D => n3546, CK => n640, RN => 
                           n6125, Q => registers_15_19_port, QN => n2607);
   registers_reg_15_18_inst : DFFR_X1 port map( D => n3545, CK => n640, RN => 
                           n6117, Q => registers_15_18_port, QN => n2606);
   registers_reg_15_17_inst : DFFR_X1 port map( D => n3544, CK => n640, RN => 
                           n6132, Q => registers_15_17_port, QN => n2605);
   registers_reg_15_16_inst : DFFR_X1 port map( D => n3543, CK => n640, RN => 
                           n6130, Q => registers_15_16_port, QN => n2604);
   registers_reg_15_15_inst : DFFR_X1 port map( D => n3542, CK => n640, RN => 
                           n6115, Q => registers_15_15_port, QN => n2603);
   registers_reg_15_14_inst : DFFR_X1 port map( D => n3541, CK => n640, RN => 
                           n6140, Q => registers_15_14_port, QN => n2602);
   registers_reg_15_13_inst : DFFR_X1 port map( D => n3540, CK => n640, RN => 
                           n6137, Q => registers_15_13_port, QN => n2601);
   registers_reg_15_12_inst : DFFR_X1 port map( D => n3539, CK => n640, RN => 
                           n6135, Q => registers_15_12_port, QN => n2600);
   registers_reg_15_11_inst : DFFR_X1 port map( D => n3538, CK => n640, RN => 
                           n6145, Q => registers_15_11_port, QN => n2599);
   registers_reg_15_10_inst : DFFR_X1 port map( D => n3537, CK => n640, RN => 
                           n6150, Q => registers_15_10_port, QN => n2598);
   registers_reg_15_9_inst : DFFR_X1 port map( D => n3536, CK => n640, RN => 
                           n6087, Q => registers_15_9_port, QN => n2597);
   registers_reg_15_8_inst : DFFR_X1 port map( D => n3535, CK => n640, RN => 
                           n6112, Q => registers_15_8_port, QN => n2596);
   registers_reg_15_7_inst : DFFR_X1 port map( D => n3534, CK => n640, RN => 
                           n6105, Q => registers_15_7_port, QN => n2594);
   registers_reg_15_6_inst : DFFR_X1 port map( D => n3533, CK => n640, RN => 
                           n6142, Q => registers_15_6_port, QN => n2593);
   registers_reg_15_5_inst : DFFR_X1 port map( D => n3532, CK => n640, RN => 
                           n6095, Q => registers_15_5_port, QN => n2592);
   registers_reg_15_4_inst : DFFR_X1 port map( D => n3531, CK => n640, RN => 
                           n6122, Q => registers_15_4_port, QN => n2591);
   registers_reg_15_3_inst : DFFR_X1 port map( D => n3530, CK => n640, RN => 
                           n6147, Q => registers_15_3_port, QN => n2590);
   registers_reg_15_2_inst : DFFR_X1 port map( D => n3529, CK => n640, RN => 
                           n6152, Q => registers_15_2_port, QN => n2589);
   registers_reg_15_1_inst : DFFR_X1 port map( D => n3528, CK => n640, RN => 
                           n6127, Q => registers_15_1_port, QN => n2588);
   registers_reg_15_0_inst : DFFR_X1 port map( D => n3527, CK => n640, RN => 
                           n6075, Q => registers_15_0_port, QN => net108355);
   registers_reg_16_31_inst : DFFR_X1 port map( D => n3526, CK => n640, RN => 
                           n6085, Q => registers_16_31_port, QN => n5204);
   registers_reg_16_30_inst : DFFR_X1 port map( D => n3525, CK => n640, RN => 
                           n6082, Q => registers_16_30_port, QN => n5203);
   registers_reg_16_29_inst : DFFR_X1 port map( D => n3524, CK => n640, RN => 
                           n6080, Q => registers_16_29_port, QN => n5214);
   registers_reg_16_28_inst : DFFR_X1 port map( D => n3523, CK => n640, RN => 
                           n6077, Q => registers_16_28_port, QN => n5202);
   registers_reg_16_27_inst : DFFR_X1 port map( D => n3522, CK => n640, RN => 
                           n6092, Q => registers_16_27_port, QN => n5201);
   registers_reg_16_26_inst : DFFR_X1 port map( D => n3521, CK => n640, RN => 
                           n6102, Q => registers_16_26_port, QN => n5213);
   registers_reg_16_25_inst : DFFR_X1 port map( D => n3520, CK => n640, RN => 
                           n6110, Q => registers_16_25_port, QN => n5200);
   registers_reg_16_24_inst : DFFR_X1 port map( D => n3519, CK => n640, RN => 
                           n6090, Q => registers_16_24_port, QN => n5199);
   registers_reg_16_23_inst : DFFR_X1 port map( D => n3518, CK => n640, RN => 
                           n6100, Q => registers_16_23_port, QN => n5212);
   registers_reg_16_22_inst : DFFR_X1 port map( D => n3517, CK => n640, RN => 
                           n6107, Q => registers_16_22_port, QN => n5198);
   registers_reg_16_21_inst : DFFR_X1 port map( D => n3516, CK => n640, RN => 
                           n6120, Q => registers_16_21_port, QN => n5197);
   registers_reg_16_20_inst : DFFR_X1 port map( D => n3515, CK => n640, RN => 
                           n6097, Q => registers_16_20_port, QN => n5211);
   registers_reg_16_19_inst : DFFR_X1 port map( D => n3514, CK => n640, RN => 
                           n6125, Q => registers_16_19_port, QN => n5196);
   registers_reg_16_18_inst : DFFR_X1 port map( D => n3513, CK => n640, RN => 
                           n6117, Q => registers_16_18_port, QN => n5195);
   registers_reg_16_17_inst : DFFR_X1 port map( D => n3512, CK => n640, RN => 
                           n6133, Q => registers_16_17_port, QN => n5210);
   registers_reg_16_16_inst : DFFR_X1 port map( D => n3511, CK => n640, RN => 
                           n6130, Q => registers_16_16_port, QN => n5194);
   registers_reg_16_15_inst : DFFR_X1 port map( D => n3510, CK => n640, RN => 
                           n6115, Q => registers_16_15_port, QN => n5193);
   registers_reg_16_14_inst : DFFR_X1 port map( D => n3509, CK => n640, RN => 
                           n6140, Q => registers_16_14_port, QN => n5209);
   registers_reg_16_13_inst : DFFR_X1 port map( D => n3508, CK => n640, RN => 
                           n6138, Q => registers_16_13_port, QN => n5192);
   registers_reg_16_12_inst : DFFR_X1 port map( D => n3507, CK => n640, RN => 
                           n6135, Q => registers_16_12_port, QN => n5191);
   registers_reg_16_11_inst : DFFR_X1 port map( D => n3506, CK => n640, RN => 
                           n6145, Q => registers_16_11_port, QN => n5208);
   registers_reg_16_10_inst : DFFR_X1 port map( D => n3505, CK => n640, RN => 
                           n6150, Q => registers_16_10_port, QN => n5190);
   registers_reg_16_9_inst : DFFR_X1 port map( D => n3504, CK => n640, RN => 
                           n6087, Q => registers_16_9_port, QN => n5189);
   registers_reg_16_8_inst : DFFR_X1 port map( D => n3503, CK => n640, RN => 
                           n6112, Q => registers_16_8_port, QN => n5207);
   registers_reg_16_7_inst : DFFR_X1 port map( D => n3502, CK => n640, RN => 
                           n6105, Q => registers_16_7_port, QN => n5188);
   registers_reg_16_6_inst : DFFR_X1 port map( D => n3501, CK => n640, RN => 
                           n6143, Q => registers_16_6_port, QN => n5187);
   registers_reg_16_5_inst : DFFR_X1 port map( D => n3500, CK => n640, RN => 
                           n6095, Q => registers_16_5_port, QN => n5206);
   registers_reg_16_4_inst : DFFR_X1 port map( D => n3499, CK => n640, RN => 
                           n6122, Q => registers_16_4_port, QN => n5186);
   registers_reg_16_3_inst : DFFR_X1 port map( D => n3498, CK => n640, RN => 
                           n6148, Q => registers_16_3_port, QN => n5185);
   registers_reg_16_2_inst : DFFR_X1 port map( D => n3497, CK => n640, RN => 
                           n6153, Q => registers_16_2_port, QN => n5205);
   registers_reg_16_1_inst : DFFR_X1 port map( D => n3496, CK => n640, RN => 
                           n6127, Q => registers_16_1_port, QN => n5184);
   registers_reg_16_0_inst : DFFR_X1 port map( D => n3495, CK => n640, RN => 
                           n6075, Q => registers_16_0_port, QN => n2154);
   registers_reg_17_31_inst : DFFR_X1 port map( D => n3494, CK => n640, RN => 
                           n6085, Q => registers_17_31_port, QN => n2444);
   registers_reg_17_30_inst : DFFR_X1 port map( D => n3493, CK => n640, RN => 
                           n6083, Q => registers_17_30_port, QN => n2443);
   registers_reg_17_29_inst : DFFR_X1 port map( D => n3492, CK => n640, RN => 
                           n6080, Q => registers_17_29_port, QN => n2454);
   registers_reg_17_28_inst : DFFR_X1 port map( D => n3491, CK => n640, RN => 
                           n6078, Q => registers_17_28_port, QN => n2442);
   registers_reg_17_27_inst : DFFR_X1 port map( D => n3490, CK => n640, RN => 
                           n6093, Q => registers_17_27_port, QN => n2441);
   registers_reg_17_26_inst : DFFR_X1 port map( D => n3489, CK => n640, RN => 
                           n6103, Q => registers_17_26_port, QN => n2453);
   registers_reg_17_25_inst : DFFR_X1 port map( D => n3488, CK => n640, RN => 
                           n6110, Q => registers_17_25_port, QN => n2440);
   registers_reg_17_24_inst : DFFR_X1 port map( D => n3487, CK => n640, RN => 
                           n6090, Q => registers_17_24_port, QN => n2439);
   registers_reg_17_23_inst : DFFR_X1 port map( D => n3486, CK => n640, RN => 
                           n6100, Q => registers_17_23_port, QN => n2452);
   registers_reg_17_22_inst : DFFR_X1 port map( D => n3485, CK => n640, RN => 
                           n6108, Q => registers_17_22_port, QN => n2438);
   registers_reg_17_21_inst : DFFR_X1 port map( D => n3484, CK => n640, RN => 
                           n6120, Q => registers_17_21_port, QN => n2437);
   registers_reg_17_20_inst : DFFR_X1 port map( D => n3483, CK => n640, RN => 
                           n6098, Q => registers_17_20_port, QN => n2451);
   registers_reg_17_19_inst : DFFR_X1 port map( D => n3482, CK => n640, RN => 
                           n6125, Q => registers_17_19_port, QN => n2436);
   registers_reg_17_18_inst : DFFR_X1 port map( D => n3481, CK => n640, RN => 
                           n6118, Q => registers_17_18_port, QN => n2435);
   registers_reg_17_17_inst : DFFR_X1 port map( D => n3480, CK => n640, RN => 
                           n6133, Q => registers_17_17_port, QN => n2450);
   registers_reg_17_16_inst : DFFR_X1 port map( D => n3479, CK => n640, RN => 
                           n6130, Q => registers_17_16_port, QN => n2434);
   registers_reg_17_15_inst : DFFR_X1 port map( D => n3478, CK => n640, RN => 
                           n6115, Q => registers_17_15_port, QN => n2433);
   registers_reg_17_14_inst : DFFR_X1 port map( D => n3477, CK => n640, RN => 
                           n6140, Q => registers_17_14_port, QN => n2449);
   registers_reg_17_13_inst : DFFR_X1 port map( D => n3476, CK => n640, RN => 
                           n6138, Q => registers_17_13_port, QN => n2432);
   registers_reg_17_12_inst : DFFR_X1 port map( D => n3475, CK => n640, RN => 
                           n6135, Q => registers_17_12_port, QN => n2431);
   registers_reg_17_11_inst : DFFR_X1 port map( D => n3474, CK => n640, RN => 
                           n6145, Q => registers_17_11_port, QN => n2448);
   registers_reg_17_10_inst : DFFR_X1 port map( D => n3473, CK => n640, RN => 
                           n6150, Q => registers_17_10_port, QN => n2430);
   registers_reg_17_9_inst : DFFR_X1 port map( D => n3472, CK => n640, RN => 
                           n6088, Q => registers_17_9_port, QN => n2429);
   registers_reg_17_8_inst : DFFR_X1 port map( D => n3471, CK => n640, RN => 
                           n6113, Q => registers_17_8_port, QN => n2447);
   registers_reg_17_7_inst : DFFR_X1 port map( D => n3470, CK => n640, RN => 
                           n6105, Q => registers_17_7_port, QN => n2428);
   registers_reg_17_6_inst : DFFR_X1 port map( D => n3469, CK => n640, RN => 
                           n6143, Q => registers_17_6_port, QN => n2427);
   registers_reg_17_5_inst : DFFR_X1 port map( D => n3468, CK => n640, RN => 
                           n6095, Q => registers_17_5_port, QN => n2446);
   registers_reg_17_4_inst : DFFR_X1 port map( D => n3467, CK => n640, RN => 
                           n6123, Q => registers_17_4_port, QN => n2426);
   registers_reg_17_3_inst : DFFR_X1 port map( D => n3466, CK => n640, RN => 
                           n6148, Q => registers_17_3_port, QN => n2425);
   registers_reg_17_2_inst : DFFR_X1 port map( D => n3465, CK => n640, RN => 
                           n6153, Q => registers_17_2_port, QN => n2445);
   registers_reg_17_1_inst : DFFR_X1 port map( D => n3464, CK => n640, RN => 
                           n6128, Q => registers_17_1_port, QN => n2423);
   registers_reg_17_0_inst : DFFR_X1 port map( D => n3463, CK => n640, RN => 
                           n6075, Q => registers_17_0_port, QN => n5238);
   registers_reg_18_31_inst : DFFR_X1 port map( D => n3462, CK => n640, RN => 
                           n6085, Q => net163875, QN => n2222);
   registers_reg_18_30_inst : DFFR_X1 port map( D => n3461, CK => n640, RN => 
                           n6083, Q => net163874, QN => n2221);
   registers_reg_18_29_inst : DFFR_X1 port map( D => n3460, CK => n640, RN => 
                           n6080, Q => net163873, QN => n2220);
   registers_reg_18_28_inst : DFFR_X1 port map( D => n3459, CK => n640, RN => 
                           n6078, Q => net163872, QN => n2219);
   registers_reg_18_27_inst : DFFR_X1 port map( D => n3458, CK => n640, RN => 
                           n6093, Q => net163871, QN => n2216);
   registers_reg_18_26_inst : DFFR_X1 port map( D => n3457, CK => n640, RN => 
                           n6103, Q => net163870, QN => n2215);
   registers_reg_18_25_inst : DFFR_X1 port map( D => n3456, CK => n640, RN => 
                           n6110, Q => net163869, QN => n2214);
   registers_reg_18_24_inst : DFFR_X1 port map( D => n3455, CK => n640, RN => 
                           n6090, Q => net163868, QN => n2213);
   registers_reg_18_23_inst : DFFR_X1 port map( D => n3454, CK => n640, RN => 
                           n6100, Q => net163867, QN => n2212);
   registers_reg_18_22_inst : DFFR_X1 port map( D => n3453, CK => n640, RN => 
                           n6108, Q => net163866, QN => n2211);
   registers_reg_18_21_inst : DFFR_X1 port map( D => n3452, CK => n640, RN => 
                           n6120, Q => net163865, QN => n2210);
   registers_reg_18_20_inst : DFFR_X1 port map( D => n3451, CK => n640, RN => 
                           n6098, Q => net163864, QN => n2209);
   registers_reg_18_19_inst : DFFR_X1 port map( D => n3450, CK => n640, RN => 
                           n6125, Q => net163863, QN => n2208);
   registers_reg_18_18_inst : DFFR_X1 port map( D => n3449, CK => n640, RN => 
                           n6118, Q => net163862, QN => n2207);
   registers_reg_18_17_inst : DFFR_X1 port map( D => n3448, CK => n640, RN => 
                           n6133, Q => net163861, QN => n2206);
   registers_reg_18_16_inst : DFFR_X1 port map( D => n3447, CK => n640, RN => 
                           n6130, Q => net163860, QN => n2205);
   registers_reg_18_15_inst : DFFR_X1 port map( D => n3446, CK => n640, RN => 
                           n6115, Q => net163859, QN => n2204);
   registers_reg_18_14_inst : DFFR_X1 port map( D => n3445, CK => n640, RN => 
                           n6140, Q => net163858, QN => n2203);
   registers_reg_18_13_inst : DFFR_X1 port map( D => n3444, CK => n640, RN => 
                           n6138, Q => net163857, QN => n2202);
   registers_reg_18_12_inst : DFFR_X1 port map( D => n3443, CK => n640, RN => 
                           n6135, Q => net163856, QN => n2201);
   registers_reg_18_11_inst : DFFR_X1 port map( D => n3442, CK => n640, RN => 
                           n6145, Q => net163855, QN => n2200);
   registers_reg_18_10_inst : DFFR_X1 port map( D => n3441, CK => n640, RN => 
                           n6150, Q => net163854, QN => n2199);
   registers_reg_18_9_inst : DFFR_X1 port map( D => n3440, CK => n640, RN => 
                           n6088, Q => net163853, QN => n2198);
   registers_reg_18_8_inst : DFFR_X1 port map( D => n3439, CK => n640, RN => 
                           n6113, Q => net163852, QN => n2197);
   registers_reg_18_7_inst : DFFR_X1 port map( D => n3438, CK => n640, RN => 
                           n6105, Q => net163851, QN => n2196);
   registers_reg_18_6_inst : DFFR_X1 port map( D => n3437, CK => n640, RN => 
                           n6143, Q => net163850, QN => n2195);
   registers_reg_18_5_inst : DFFR_X1 port map( D => n3436, CK => n640, RN => 
                           n6095, Q => net163849, QN => n2194);
   registers_reg_18_4_inst : DFFR_X1 port map( D => n3435, CK => n640, RN => 
                           n6123, Q => net163848, QN => n2193);
   registers_reg_18_3_inst : DFFR_X1 port map( D => n3434, CK => n640, RN => 
                           n6148, Q => net163847, QN => n2192);
   registers_reg_18_2_inst : DFFR_X1 port map( D => n3433, CK => n640, RN => 
                           n6153, Q => net163846, QN => n2191);
   registers_reg_18_1_inst : DFFR_X1 port map( D => n3432, CK => n640, RN => 
                           n6128, Q => net163845, QN => n2190);
   registers_reg_18_0_inst : DFFR_X1 port map( D => n3431, CK => n640, RN => 
                           n6075, Q => net163844, QN => n2225);
   registers_reg_19_31_inst : DFFR_X1 port map( D => n3430, CK => n640, RN => 
                           n6085, Q => registers_19_31_port, QN => n2421);
   registers_reg_19_30_inst : DFFR_X1 port map( D => n3429, CK => n640, RN => 
                           n6083, Q => registers_19_30_port, QN => n2420);
   registers_reg_19_29_inst : DFFR_X1 port map( D => n3428, CK => n640, RN => 
                           n6080, Q => registers_19_29_port, QN => n2419);
   registers_reg_19_28_inst : DFFR_X1 port map( D => n3427, CK => n640, RN => 
                           n6078, Q => registers_19_28_port, QN => n2418);
   registers_reg_19_27_inst : DFFR_X1 port map( D => n3426, CK => n640, RN => 
                           n6093, Q => registers_19_27_port, QN => n2417);
   registers_reg_19_26_inst : DFFR_X1 port map( D => n3425, CK => n640, RN => 
                           n6103, Q => registers_19_26_port, QN => n2416);
   registers_reg_19_25_inst : DFFR_X1 port map( D => n3424, CK => n640, RN => 
                           n6110, Q => registers_19_25_port, QN => n2415);
   registers_reg_19_24_inst : DFFR_X1 port map( D => n3423, CK => n640, RN => 
                           n6090, Q => registers_19_24_port, QN => n2414);
   registers_reg_19_23_inst : DFFR_X1 port map( D => n3422, CK => n640, RN => 
                           n6100, Q => registers_19_23_port, QN => n2413);
   registers_reg_19_22_inst : DFFR_X1 port map( D => n3421, CK => n640, RN => 
                           n6108, Q => registers_19_22_port, QN => n2412);
   registers_reg_19_21_inst : DFFR_X1 port map( D => n3420, CK => n640, RN => 
                           n6120, Q => registers_19_21_port, QN => n2411);
   registers_reg_19_20_inst : DFFR_X1 port map( D => n3419, CK => n640, RN => 
                           n6098, Q => registers_19_20_port, QN => n2410);
   registers_reg_19_19_inst : DFFR_X1 port map( D => n3418, CK => n640, RN => 
                           n6125, Q => registers_19_19_port, QN => n2409);
   registers_reg_19_18_inst : DFFR_X1 port map( D => n3417, CK => n640, RN => 
                           n6118, Q => registers_19_18_port, QN => n2408);
   registers_reg_19_17_inst : DFFR_X1 port map( D => n3416, CK => n640, RN => 
                           n6133, Q => registers_19_17_port, QN => n2407);
   registers_reg_19_16_inst : DFFR_X1 port map( D => n3415, CK => n640, RN => 
                           n6130, Q => registers_19_16_port, QN => n2406);
   registers_reg_19_15_inst : DFFR_X1 port map( D => n3414, CK => n640, RN => 
                           n6115, Q => registers_19_15_port, QN => n2405);
   registers_reg_19_14_inst : DFFR_X1 port map( D => n3413, CK => n640, RN => 
                           n6140, Q => registers_19_14_port, QN => n2404);
   registers_reg_19_13_inst : DFFR_X1 port map( D => n3412, CK => n640, RN => 
                           n6138, Q => registers_19_13_port, QN => n2403);
   registers_reg_19_12_inst : DFFR_X1 port map( D => n3411, CK => n640, RN => 
                           n6135, Q => registers_19_12_port, QN => n2402);
   registers_reg_19_11_inst : DFFR_X1 port map( D => n3410, CK => n640, RN => 
                           n6145, Q => registers_19_11_port, QN => n2401);
   registers_reg_19_10_inst : DFFR_X1 port map( D => n3409, CK => n640, RN => 
                           n6150, Q => registers_19_10_port, QN => n2400);
   registers_reg_19_9_inst : DFFR_X1 port map( D => n3408, CK => n640, RN => 
                           n6088, Q => registers_19_9_port, QN => n2399);
   registers_reg_19_8_inst : DFFR_X1 port map( D => n3407, CK => n640, RN => 
                           n6113, Q => registers_19_8_port, QN => n2398);
   registers_reg_19_7_inst : DFFR_X1 port map( D => n3406, CK => n640, RN => 
                           n6105, Q => registers_19_7_port, QN => n2397);
   registers_reg_19_6_inst : DFFR_X1 port map( D => n3405, CK => n640, RN => 
                           n6143, Q => registers_19_6_port, QN => n2396);
   registers_reg_19_5_inst : DFFR_X1 port map( D => n3404, CK => n640, RN => 
                           n6095, Q => registers_19_5_port, QN => n2395);
   registers_reg_19_4_inst : DFFR_X1 port map( D => n3403, CK => n640, RN => 
                           n6123, Q => registers_19_4_port, QN => n2394);
   registers_reg_19_3_inst : DFFR_X1 port map( D => n3402, CK => n640, RN => 
                           n6148, Q => registers_19_3_port, QN => n2393);
   registers_reg_19_2_inst : DFFR_X1 port map( D => n3401, CK => n640, RN => 
                           n6153, Q => registers_19_2_port, QN => n2392);
   registers_reg_19_1_inst : DFFR_X1 port map( D => n3400, CK => n640, RN => 
                           n6128, Q => registers_19_1_port, QN => n2391);
   registers_reg_19_0_inst : DFFR_X1 port map( D => n3399, CK => n640, RN => 
                           n6075, Q => registers_19_0_port, QN => n2389);
   registers_reg_20_31_inst : DFFR_X1 port map( D => n3398, CK => n640, RN => 
                           n6085, Q => registers_20_31_port, QN => n2948);
   registers_reg_20_30_inst : DFFR_X1 port map( D => n3397, CK => n640, RN => 
                           n6083, Q => registers_20_30_port, QN => n2947);
   registers_reg_20_29_inst : DFFR_X1 port map( D => n3396, CK => n640, RN => 
                           n6080, Q => registers_20_29_port, QN => n4204);
   registers_reg_20_28_inst : DFFR_X1 port map( D => n3395, CK => n640, RN => 
                           n6078, Q => registers_20_28_port, QN => n4147);
   registers_reg_20_27_inst : DFFR_X1 port map( D => n3394, CK => n640, RN => 
                           n6093, Q => registers_20_27_port, QN => n4128);
   registers_reg_20_26_inst : DFFR_X1 port map( D => n3393, CK => n640, RN => 
                           n6103, Q => registers_20_26_port, QN => n4185);
   registers_reg_20_25_inst : DFFR_X1 port map( D => n3392, CK => n640, RN => 
                           n6110, Q => registers_20_25_port, QN => n4109);
   registers_reg_20_24_inst : DFFR_X1 port map( D => n3391, CK => n640, RN => 
                           n6090, Q => registers_20_24_port, QN => n4090);
   registers_reg_20_23_inst : DFFR_X1 port map( D => n3390, CK => n640, RN => 
                           n6100, Q => registers_20_23_port, QN => n4071);
   registers_reg_20_22_inst : DFFR_X1 port map( D => n3389, CK => n640, RN => 
                           n6108, Q => registers_20_22_port, QN => n4052);
   registers_reg_20_21_inst : DFFR_X1 port map( D => n3388, CK => n640, RN => 
                           n6120, Q => registers_20_21_port, QN => n4033);
   registers_reg_20_20_inst : DFFR_X1 port map( D => n3387, CK => n640, RN => 
                           n6098, Q => registers_20_20_port, QN => n4014);
   registers_reg_20_19_inst : DFFR_X1 port map( D => n3386, CK => n640, RN => 
                           n6125, Q => registers_20_19_port, QN => n2946);
   registers_reg_20_18_inst : DFFR_X1 port map( D => n3385, CK => n640, RN => 
                           n6118, Q => registers_20_18_port, QN => n2945);
   registers_reg_20_17_inst : DFFR_X1 port map( D => n3384, CK => n640, RN => 
                           n6133, Q => registers_20_17_port, QN => n4166);
   registers_reg_20_16_inst : DFFR_X1 port map( D => n3383, CK => n640, RN => 
                           n6130, Q => registers_20_16_port, QN => n2944);
   registers_reg_20_15_inst : DFFR_X1 port map( D => n3382, CK => n640, RN => 
                           n6115, Q => registers_20_15_port, QN => n2943);
   registers_reg_20_14_inst : DFFR_X1 port map( D => n3381, CK => n640, RN => 
                           n6140, Q => registers_20_14_port, QN => n2942);
   registers_reg_20_13_inst : DFFR_X1 port map( D => n3380, CK => n640, RN => 
                           n6138, Q => registers_20_13_port, QN => n2941);
   registers_reg_20_12_inst : DFFR_X1 port map( D => n3379, CK => n640, RN => 
                           n6135, Q => registers_20_12_port, QN => n2940);
   registers_reg_20_11_inst : DFFR_X1 port map( D => n3378, CK => n640, RN => 
                           n6145, Q => registers_20_11_port, QN => n2939);
   registers_reg_20_10_inst : DFFR_X1 port map( D => n3377, CK => n640, RN => 
                           n6150, Q => registers_20_10_port, QN => n2938);
   registers_reg_20_9_inst : DFFR_X1 port map( D => n3376, CK => n640, RN => 
                           n6088, Q => registers_20_9_port, QN => n2937);
   registers_reg_20_8_inst : DFFR_X1 port map( D => n3375, CK => n640, RN => 
                           n6113, Q => registers_20_8_port, QN => n2949);
   registers_reg_20_7_inst : DFFR_X1 port map( D => n3374, CK => n640, RN => 
                           n6105, Q => registers_20_7_port, QN => n2936);
   registers_reg_20_6_inst : DFFR_X1 port map( D => n3373, CK => n640, RN => 
                           n6143, Q => registers_20_6_port, QN => n2935);
   registers_reg_20_5_inst : DFFR_X1 port map( D => n3372, CK => n640, RN => 
                           n6095, Q => registers_20_5_port, QN => n2934);
   registers_reg_20_4_inst : DFFR_X1 port map( D => n3371, CK => n640, RN => 
                           n6123, Q => registers_20_4_port, QN => n2933);
   registers_reg_20_3_inst : DFFR_X1 port map( D => n3370, CK => n640, RN => 
                           n6148, Q => registers_20_3_port, QN => n2932);
   registers_reg_20_2_inst : DFFR_X1 port map( D => n3369, CK => n640, RN => 
                           n6153, Q => registers_20_2_port, QN => n2931);
   registers_reg_20_1_inst : DFFR_X1 port map( D => n3368, CK => n640, RN => 
                           n6128, Q => registers_20_1_port, QN => n2930);
   registers_reg_20_0_inst : DFFR_X1 port map( D => n3367, CK => n640, RN => 
                           n6075, Q => net163843, QN => n2224);
   registers_reg_21_31_inst : DFFR_X1 port map( D => n3366, CK => n640, RN => 
                           n6085, Q => registers_21_31_port, QN => n5246);
   registers_reg_21_30_inst : DFFR_X1 port map( D => n3365, CK => n640, RN => 
                           n6083, Q => registers_21_30_port, QN => n5245);
   registers_reg_21_29_inst : DFFR_X1 port map( D => n3364, CK => n640, RN => 
                           n6080, Q => registers_21_29_port, QN => n5244);
   registers_reg_21_28_inst : DFFR_X1 port map( D => n3363, CK => n640, RN => 
                           n6078, Q => registers_21_28_port, QN => n5243);
   registers_reg_21_27_inst : DFFR_X1 port map( D => n3362, CK => n640, RN => 
                           n6093, Q => registers_21_27_port, QN => n5242);
   registers_reg_21_26_inst : DFFR_X1 port map( D => n3361, CK => n640, RN => 
                           n6103, Q => registers_21_26_port, QN => n5241);
   registers_reg_21_25_inst : DFFR_X1 port map( D => n3360, CK => n640, RN => 
                           n6110, Q => registers_21_25_port, QN => n5240);
   registers_reg_21_24_inst : DFFR_X1 port map( D => n3359, CK => n640, RN => 
                           n6090, Q => registers_21_24_port, QN => n5239);
   registers_reg_21_23_inst : DFFR_X1 port map( D => n3358, CK => n640, RN => 
                           n6100, Q => registers_21_23_port, QN => n5237);
   registers_reg_21_22_inst : DFFR_X1 port map( D => n3357, CK => n640, RN => 
                           n6108, Q => registers_21_22_port, QN => n5236);
   registers_reg_21_21_inst : DFFR_X1 port map( D => n3356, CK => n640, RN => 
                           n6120, Q => registers_21_21_port, QN => n5235);
   registers_reg_21_20_inst : DFFR_X1 port map( D => n3355, CK => n640, RN => 
                           n6098, Q => registers_21_20_port, QN => n5234);
   registers_reg_21_19_inst : DFFR_X1 port map( D => n3354, CK => n640, RN => 
                           n6125, Q => registers_21_19_port, QN => n5233);
   registers_reg_21_18_inst : DFFR_X1 port map( D => n3353, CK => n640, RN => 
                           n6118, Q => registers_21_18_port, QN => n5232);
   registers_reg_21_17_inst : DFFR_X1 port map( D => n3352, CK => n640, RN => 
                           n6133, Q => registers_21_17_port, QN => n5231);
   registers_reg_21_16_inst : DFFR_X1 port map( D => n3351, CK => n640, RN => 
                           n6130, Q => registers_21_16_port, QN => n5230);
   registers_reg_21_15_inst : DFFR_X1 port map( D => n3350, CK => n640, RN => 
                           n6115, Q => registers_21_15_port, QN => n5229);
   registers_reg_21_14_inst : DFFR_X1 port map( D => n3349, CK => n640, RN => 
                           n6140, Q => registers_21_14_port, QN => n5228);
   registers_reg_21_13_inst : DFFR_X1 port map( D => n3348, CK => n640, RN => 
                           n6138, Q => registers_21_13_port, QN => n5227);
   registers_reg_21_12_inst : DFFR_X1 port map( D => n3347, CK => n640, RN => 
                           n6135, Q => registers_21_12_port, QN => n5226);
   registers_reg_21_11_inst : DFFR_X1 port map( D => n3346, CK => n640, RN => 
                           n6145, Q => registers_21_11_port, QN => n5225);
   registers_reg_21_10_inst : DFFR_X1 port map( D => n3345, CK => n640, RN => 
                           n6150, Q => registers_21_10_port, QN => n5224);
   registers_reg_21_9_inst : DFFR_X1 port map( D => n3344, CK => n640, RN => 
                           n6088, Q => registers_21_9_port, QN => n5223);
   registers_reg_21_8_inst : DFFR_X1 port map( D => n3343, CK => n640, RN => 
                           n6113, Q => registers_21_8_port, QN => n5222);
   registers_reg_21_7_inst : DFFR_X1 port map( D => n3342, CK => n640, RN => 
                           n6105, Q => registers_21_7_port, QN => n5221);
   registers_reg_21_6_inst : DFFR_X1 port map( D => n3341, CK => n640, RN => 
                           n6143, Q => registers_21_6_port, QN => n5220);
   registers_reg_21_5_inst : DFFR_X1 port map( D => n3340, CK => n640, RN => 
                           n6095, Q => registers_21_5_port, QN => n5219);
   registers_reg_21_4_inst : DFFR_X1 port map( D => n3339, CK => n640, RN => 
                           n6123, Q => registers_21_4_port, QN => n5218);
   registers_reg_21_3_inst : DFFR_X1 port map( D => n3338, CK => n640, RN => 
                           n6148, Q => registers_21_3_port, QN => n5217);
   registers_reg_21_2_inst : DFFR_X1 port map( D => n3337, CK => n640, RN => 
                           n6153, Q => registers_21_2_port, QN => n5216);
   registers_reg_21_1_inst : DFFR_X1 port map( D => n3336, CK => n640, RN => 
                           n6128, Q => registers_21_1_port, QN => n5215);
   registers_reg_21_0_inst : DFFR_X1 port map( D => n3335, CK => n640, RN => 
                           n6075, Q => registers_21_0_port, QN => n2422);
   registers_reg_22_31_inst : DFFR_X1 port map( D => n3334, CK => n640, RN => 
                           n6085, Q => registers_22_31_port, QN => n5278);
   registers_reg_22_30_inst : DFFR_X1 port map( D => n3333, CK => n640, RN => 
                           n6083, Q => registers_22_30_port, QN => n5277);
   registers_reg_22_29_inst : DFFR_X1 port map( D => n3332, CK => n640, RN => 
                           n6080, Q => registers_22_29_port, QN => n5276);
   registers_reg_22_28_inst : DFFR_X1 port map( D => n3331, CK => n640, RN => 
                           n6078, Q => registers_22_28_port, QN => n5275);
   registers_reg_22_27_inst : DFFR_X1 port map( D => n3330, CK => n640, RN => 
                           n6093, Q => registers_22_27_port, QN => n5274);
   registers_reg_22_26_inst : DFFR_X1 port map( D => n3329, CK => n640, RN => 
                           n6103, Q => registers_22_26_port, QN => n5273);
   registers_reg_22_25_inst : DFFR_X1 port map( D => n3328, CK => n640, RN => 
                           n6110, Q => registers_22_25_port, QN => n5272);
   registers_reg_22_24_inst : DFFR_X1 port map( D => n3327, CK => n640, RN => 
                           n6090, Q => registers_22_24_port, QN => n5271);
   registers_reg_22_23_inst : DFFR_X1 port map( D => n3326, CK => n640, RN => 
                           n6100, Q => registers_22_23_port, QN => n5270);
   registers_reg_22_22_inst : DFFR_X1 port map( D => n3325, CK => n640, RN => 
                           n6108, Q => registers_22_22_port, QN => n5269);
   registers_reg_22_21_inst : DFFR_X1 port map( D => n3324, CK => n640, RN => 
                           n6120, Q => registers_22_21_port, QN => n5268);
   registers_reg_22_20_inst : DFFR_X1 port map( D => n3323, CK => n640, RN => 
                           n6098, Q => registers_22_20_port, QN => n5267);
   registers_reg_22_19_inst : DFFR_X1 port map( D => n3322, CK => n640, RN => 
                           n6125, Q => registers_22_19_port, QN => n5266);
   registers_reg_22_18_inst : DFFR_X1 port map( D => n3321, CK => n640, RN => 
                           n6118, Q => registers_22_18_port, QN => n5265);
   registers_reg_22_17_inst : DFFR_X1 port map( D => n3320, CK => n640, RN => 
                           n6133, Q => registers_22_17_port, QN => n5264);
   registers_reg_22_16_inst : DFFR_X1 port map( D => n3319, CK => n640, RN => 
                           n6131, Q => registers_22_16_port, QN => n5263);
   registers_reg_22_15_inst : DFFR_X1 port map( D => n3318, CK => n640, RN => 
                           n6115, Q => registers_22_15_port, QN => n5262);
   registers_reg_22_14_inst : DFFR_X1 port map( D => n3317, CK => n640, RN => 
                           n6141, Q => registers_22_14_port, QN => n5261);
   registers_reg_22_13_inst : DFFR_X1 port map( D => n3316, CK => n640, RN => 
                           n6138, Q => registers_22_13_port, QN => n5260);
   registers_reg_22_12_inst : DFFR_X1 port map( D => n3315, CK => n640, RN => 
                           n6136, Q => registers_22_12_port, QN => n5259);
   registers_reg_22_11_inst : DFFR_X1 port map( D => n3314, CK => n640, RN => 
                           n6146, Q => registers_22_11_port, QN => n5258);
   registers_reg_22_10_inst : DFFR_X1 port map( D => n3313, CK => n640, RN => 
                           n6151, Q => registers_22_10_port, QN => n5257);
   registers_reg_22_9_inst : DFFR_X1 port map( D => n3312, CK => n640, RN => 
                           n6088, Q => registers_22_9_port, QN => n5256);
   registers_reg_22_8_inst : DFFR_X1 port map( D => n3311, CK => n640, RN => 
                           n6113, Q => registers_22_8_port, QN => n5255);
   registers_reg_22_7_inst : DFFR_X1 port map( D => n3310, CK => n640, RN => 
                           n6105, Q => registers_22_7_port, QN => n5254);
   registers_reg_22_6_inst : DFFR_X1 port map( D => n3309, CK => n640, RN => 
                           n6143, Q => registers_22_6_port, QN => n5253);
   registers_reg_22_5_inst : DFFR_X1 port map( D => n3308, CK => n640, RN => 
                           n6095, Q => registers_22_5_port, QN => n5252);
   registers_reg_22_4_inst : DFFR_X1 port map( D => n3307, CK => n640, RN => 
                           n6123, Q => registers_22_4_port, QN => n5251);
   registers_reg_22_3_inst : DFFR_X1 port map( D => n3306, CK => n640, RN => 
                           n6148, Q => registers_22_3_port, QN => n5250);
   registers_reg_22_2_inst : DFFR_X1 port map( D => n3305, CK => n640, RN => 
                           n6153, Q => registers_22_2_port, QN => n5249);
   registers_reg_22_1_inst : DFFR_X1 port map( D => n3304, CK => n640, RN => 
                           n6128, Q => registers_22_1_port, QN => n5248);
   registers_reg_22_0_inst : DFFR_X1 port map( D => n3303, CK => n640, RN => 
                           n6075, Q => registers_22_0_port, QN => n5247);
   registers_reg_23_31_inst : DFFR_X1 port map( D => n3302, CK => n640, RN => 
                           n6086, Q => net163842, QN => n2175);
   registers_reg_23_30_inst : DFFR_X1 port map( D => n3301, CK => n640, RN => 
                           n6083, Q => net163841, QN => n2174);
   registers_reg_23_29_inst : DFFR_X1 port map( D => n3300, CK => n640, RN => 
                           n6081, Q => net163840, QN => n2189);
   registers_reg_23_28_inst : DFFR_X1 port map( D => n3299, CK => n640, RN => 
                           n6078, Q => net163839, QN => n2173);
   registers_reg_23_27_inst : DFFR_X1 port map( D => n3298, CK => n640, RN => 
                           n6093, Q => net163838, QN => n2172);
   registers_reg_23_26_inst : DFFR_X1 port map( D => n3297, CK => n640, RN => 
                           n6103, Q => net163837, QN => n2188);
   registers_reg_23_25_inst : DFFR_X1 port map( D => n3296, CK => n640, RN => 
                           n6111, Q => net163836, QN => n2171);
   registers_reg_23_24_inst : DFFR_X1 port map( D => n3295, CK => n640, RN => 
                           n6091, Q => net163835, QN => n2170);
   registers_reg_23_23_inst : DFFR_X1 port map( D => n3294, CK => n640, RN => 
                           n6101, Q => net163834, QN => n2187);
   registers_reg_23_22_inst : DFFR_X1 port map( D => n3293, CK => n640, RN => 
                           n6108, Q => net163833, QN => n2169);
   registers_reg_23_21_inst : DFFR_X1 port map( D => n3292, CK => n640, RN => 
                           n6121, Q => net163832, QN => n2168);
   registers_reg_23_20_inst : DFFR_X1 port map( D => n3291, CK => n640, RN => 
                           n6098, Q => net163831, QN => n2186);
   registers_reg_23_19_inst : DFFR_X1 port map( D => n3290, CK => n640, RN => 
                           n6126, Q => net163830, QN => n2167);
   registers_reg_23_18_inst : DFFR_X1 port map( D => n3289, CK => n640, RN => 
                           n6118, Q => net163829, QN => n2166);
   registers_reg_23_17_inst : DFFR_X1 port map( D => n3288, CK => n640, RN => 
                           n6133, Q => net163828, QN => n2185);
   registers_reg_23_16_inst : DFFR_X1 port map( D => n3287, CK => n640, RN => 
                           n6131, Q => net163827, QN => n2165);
   registers_reg_23_15_inst : DFFR_X1 port map( D => n3286, CK => n640, RN => 
                           n6116, Q => net163826, QN => n2164);
   registers_reg_23_14_inst : DFFR_X1 port map( D => n3285, CK => n640, RN => 
                           n6141, Q => net163825, QN => n2184);
   registers_reg_23_13_inst : DFFR_X1 port map( D => n3284, CK => n640, RN => 
                           n6138, Q => net163824, QN => n2163);
   registers_reg_23_12_inst : DFFR_X1 port map( D => n3283, CK => n640, RN => 
                           n6136, Q => net163823, QN => n2162);
   registers_reg_23_11_inst : DFFR_X1 port map( D => n3282, CK => n640, RN => 
                           n6146, Q => net163822, QN => n2179);
   registers_reg_23_10_inst : DFFR_X1 port map( D => n3281, CK => n640, RN => 
                           n6151, Q => net163821, QN => n2161);
   registers_reg_23_9_inst : DFFR_X1 port map( D => n3280, CK => n640, RN => 
                           n6088, Q => net163820, QN => n2160);
   registers_reg_23_8_inst : DFFR_X1 port map( D => n3279, CK => n640, RN => 
                           n6113, Q => net163819, QN => n2178);
   registers_reg_23_7_inst : DFFR_X1 port map( D => n3278, CK => n640, RN => 
                           n6106, Q => net163818, QN => n2159);
   registers_reg_23_6_inst : DFFR_X1 port map( D => n3277, CK => n640, RN => 
                           n6143, Q => net163817, QN => n2158);
   registers_reg_23_5_inst : DFFR_X1 port map( D => n3276, CK => n640, RN => 
                           n6096, Q => net163816, QN => n2177);
   registers_reg_23_4_inst : DFFR_X1 port map( D => n3275, CK => n640, RN => 
                           n6123, Q => net163815, QN => n2157);
   registers_reg_23_3_inst : DFFR_X1 port map( D => n3274, CK => n640, RN => 
                           n6148, Q => net163814, QN => n2156);
   registers_reg_23_2_inst : DFFR_X1 port map( D => n3273, CK => n640, RN => 
                           n6153, Q => net163813, QN => n2176);
   registers_reg_23_1_inst : DFFR_X1 port map( D => n3272, CK => n640, RN => 
                           n6128, Q => net163812, QN => n2155);
   registers_reg_23_0_inst : DFFR_X1 port map( D => n3271, CK => n640, RN => 
                           n6075, Q => net163811, QN => n2223);
   registers_reg_24_31_inst : DFFR_X1 port map( D => n3270, CK => n640, RN => 
                           n6086, Q => net163810, QN => n2510);
   registers_reg_24_30_inst : DFFR_X1 port map( D => n3269, CK => n640, RN => 
                           n6083, Q => net163809, QN => n2509);
   registers_reg_24_29_inst : DFFR_X1 port map( D => n3268, CK => n640, RN => 
                           n6081, Q => net163808, QN => n2522);
   registers_reg_24_28_inst : DFFR_X1 port map( D => n3267, CK => n640, RN => 
                           n6078, Q => net163807, QN => n2508);
   registers_reg_24_27_inst : DFFR_X1 port map( D => n3266, CK => n640, RN => 
                           n6093, Q => net163806, QN => n2507);
   registers_reg_24_26_inst : DFFR_X1 port map( D => n3265, CK => n640, RN => 
                           n6103, Q => net163805, QN => n2521);
   registers_reg_24_25_inst : DFFR_X1 port map( D => n3264, CK => n640, RN => 
                           n6111, Q => net163804, QN => n2506);
   registers_reg_24_24_inst : DFFR_X1 port map( D => n3263, CK => n640, RN => 
                           n6091, Q => net163803, QN => n2505);
   registers_reg_24_23_inst : DFFR_X1 port map( D => n3262, CK => n640, RN => 
                           n6101, Q => net163802, QN => n2520);
   registers_reg_24_22_inst : DFFR_X1 port map( D => n3261, CK => n640, RN => 
                           n6108, Q => net163801, QN => n2504);
   registers_reg_24_21_inst : DFFR_X1 port map( D => n3260, CK => n640, RN => 
                           n6121, Q => net163800, QN => n2503);
   registers_reg_24_20_inst : DFFR_X1 port map( D => n3259, CK => n640, RN => 
                           n6098, Q => net163799, QN => n2519);
   registers_reg_24_19_inst : DFFR_X1 port map( D => n3258, CK => n640, RN => 
                           n6126, Q => net163798, QN => n2502);
   registers_reg_24_18_inst : DFFR_X1 port map( D => n3257, CK => n640, RN => 
                           n6118, Q => net163797, QN => n2501);
   registers_reg_24_17_inst : DFFR_X1 port map( D => n3256, CK => n640, RN => 
                           n6133, Q => net163796, QN => n2518);
   registers_reg_24_16_inst : DFFR_X1 port map( D => n3255, CK => n640, RN => 
                           n6131, Q => net163795, QN => n2500);
   registers_reg_24_15_inst : DFFR_X1 port map( D => n3254, CK => n640, RN => 
                           n6116, Q => net163794, QN => n2499);
   registers_reg_24_14_inst : DFFR_X1 port map( D => n3253, CK => n640, RN => 
                           n6141, Q => net163793, QN => n2517);
   registers_reg_24_13_inst : DFFR_X1 port map( D => n3252, CK => n640, RN => 
                           n6138, Q => net163792, QN => n2498);
   registers_reg_24_12_inst : DFFR_X1 port map( D => n3251, CK => n640, RN => 
                           n6136, Q => net163791, QN => n2497);
   registers_reg_24_11_inst : DFFR_X1 port map( D => n3250, CK => n640, RN => 
                           n6146, Q => net163790, QN => n2516);
   registers_reg_24_10_inst : DFFR_X1 port map( D => n3249, CK => n640, RN => 
                           n6151, Q => net163789, QN => n2496);
   registers_reg_24_9_inst : DFFR_X1 port map( D => n3248, CK => n640, RN => 
                           n6088, Q => net163788, QN => n2495);
   registers_reg_24_8_inst : DFFR_X1 port map( D => n3247, CK => n640, RN => 
                           n6113, Q => net163787, QN => n2515);
   registers_reg_24_7_inst : DFFR_X1 port map( D => n3246, CK => n640, RN => 
                           n6106, Q => net163786, QN => n2494);
   registers_reg_24_6_inst : DFFR_X1 port map( D => n3245, CK => n640, RN => 
                           n6143, Q => net163785, QN => n2491);
   registers_reg_24_5_inst : DFFR_X1 port map( D => n3244, CK => n640, RN => 
                           n6096, Q => net163784, QN => n2514);
   registers_reg_24_4_inst : DFFR_X1 port map( D => n3243, CK => n640, RN => 
                           n6123, Q => net163783, QN => n2490);
   registers_reg_24_3_inst : DFFR_X1 port map( D => n3242, CK => n640, RN => 
                           n6148, Q => net163782, QN => n2489);
   registers_reg_24_2_inst : DFFR_X1 port map( D => n3241, CK => n640, RN => 
                           n6153, Q => net163781, QN => n2513);
   registers_reg_24_1_inst : DFFR_X1 port map( D => n3240, CK => n640, RN => 
                           n6128, Q => net163780, QN => n2488);
   registers_reg_24_0_inst : DFFR_X1 port map( D => n3239, CK => n640, RN => 
                           n6075, Q => net163779, QN => n2512);
   registers_reg_25_31_inst : DFFR_X1 port map( D => n3238, CK => n640, RN => 
                           n6086, Q => registers_25_31_port, QN => n2587);
   registers_reg_25_30_inst : DFFR_X1 port map( D => n3237, CK => n640, RN => 
                           n6083, Q => registers_25_30_port, QN => n2586);
   registers_reg_25_29_inst : DFFR_X1 port map( D => n3236, CK => n640, RN => 
                           n6081, Q => registers_25_29_port, QN => n2585);
   registers_reg_25_28_inst : DFFR_X1 port map( D => n3235, CK => n640, RN => 
                           n6078, Q => registers_25_28_port, QN => n2584);
   registers_reg_25_27_inst : DFFR_X1 port map( D => n3234, CK => n640, RN => 
                           n6093, Q => registers_25_27_port, QN => n2583);
   registers_reg_25_26_inst : DFFR_X1 port map( D => n3233, CK => n640, RN => 
                           n6103, Q => registers_25_26_port, QN => n2582);
   registers_reg_25_25_inst : DFFR_X1 port map( D => n3232, CK => n640, RN => 
                           n6111, Q => registers_25_25_port, QN => n2581);
   registers_reg_25_24_inst : DFFR_X1 port map( D => n3231, CK => n640, RN => 
                           n6091, Q => registers_25_24_port, QN => n2580);
   registers_reg_25_23_inst : DFFR_X1 port map( D => n3230, CK => n640, RN => 
                           n6101, Q => registers_25_23_port, QN => n2579);
   registers_reg_25_22_inst : DFFR_X1 port map( D => n3229, CK => n640, RN => 
                           n6108, Q => registers_25_22_port, QN => n2578);
   registers_reg_25_21_inst : DFFR_X1 port map( D => n3228, CK => n640, RN => 
                           n6121, Q => registers_25_21_port, QN => n2577);
   registers_reg_25_20_inst : DFFR_X1 port map( D => n3227, CK => n640, RN => 
                           n6098, Q => registers_25_20_port, QN => n2576);
   registers_reg_25_19_inst : DFFR_X1 port map( D => n3226, CK => n640, RN => 
                           n6126, Q => registers_25_19_port, QN => n2575);
   registers_reg_25_18_inst : DFFR_X1 port map( D => n3225, CK => n640, RN => 
                           n6118, Q => registers_25_18_port, QN => n2574);
   registers_reg_25_17_inst : DFFR_X1 port map( D => n3224, CK => n640, RN => 
                           n6133, Q => registers_25_17_port, QN => n2573);
   registers_reg_25_16_inst : DFFR_X1 port map( D => n3223, CK => n640, RN => 
                           n6131, Q => registers_25_16_port, QN => n2572);
   registers_reg_25_15_inst : DFFR_X1 port map( D => n3222, CK => n640, RN => 
                           n6116, Q => registers_25_15_port, QN => n2571);
   registers_reg_25_14_inst : DFFR_X1 port map( D => n3221, CK => n640, RN => 
                           n6141, Q => registers_25_14_port, QN => n2570);
   registers_reg_25_13_inst : DFFR_X1 port map( D => n3220, CK => n640, RN => 
                           n6138, Q => registers_25_13_port, QN => n2569);
   registers_reg_25_12_inst : DFFR_X1 port map( D => n3219, CK => n640, RN => 
                           n6136, Q => registers_25_12_port, QN => n2568);
   registers_reg_25_11_inst : DFFR_X1 port map( D => n3218, CK => n640, RN => 
                           n6146, Q => registers_25_11_port, QN => n2567);
   registers_reg_25_10_inst : DFFR_X1 port map( D => n3217, CK => n640, RN => 
                           n6151, Q => registers_25_10_port, QN => n2566);
   registers_reg_25_9_inst : DFFR_X1 port map( D => n3216, CK => n640, RN => 
                           n6088, Q => registers_25_9_port, QN => n2565);
   registers_reg_25_8_inst : DFFR_X1 port map( D => n3215, CK => n640, RN => 
                           n6113, Q => registers_25_8_port, QN => n2564);
   registers_reg_25_7_inst : DFFR_X1 port map( D => n3214, CK => n640, RN => 
                           n6106, Q => registers_25_7_port, QN => n2563);
   registers_reg_25_6_inst : DFFR_X1 port map( D => n3213, CK => n640, RN => 
                           n6143, Q => registers_25_6_port, QN => n2562);
   registers_reg_25_5_inst : DFFR_X1 port map( D => n3212, CK => n640, RN => 
                           n6096, Q => registers_25_5_port, QN => n2560);
   registers_reg_25_4_inst : DFFR_X1 port map( D => n3211, CK => n640, RN => 
                           n6123, Q => registers_25_4_port, QN => n2559);
   registers_reg_25_3_inst : DFFR_X1 port map( D => n3210, CK => n640, RN => 
                           n6148, Q => registers_25_3_port, QN => n2558);
   registers_reg_25_2_inst : DFFR_X1 port map( D => n3209, CK => n640, RN => 
                           n6153, Q => registers_25_2_port, QN => n2557);
   registers_reg_25_1_inst : DFFR_X1 port map( D => n3208, CK => n640, RN => 
                           n6128, Q => registers_25_1_port, QN => n2556);
   registers_reg_25_0_inst : DFFR_X1 port map( D => n3207, CK => n640, RN => 
                           n6076, Q => registers_25_0_port, QN => n2555);
   registers_reg_26_31_inst : DFFR_X1 port map( D => n3206, CK => n640, RN => 
                           n6086, Q => registers_26_31_port, QN => n2487);
   registers_reg_26_30_inst : DFFR_X1 port map( D => n3205, CK => n640, RN => 
                           n6083, Q => registers_26_30_port, QN => n2486);
   registers_reg_26_29_inst : DFFR_X1 port map( D => n3204, CK => n640, RN => 
                           n6081, Q => registers_26_29_port, QN => n2485);
   registers_reg_26_28_inst : DFFR_X1 port map( D => n3203, CK => n640, RN => 
                           n6078, Q => registers_26_28_port, QN => n2484);
   registers_reg_26_27_inst : DFFR_X1 port map( D => n3202, CK => n640, RN => 
                           n6093, Q => registers_26_27_port, QN => n2483);
   registers_reg_26_26_inst : DFFR_X1 port map( D => n3201, CK => n640, RN => 
                           n6103, Q => registers_26_26_port, QN => n2482);
   registers_reg_26_25_inst : DFFR_X1 port map( D => n3200, CK => n640, RN => 
                           n6111, Q => registers_26_25_port, QN => n2481);
   registers_reg_26_24_inst : DFFR_X1 port map( D => n3199, CK => n640, RN => 
                           n6091, Q => registers_26_24_port, QN => n2480);
   registers_reg_26_23_inst : DFFR_X1 port map( D => n3198, CK => n640, RN => 
                           n6101, Q => registers_26_23_port, QN => n2478);
   registers_reg_26_22_inst : DFFR_X1 port map( D => n3197, CK => n640, RN => 
                           n6108, Q => registers_26_22_port, QN => n2477);
   registers_reg_26_21_inst : DFFR_X1 port map( D => n3196, CK => n640, RN => 
                           n6121, Q => registers_26_21_port, QN => n2476);
   registers_reg_26_20_inst : DFFR_X1 port map( D => n3195, CK => n640, RN => 
                           n6098, Q => registers_26_20_port, QN => n2475);
   registers_reg_26_19_inst : DFFR_X1 port map( D => n3194, CK => n640, RN => 
                           n6126, Q => registers_26_19_port, QN => n2474);
   registers_reg_26_18_inst : DFFR_X1 port map( D => n3193, CK => n640, RN => 
                           n6118, Q => registers_26_18_port, QN => n2473);
   registers_reg_26_17_inst : DFFR_X1 port map( D => n3192, CK => n640, RN => 
                           n6133, Q => registers_26_17_port, QN => n2472);
   registers_reg_26_16_inst : DFFR_X1 port map( D => n3191, CK => n640, RN => 
                           n6131, Q => registers_26_16_port, QN => n2471);
   registers_reg_26_15_inst : DFFR_X1 port map( D => n3190, CK => n640, RN => 
                           n6116, Q => registers_26_15_port, QN => n2470);
   registers_reg_26_14_inst : DFFR_X1 port map( D => n3189, CK => n640, RN => 
                           n6141, Q => registers_26_14_port, QN => n2469);
   registers_reg_26_13_inst : DFFR_X1 port map( D => n3188, CK => n640, RN => 
                           n6138, Q => registers_26_13_port, QN => n2468);
   registers_reg_26_12_inst : DFFR_X1 port map( D => n3187, CK => n640, RN => 
                           n6136, Q => registers_26_12_port, QN => n2467);
   registers_reg_26_11_inst : DFFR_X1 port map( D => n3186, CK => n640, RN => 
                           n6146, Q => registers_26_11_port, QN => n2466);
   registers_reg_26_10_inst : DFFR_X1 port map( D => n3185, CK => n640, RN => 
                           n6151, Q => registers_26_10_port, QN => n2465);
   registers_reg_26_9_inst : DFFR_X1 port map( D => n3184, CK => n640, RN => 
                           n6088, Q => registers_26_9_port, QN => n2464);
   registers_reg_26_8_inst : DFFR_X1 port map( D => n3183, CK => n640, RN => 
                           n6113, Q => registers_26_8_port, QN => n2463);
   registers_reg_26_7_inst : DFFR_X1 port map( D => n3182, CK => n640, RN => 
                           n6106, Q => registers_26_7_port, QN => n2462);
   registers_reg_26_6_inst : DFFR_X1 port map( D => n3181, CK => n640, RN => 
                           n6143, Q => registers_26_6_port, QN => n2461);
   registers_reg_26_5_inst : DFFR_X1 port map( D => n3180, CK => n640, RN => 
                           n6096, Q => registers_26_5_port, QN => n2460);
   registers_reg_26_4_inst : DFFR_X1 port map( D => n3179, CK => n640, RN => 
                           n6123, Q => registers_26_4_port, QN => n2459);
   registers_reg_26_3_inst : DFFR_X1 port map( D => n3178, CK => n640, RN => 
                           n6148, Q => registers_26_3_port, QN => n2457);
   registers_reg_26_2_inst : DFFR_X1 port map( D => n3177, CK => n640, RN => 
                           n6153, Q => registers_26_2_port, QN => n2456);
   registers_reg_26_1_inst : DFFR_X1 port map( D => n3176, CK => n640, RN => 
                           n6128, Q => registers_26_1_port, QN => n2455);
   registers_reg_26_0_inst : DFFR_X1 port map( D => n3175, CK => n640, RN => 
                           n6076, Q => registers_26_0_port, QN => n5279);
   registers_reg_27_31_inst : DFFR_X1 port map( D => n3174, CK => n640, RN => 
                           n6086, Q => registers_27_31_port, QN => n2373);
   registers_reg_27_30_inst : DFFR_X1 port map( D => n3173, CK => n640, RN => 
                           n6083, Q => registers_27_30_port, QN => n2372);
   registers_reg_27_29_inst : DFFR_X1 port map( D => n3172, CK => n640, RN => 
                           n6081, Q => registers_27_29_port, QN => n2385);
   registers_reg_27_28_inst : DFFR_X1 port map( D => n3171, CK => n640, RN => 
                           n6078, Q => registers_27_28_port, QN => n2382);
   registers_reg_27_27_inst : DFFR_X1 port map( D => n3170, CK => n640, RN => 
                           n6093, Q => registers_27_27_port, QN => n2381);
   registers_reg_27_26_inst : DFFR_X1 port map( D => n3169, CK => n640, RN => 
                           n6103, Q => registers_27_26_port, QN => n2384);
   registers_reg_27_25_inst : DFFR_X1 port map( D => n3168, CK => n640, RN => 
                           n6111, Q => registers_27_25_port, QN => n2380);
   registers_reg_27_24_inst : DFFR_X1 port map( D => n3167, CK => n640, RN => 
                           n6091, Q => registers_27_24_port, QN => n2379);
   registers_reg_27_23_inst : DFFR_X1 port map( D => n3166, CK => n640, RN => 
                           n6101, Q => registers_27_23_port, QN => n2378);
   registers_reg_27_22_inst : DFFR_X1 port map( D => n3165, CK => n640, RN => 
                           n6108, Q => registers_27_22_port, QN => n2377);
   registers_reg_27_21_inst : DFFR_X1 port map( D => n3164, CK => n640, RN => 
                           n6121, Q => registers_27_21_port, QN => n2376);
   registers_reg_27_20_inst : DFFR_X1 port map( D => n3163, CK => n640, RN => 
                           n6098, Q => registers_27_20_port, QN => n2375);
   registers_reg_27_19_inst : DFFR_X1 port map( D => n3162, CK => n640, RN => 
                           n6126, Q => registers_27_19_port, QN => n2371);
   registers_reg_27_18_inst : DFFR_X1 port map( D => n3161, CK => n640, RN => 
                           n6118, Q => registers_27_18_port, QN => n2370);
   registers_reg_27_17_inst : DFFR_X1 port map( D => n3160, CK => n640, RN => 
                           n6133, Q => registers_27_17_port, QN => n2383);
   registers_reg_27_16_inst : DFFR_X1 port map( D => n3159, CK => n640, RN => 
                           n6131, Q => registers_27_16_port, QN => n2369);
   registers_reg_27_15_inst : DFFR_X1 port map( D => n3158, CK => n640, RN => 
                           n6116, Q => registers_27_15_port, QN => n2368);
   registers_reg_27_14_inst : DFFR_X1 port map( D => n3157, CK => n640, RN => 
                           n6141, Q => registers_27_14_port, QN => n2367);
   registers_reg_27_13_inst : DFFR_X1 port map( D => n3156, CK => n640, RN => 
                           n6138, Q => registers_27_13_port, QN => n2366);
   registers_reg_27_12_inst : DFFR_X1 port map( D => n3155, CK => n640, RN => 
                           n6136, Q => registers_27_12_port, QN => n2365);
   registers_reg_27_11_inst : DFFR_X1 port map( D => n3154, CK => n640, RN => 
                           n6146, Q => registers_27_11_port, QN => n2364);
   registers_reg_27_10_inst : DFFR_X1 port map( D => n3153, CK => n640, RN => 
                           n6151, Q => registers_27_10_port, QN => n2363);
   registers_reg_27_9_inst : DFFR_X1 port map( D => n3152, CK => n640, RN => 
                           n6088, Q => registers_27_9_port, QN => n2362);
   registers_reg_27_8_inst : DFFR_X1 port map( D => n3151, CK => n640, RN => 
                           n6113, Q => registers_27_8_port, QN => n2374);
   registers_reg_27_7_inst : DFFR_X1 port map( D => n3150, CK => n640, RN => 
                           n6106, Q => registers_27_7_port, QN => n2361);
   registers_reg_27_6_inst : DFFR_X1 port map( D => n3149, CK => n640, RN => 
                           n6143, Q => registers_27_6_port, QN => n2360);
   registers_reg_27_5_inst : DFFR_X1 port map( D => n3148, CK => n640, RN => 
                           n6096, Q => registers_27_5_port, QN => n2359);
   registers_reg_27_4_inst : DFFR_X1 port map( D => n3147, CK => n640, RN => 
                           n6123, Q => registers_27_4_port, QN => n2358);
   registers_reg_27_3_inst : DFFR_X1 port map( D => n3146, CK => n640, RN => 
                           n6148, Q => registers_27_3_port, QN => n2357);
   registers_reg_27_2_inst : DFFR_X1 port map( D => n3145, CK => n640, RN => 
                           n6153, Q => registers_27_2_port, QN => n2354);
   registers_reg_27_1_inst : DFFR_X1 port map( D => n3144, CK => n640, RN => 
                           n6128, Q => registers_27_1_port, QN => n2353);
   registers_reg_27_0_inst : DFFR_X1 port map( D => n3143, CK => n640, RN => 
                           n6076, Q => net163778, QN => n2116);
   registers_reg_28_31_inst : DFFR_X1 port map( D => n3142, CK => n640, RN => 
                           n6086, Q => registers_28_31_port, QN => n2647);
   registers_reg_28_30_inst : DFFR_X1 port map( D => n3141, CK => n640, RN => 
                           n6083, Q => registers_28_30_port, QN => n2646);
   registers_reg_28_29_inst : DFFR_X1 port map( D => n3140, CK => n640, RN => 
                           n6081, Q => registers_28_29_port, QN => n2645);
   registers_reg_28_28_inst : DFFR_X1 port map( D => n3139, CK => n640, RN => 
                           n6078, Q => registers_28_28_port, QN => n2644);
   registers_reg_28_27_inst : DFFR_X1 port map( D => n3138, CK => n640, RN => 
                           n6093, Q => registers_28_27_port, QN => n2643);
   registers_reg_28_26_inst : DFFR_X1 port map( D => n3137, CK => n640, RN => 
                           n6103, Q => registers_28_26_port, QN => n2642);
   registers_reg_28_25_inst : DFFR_X1 port map( D => n3136, CK => n640, RN => 
                           n6111, Q => registers_28_25_port, QN => n2641);
   registers_reg_28_24_inst : DFFR_X1 port map( D => n3135, CK => n640, RN => 
                           n6091, Q => registers_28_24_port, QN => n2640);
   registers_reg_28_23_inst : DFFR_X1 port map( D => n3134, CK => n640, RN => 
                           n6101, Q => registers_28_23_port, QN => n2639);
   registers_reg_28_22_inst : DFFR_X1 port map( D => n3133, CK => n640, RN => 
                           n6108, Q => registers_28_22_port, QN => n2638);
   registers_reg_28_21_inst : DFFR_X1 port map( D => n3132, CK => n640, RN => 
                           n6121, Q => registers_28_21_port, QN => n2637);
   registers_reg_28_20_inst : DFFR_X1 port map( D => n3131, CK => n640, RN => 
                           n6098, Q => registers_28_20_port, QN => n2636);
   registers_reg_28_19_inst : DFFR_X1 port map( D => n3130, CK => n640, RN => 
                           n6126, Q => registers_28_19_port, QN => n2635);
   registers_reg_28_18_inst : DFFR_X1 port map( D => n3129, CK => n640, RN => 
                           n6118, Q => registers_28_18_port, QN => n2634);
   registers_reg_28_17_inst : DFFR_X1 port map( D => n3128, CK => n640, RN => 
                           n6134, Q => registers_28_17_port, QN => n2633);
   registers_reg_28_16_inst : DFFR_X1 port map( D => n3127, CK => n640, RN => 
                           n6131, Q => registers_28_16_port, QN => n2632);
   registers_reg_28_15_inst : DFFR_X1 port map( D => n3126, CK => n640, RN => 
                           n6116, Q => registers_28_15_port, QN => n2631);
   registers_reg_28_14_inst : DFFR_X1 port map( D => n3125, CK => n640, RN => 
                           n6141, Q => registers_28_14_port, QN => n2628);
   registers_reg_28_13_inst : DFFR_X1 port map( D => n3124, CK => n640, RN => 
                           n6139, Q => registers_28_13_port, QN => n2627);
   registers_reg_28_12_inst : DFFR_X1 port map( D => n3123, CK => n640, RN => 
                           n6136, Q => registers_28_12_port, QN => n2626);
   registers_reg_28_11_inst : DFFR_X1 port map( D => n3122, CK => n640, RN => 
                           n6146, Q => registers_28_11_port, QN => n2625);
   registers_reg_28_10_inst : DFFR_X1 port map( D => n3121, CK => n640, RN => 
                           n6151, Q => registers_28_10_port, QN => n2624);
   registers_reg_28_9_inst : DFFR_X1 port map( D => n3120, CK => n640, RN => 
                           n6088, Q => registers_28_9_port, QN => n2623);
   registers_reg_28_8_inst : DFFR_X1 port map( D => n3119, CK => n640, RN => 
                           n6113, Q => registers_28_8_port, QN => n2622);
   registers_reg_28_7_inst : DFFR_X1 port map( D => n3118, CK => n640, RN => 
                           n6106, Q => registers_28_7_port, QN => n2621);
   registers_reg_28_6_inst : DFFR_X1 port map( D => n3117, CK => n640, RN => 
                           n6144, Q => registers_28_6_port, QN => n2620);
   registers_reg_28_5_inst : DFFR_X1 port map( D => n3116, CK => n640, RN => 
                           n6096, Q => registers_28_5_port, QN => n2619);
   registers_reg_28_4_inst : DFFR_X1 port map( D => n3115, CK => n640, RN => 
                           n6123, Q => registers_28_4_port, QN => n2618);
   registers_reg_28_3_inst : DFFR_X1 port map( D => n3114, CK => n640, RN => 
                           n6149, Q => registers_28_3_port, QN => n2617);
   registers_reg_28_2_inst : DFFR_X1 port map( D => n3113, CK => n640, RN => 
                           n6154, Q => registers_28_2_port, QN => n2616);
   registers_reg_28_1_inst : DFFR_X1 port map( D => n3112, CK => n640, RN => 
                           n6128, Q => registers_28_1_port, QN => n2615);
   registers_reg_28_0_inst : DFFR_X1 port map( D => n3111, CK => n640, RN => 
                           n6076, Q => registers_28_0_port, QN => n2614);
   registers_reg_29_31_inst : DFFR_X1 port map( D => n3110, CK => n640, RN => 
                           n6086, Q => registers_29_31_port, QN => n2921);
   registers_reg_29_30_inst : DFFR_X1 port map( D => n3109, CK => n640, RN => 
                           n6084, Q => registers_29_30_port, QN => n2920);
   registers_reg_29_29_inst : DFFR_X1 port map( D => n3108, CK => n640, RN => 
                           n6081, Q => registers_29_29_port, QN => n2919);
   registers_reg_29_28_inst : DFFR_X1 port map( D => n3107, CK => n640, RN => 
                           n6079, Q => registers_29_28_port, QN => n2908);
   registers_reg_29_27_inst : DFFR_X1 port map( D => n3106, CK => n640, RN => 
                           n6094, Q => registers_29_27_port, QN => n2889);
   registers_reg_29_26_inst : DFFR_X1 port map( D => n3105, CK => n640, RN => 
                           n6104, Q => registers_29_26_port, QN => n2870);
   registers_reg_29_25_inst : DFFR_X1 port map( D => n3104, CK => n640, RN => 
                           n6111, Q => registers_29_25_port, QN => n2851);
   registers_reg_29_24_inst : DFFR_X1 port map( D => n3103, CK => n640, RN => 
                           n6091, Q => registers_29_24_port, QN => n2832);
   registers_reg_29_23_inst : DFFR_X1 port map( D => n3102, CK => n640, RN => 
                           n6101, Q => registers_29_23_port, QN => n2679);
   registers_reg_29_22_inst : DFFR_X1 port map( D => n3101, CK => n640, RN => 
                           n6109, Q => registers_29_22_port, QN => n2678);
   registers_reg_29_21_inst : DFFR_X1 port map( D => n3100, CK => n640, RN => 
                           n6121, Q => registers_29_21_port, QN => n2677);
   registers_reg_29_20_inst : DFFR_X1 port map( D => n3099, CK => n640, RN => 
                           n6099, Q => registers_29_20_port, QN => n2676);
   registers_reg_29_19_inst : DFFR_X1 port map( D => n3098, CK => n640, RN => 
                           n6126, Q => registers_29_19_port, QN => n2675);
   registers_reg_29_18_inst : DFFR_X1 port map( D => n3097, CK => n640, RN => 
                           n6119, Q => registers_29_18_port, QN => n2674);
   registers_reg_29_17_inst : DFFR_X1 port map( D => n3096, CK => n640, RN => 
                           n6134, Q => registers_29_17_port, QN => n2673);
   registers_reg_29_16_inst : DFFR_X1 port map( D => n3095, CK => n640, RN => 
                           n6131, Q => registers_29_16_port, QN => n2672);
   registers_reg_29_15_inst : DFFR_X1 port map( D => n3094, CK => n640, RN => 
                           n6116, Q => registers_29_15_port, QN => n2671);
   registers_reg_29_14_inst : DFFR_X1 port map( D => n3093, CK => n640, RN => 
                           n6141, Q => registers_29_14_port, QN => n2670);
   registers_reg_29_13_inst : DFFR_X1 port map( D => n3092, CK => n640, RN => 
                           n6139, Q => registers_29_13_port, QN => n2669);
   registers_reg_29_12_inst : DFFR_X1 port map( D => n3091, CK => n640, RN => 
                           n6136, Q => registers_29_12_port, QN => n2668);
   registers_reg_29_11_inst : DFFR_X1 port map( D => n3090, CK => n640, RN => 
                           n6146, Q => registers_29_11_port, QN => n2667);
   registers_reg_29_10_inst : DFFR_X1 port map( D => n3089, CK => n640, RN => 
                           n6151, Q => registers_29_10_port, QN => n2666);
   registers_reg_29_9_inst : DFFR_X1 port map( D => n3088, CK => n640, RN => 
                           n6089, Q => registers_29_9_port, QN => n2663);
   registers_reg_29_8_inst : DFFR_X1 port map( D => n3087, CK => n640, RN => 
                           n6114, Q => registers_29_8_port, QN => n2662);
   registers_reg_29_7_inst : DFFR_X1 port map( D => n3086, CK => n640, RN => 
                           n6106, Q => registers_29_7_port, QN => n2661);
   registers_reg_29_6_inst : DFFR_X1 port map( D => n3085, CK => n640, RN => 
                           n6144, Q => registers_29_6_port, QN => n2660);
   registers_reg_29_5_inst : DFFR_X1 port map( D => n3084, CK => n640, RN => 
                           n6096, Q => registers_29_5_port, QN => n2659);
   registers_reg_29_4_inst : DFFR_X1 port map( D => n3083, CK => n640, RN => 
                           n6124, Q => registers_29_4_port, QN => n2658);
   registers_reg_29_3_inst : DFFR_X1 port map( D => n3082, CK => n640, RN => 
                           n6149, Q => registers_29_3_port, QN => n2657);
   registers_reg_29_2_inst : DFFR_X1 port map( D => n3081, CK => n640, RN => 
                           n6154, Q => registers_29_2_port, QN => n2656);
   registers_reg_29_1_inst : DFFR_X1 port map( D => n3080, CK => n640, RN => 
                           n6129, Q => registers_29_1_port, QN => n2655);
   registers_reg_29_0_inst : DFFR_X1 port map( D => n3079, CK => n640, RN => 
                           n6076, Q => registers_29_0_port, QN => n2654);
   registers_reg_30_31_inst : DFFR_X1 port map( D => n3078, CK => n640, RN => 
                           n6086, Q => registers_30_31_port, QN => n5298);
   registers_reg_30_30_inst : DFFR_X1 port map( D => n3077, CK => n640, RN => 
                           n6084, Q => registers_30_30_port, QN => n5297);
   registers_reg_30_29_inst : DFFR_X1 port map( D => n3076, CK => n640, RN => 
                           n6081, Q => registers_30_29_port, QN => n5310);
   registers_reg_30_28_inst : DFFR_X1 port map( D => n3075, CK => n640, RN => 
                           n6079, Q => registers_30_28_port, QN => n5307);
   registers_reg_30_27_inst : DFFR_X1 port map( D => n3074, CK => n640, RN => 
                           n6094, Q => registers_30_27_port, QN => n5306);
   registers_reg_30_26_inst : DFFR_X1 port map( D => n3073, CK => n640, RN => 
                           n6104, Q => registers_30_26_port, QN => n5309);
   registers_reg_30_25_inst : DFFR_X1 port map( D => n3072, CK => n640, RN => 
                           n6111, Q => registers_30_25_port, QN => n5305);
   registers_reg_30_24_inst : DFFR_X1 port map( D => n3071, CK => n640, RN => 
                           n6091, Q => registers_30_24_port, QN => n5304);
   registers_reg_30_23_inst : DFFR_X1 port map( D => n3070, CK => n640, RN => 
                           n6101, Q => registers_30_23_port, QN => n5303);
   registers_reg_30_22_inst : DFFR_X1 port map( D => n3069, CK => n640, RN => 
                           n6109, Q => registers_30_22_port, QN => n5302);
   registers_reg_30_21_inst : DFFR_X1 port map( D => n3068, CK => n640, RN => 
                           n6121, Q => registers_30_21_port, QN => n5301);
   registers_reg_30_20_inst : DFFR_X1 port map( D => n3067, CK => n640, RN => 
                           n6099, Q => registers_30_20_port, QN => n5300);
   registers_reg_30_19_inst : DFFR_X1 port map( D => n3066, CK => n640, RN => 
                           n6126, Q => registers_30_19_port, QN => n5296);
   registers_reg_30_18_inst : DFFR_X1 port map( D => n3065, CK => n640, RN => 
                           n6119, Q => registers_30_18_port, QN => n5295);
   registers_reg_30_17_inst : DFFR_X1 port map( D => n3064, CK => n640, RN => 
                           n6134, Q => registers_30_17_port, QN => n5308);
   registers_reg_30_16_inst : DFFR_X1 port map( D => n3063, CK => n640, RN => 
                           n6131, Q => registers_30_16_port, QN => n5294);
   registers_reg_30_15_inst : DFFR_X1 port map( D => n3062, CK => n640, RN => 
                           n6116, Q => registers_30_15_port, QN => n5293);
   registers_reg_30_14_inst : DFFR_X1 port map( D => n3061, CK => n640, RN => 
                           n6141, Q => registers_30_14_port, QN => n5292);
   registers_reg_30_13_inst : DFFR_X1 port map( D => n3060, CK => n640, RN => 
                           n6139, Q => registers_30_13_port, QN => n5291);
   registers_reg_30_12_inst : DFFR_X1 port map( D => n3059, CK => n640, RN => 
                           n6136, Q => registers_30_12_port, QN => n5290);
   registers_reg_30_11_inst : DFFR_X1 port map( D => n3058, CK => n640, RN => 
                           n6146, Q => registers_30_11_port, QN => n5289);
   registers_reg_30_10_inst : DFFR_X1 port map( D => n3057, CK => n640, RN => 
                           n6151, Q => registers_30_10_port, QN => n5288);
   registers_reg_30_9_inst : DFFR_X1 port map( D => n3056, CK => n640, RN => 
                           n6089, Q => registers_30_9_port, QN => n5287);
   registers_reg_30_8_inst : DFFR_X1 port map( D => n3055, CK => n640, RN => 
                           n6114, Q => registers_30_8_port, QN => n5299);
   registers_reg_30_7_inst : DFFR_X1 port map( D => n3054, CK => n640, RN => 
                           n6106, Q => registers_30_7_port, QN => n5286);
   registers_reg_30_6_inst : DFFR_X1 port map( D => n3053, CK => n640, RN => 
                           n6144, Q => registers_30_6_port, QN => n5285);
   registers_reg_30_5_inst : DFFR_X1 port map( D => n3052, CK => n640, RN => 
                           n6096, Q => registers_30_5_port, QN => n5284);
   registers_reg_30_4_inst : DFFR_X1 port map( D => n3051, CK => n640, RN => 
                           n6124, Q => registers_30_4_port, QN => n5283);
   registers_reg_30_3_inst : DFFR_X1 port map( D => n3050, CK => n640, RN => 
                           n6149, Q => registers_30_3_port, QN => n5282);
   registers_reg_30_2_inst : DFFR_X1 port map( D => n3049, CK => n640, RN => 
                           n6154, Q => registers_30_2_port, QN => n5281);
   registers_reg_30_1_inst : DFFR_X1 port map( D => n3048, CK => n640, RN => 
                           n6129, Q => registers_30_1_port, QN => n5280);
   registers_reg_30_0_inst : DFFR_X1 port map( D => n3047, CK => n640, RN => 
                           n6076, Q => registers_30_0_port, QN => n5312);
   registers_reg_31_31_inst : DFFR_X1 port map( D => n3046, CK => n640, RN => 
                           n6156, Q => net108162, QN => n5313);
   d_out2_reg_31_inst : DFF_X1 port map( D => n3045, CK => n640, Q => 
                           d_out2_31_port, QN => net108161);
   registers_reg_31_30_inst : DFFR_X1 port map( D => n3044, CK => n640, RN => 
                           n6156, Q => registers_31_30_port, QN => n5344);
   d_out2_reg_30_inst : DFF_X1 port map( D => n3043, CK => n640, Q => 
                           d_out2_30_port, QN => net163777);
   registers_reg_31_29_inst : DFFR_X1 port map( D => n3042, CK => n640, RN => 
                           n6156, Q => registers_31_29_port, QN => n5343);
   d_out2_reg_29_inst : DFF_X1 port map( D => n3041, CK => n640, Q => 
                           d_out2_29_port, QN => net163776);
   registers_reg_31_28_inst : DFFR_X1 port map( D => n3040, CK => n640, RN => 
                           n6076, Q => registers_31_28_port, QN => n5342);
   d_out2_reg_28_inst : DFF_X1 port map( D => n3039, CK => n640, Q => 
                           d_out2_28_port, QN => net163775);
   registers_reg_31_27_inst : DFFR_X1 port map( D => n3038, CK => n640, RN => 
                           n6156, Q => registers_31_27_port, QN => n5341);
   d_out2_reg_27_inst : DFF_X1 port map( D => n3037, CK => n640, Q => 
                           d_out2_27_port, QN => net163774);
   registers_reg_31_26_inst : DFFR_X1 port map( D => n3036, CK => n640, RN => 
                           n6156, Q => registers_31_26_port, QN => n5340);
   d_out2_reg_26_inst : DFF_X1 port map( D => n3035, CK => n640, Q => 
                           d_out2_26_port, QN => net163773);
   registers_reg_31_25_inst : DFFR_X1 port map( D => n3034, CK => n640, RN => 
                           n6156, Q => registers_31_25_port, QN => n5339);
   d_out2_reg_25_inst : DFF_X1 port map( D => n3033, CK => n640, Q => 
                           d_out2_25_port, QN => net163772);
   registers_reg_31_24_inst : DFFR_X1 port map( D => n3032, CK => n640, RN => 
                           n6156, Q => registers_31_24_port, QN => n5338);
   d_out2_reg_24_inst : DFF_X1 port map( D => n3031, CK => n640, Q => 
                           d_out2_24_port, QN => net163771);
   registers_reg_31_23_inst : DFFR_X1 port map( D => n3030, CK => n640, RN => 
                           n6155, Q => registers_31_23_port, QN => n5337);
   d_out2_reg_23_inst : DFF_X1 port map( D => n3029, CK => n640, Q => 
                           d_out2_23_port, QN => net163770);
   registers_reg_31_22_inst : DFFR_X1 port map( D => n3028, CK => n640, RN => 
                           n6155, Q => registers_31_22_port, QN => n5336);
   d_out2_reg_22_inst : DFF_X1 port map( D => n3027, CK => n640, Q => 
                           d_out2_22_port, QN => net163769);
   registers_reg_31_21_inst : DFFR_X1 port map( D => n3026, CK => n640, RN => 
                           n6155, Q => registers_31_21_port, QN => n5335);
   d_out2_reg_21_inst : DFF_X1 port map( D => n3025, CK => n640, Q => 
                           d_out2_21_port, QN => net163768);
   registers_reg_31_20_inst : DFFR_X1 port map( D => n3024, CK => n640, RN => 
                           n6155, Q => registers_31_20_port, QN => n5334);
   d_out2_reg_20_inst : DFF_X1 port map( D => n3023, CK => n640, Q => 
                           d_out2_20_port, QN => net163767);
   registers_reg_31_19_inst : DFFR_X1 port map( D => n3022, CK => n640, RN => 
                           n6155, Q => registers_31_19_port, QN => n5333);
   d_out2_reg_19_inst : DFF_X1 port map( D => n3021, CK => n640, Q => 
                           d_out2_19_port, QN => net163766);
   registers_reg_31_18_inst : DFFR_X1 port map( D => n3020, CK => n640, RN => 
                           n6155, Q => registers_31_18_port, QN => n5332);
   d_out2_reg_18_inst : DFF_X1 port map( D => n3019, CK => n640, Q => 
                           d_out2_18_port, QN => net163765);
   registers_reg_31_17_inst : DFFR_X1 port map( D => n3018, CK => n640, RN => 
                           n6155, Q => registers_31_17_port, QN => n5331);
   d_out2_reg_17_inst : DFF_X1 port map( D => n3017, CK => n640, Q => 
                           d_out2_17_port, QN => net163764);
   registers_reg_31_16_inst : DFFR_X1 port map( D => n3016, CK => n640, RN => 
                           n6155, Q => registers_31_16_port, QN => n5330);
   d_out2_reg_16_inst : DFF_X1 port map( D => n3015, CK => n640, Q => 
                           d_out2_16_port, QN => net163763);
   registers_reg_31_15_inst : DFFR_X1 port map( D => n3014, CK => n640, RN => 
                           n6155, Q => registers_31_15_port, QN => n5329);
   d_out2_reg_15_inst : DFF_X1 port map( D => n3013, CK => n640, Q => 
                           d_out2_15_port, QN => net163762);
   registers_reg_31_14_inst : DFFR_X1 port map( D => n3012, CK => n640, RN => 
                           n6155, Q => registers_31_14_port, QN => n5328);
   d_out2_reg_14_inst : DFF_X1 port map( D => n3011, CK => n640, Q => 
                           d_out2_14_port, QN => net163761);
   registers_reg_31_13_inst : DFFR_X1 port map( D => n3010, CK => n640, RN => 
                           n6155, Q => registers_31_13_port, QN => n5327);
   d_out2_reg_13_inst : DFF_X1 port map( D => n3009, CK => n640, Q => 
                           d_out2_13_port, QN => net163760);
   registers_reg_31_12_inst : DFFR_X1 port map( D => n3008, CK => n640, RN => 
                           n6155, Q => registers_31_12_port, QN => n5314);
   d_out2_reg_12_inst : DFF_X1 port map( D => n3007, CK => n640, Q => 
                           d_out2_12_port, QN => net163759);
   registers_reg_31_11_inst : DFFR_X1 port map( D => n3006, CK => n640, RN => 
                           n6154, Q => registers_31_11_port, QN => n5326);
   d_out2_reg_11_inst : DFF_X1 port map( D => n3005, CK => n640, Q => 
                           d_out2_11_port, QN => net163758);
   registers_reg_31_10_inst : DFFR_X1 port map( D => n3004, CK => n640, RN => 
                           n6154, Q => registers_31_10_port, QN => n5325);
   d_out2_reg_10_inst : DFF_X1 port map( D => n3003, CK => n640, Q => 
                           d_out2_10_port, QN => net163757);
   registers_reg_31_9_inst : DFFR_X1 port map( D => n3002, CK => n640, RN => 
                           n6154, Q => registers_31_9_port, QN => n5324);
   d_out2_reg_9_inst : DFF_X1 port map( D => n3001, CK => n640, Q => 
                           d_out2_9_port, QN => net163756);
   registers_reg_31_8_inst : DFFR_X1 port map( D => n3000, CK => n640, RN => 
                           n6154, Q => registers_31_8_port, QN => n5323);
   d_out2_reg_8_inst : DFF_X1 port map( D => n2999, CK => n640, Q => 
                           d_out2_8_port, QN => net163755);
   registers_reg_31_7_inst : DFFR_X1 port map( D => n2998, CK => n640, RN => 
                           n6154, Q => registers_31_7_port, QN => n5322);
   d_out2_reg_7_inst : DFF_X1 port map( D => n2997, CK => n640, Q => 
                           d_out2_7_port, QN => net163754);
   registers_reg_31_6_inst : DFFR_X1 port map( D => n2996, CK => n640, RN => 
                           n6154, Q => registers_31_6_port, QN => n5321);
   d_out2_reg_6_inst : DFF_X1 port map( D => n2995, CK => n640, Q => 
                           d_out2_6_port, QN => net163753);
   registers_reg_31_5_inst : DFFR_X1 port map( D => n2994, CK => n640, RN => 
                           n6154, Q => registers_31_5_port, QN => n5315);
   d_out2_reg_5_inst : DFF_X1 port map( D => n2993, CK => n640, Q => 
                           d_out2_5_port, QN => net163752);
   registers_reg_31_4_inst : DFFR_X1 port map( D => n2992, CK => n640, RN => 
                           n6154, Q => registers_31_4_port, QN => n5320);
   d_out2_reg_4_inst : DFF_X1 port map( D => n2991, CK => n640, Q => 
                           d_out2_4_port, QN => net163751);
   registers_reg_31_3_inst : DFFR_X1 port map( D => n2990, CK => n640, RN => 
                           n6154, Q => registers_31_3_port, QN => n5319);
   d_out2_reg_3_inst : DFF_X1 port map( D => n2989, CK => n640, Q => 
                           d_out2_3_port, QN => net163750);
   registers_reg_31_2_inst : DFFR_X1 port map( D => n2988, CK => n640, RN => 
                           n6156, Q => registers_31_2_port, QN => n5318);
   d_out2_reg_2_inst : DFF_X1 port map( D => n2987, CK => n640, Q => 
                           d_out2_2_port, QN => net163749);
   registers_reg_31_1_inst : DFFR_X1 port map( D => n2986, CK => n640, RN => 
                           n6129, Q => registers_31_1_port, QN => n5317);
   d_out2_reg_1_inst : DFF_X1 port map( D => n2985, CK => n640, Q => 
                           d_out2_1_port, QN => net163748);
   registers_reg_31_0_inst : DFFR_X1 port map( D => n2984, CK => n640, RN => 
                           n6076, Q => registers_31_0_port, QN => n5316);
   d_out2_reg_0_inst : DFF_X1 port map( D => n2983, CK => n640, Q => 
                           d_out2_0_port, QN => net163747);
   d_out1_reg_31_inst : DFF_X1 port map( D => n2982, CK => n640, Q => 
                           d_out1(31), QN => net108160);
   d_out1_reg_30_inst : DFF_X1 port map( D => n2981, CK => n640, Q => 
                           d_out1(30), QN => net108159);
   d_out1_reg_29_inst : DFF_X1 port map( D => n2980, CK => n640, Q => 
                           d_out1(29), QN => net108158);
   d_out1_reg_28_inst : DFF_X1 port map( D => n2979, CK => n640, Q => 
                           d_out1(28), QN => net108157);
   d_out1_reg_27_inst : DFF_X1 port map( D => n2978, CK => n640, Q => 
                           d_out1(27), QN => net108156);
   d_out1_reg_26_inst : DFF_X1 port map( D => n2977, CK => n640, Q => 
                           d_out1(26), QN => net108155);
   d_out1_reg_25_inst : DFF_X1 port map( D => n2976, CK => n640, Q => 
                           d_out1(25), QN => net108154);
   d_out1_reg_24_inst : DFF_X1 port map( D => n2975, CK => n640, Q => 
                           d_out1(24), QN => net108153);
   d_out1_reg_23_inst : DFF_X1 port map( D => n2974, CK => n640, Q => 
                           d_out1(23), QN => net108152);
   d_out1_reg_22_inst : DFF_X1 port map( D => n2973, CK => n640, Q => 
                           d_out1(22), QN => net108151);
   d_out1_reg_21_inst : DFF_X1 port map( D => n2972, CK => n640, Q => 
                           d_out1(21), QN => net108150);
   d_out1_reg_20_inst : DFF_X1 port map( D => n2971, CK => n640, Q => 
                           d_out1(20), QN => net108149);
   d_out1_reg_19_inst : DFF_X1 port map( D => n2970, CK => n640, Q => 
                           d_out1(19), QN => net108148);
   d_out1_reg_18_inst : DFF_X1 port map( D => n2969, CK => n640, Q => 
                           d_out1(18), QN => net108147);
   d_out1_reg_17_inst : DFF_X1 port map( D => n2968, CK => n640, Q => 
                           d_out1(17), QN => net108146);
   d_out1_reg_16_inst : DFF_X1 port map( D => n2967, CK => n640, Q => 
                           d_out1(16), QN => net108145);
   d_out1_reg_15_inst : DFF_X1 port map( D => n2966, CK => n640, Q => 
                           d_out1(15), QN => net108144);
   d_out1_reg_14_inst : DFF_X1 port map( D => n2965, CK => n640, Q => 
                           d_out1(14), QN => net108143);
   d_out1_reg_13_inst : DFF_X1 port map( D => n2964, CK => n640, Q => 
                           d_out1(13), QN => net108142);
   d_out1_reg_12_inst : DFF_X1 port map( D => n2963, CK => n640, Q => 
                           d_out1(12), QN => net108141);
   d_out1_reg_11_inst : DFF_X1 port map( D => n2962, CK => n640, Q => 
                           d_out1(11), QN => net108140);
   d_out1_reg_10_inst : DFF_X1 port map( D => n2961, CK => n640, Q => 
                           d_out1(10), QN => net108139);
   d_out1_reg_9_inst : DFF_X1 port map( D => n2960, CK => n640, Q => d_out1(9),
                           QN => net108138);
   d_out1_reg_8_inst : DFF_X1 port map( D => n2959, CK => n640, Q => d_out1(8),
                           QN => net108137);
   d_out1_reg_7_inst : DFF_X1 port map( D => n2958, CK => n640, Q => d_out1(7),
                           QN => net108136);
   d_out1_reg_6_inst : DFF_X1 port map( D => n2957, CK => n640, Q => d_out1(6),
                           QN => net108135);
   d_out1_reg_5_inst : DFF_X1 port map( D => n2956, CK => n640, Q => d_out1(5),
                           QN => net108134);
   d_out1_reg_4_inst : DFF_X1 port map( D => n2955, CK => n640, Q => d_out1(4),
                           QN => net108133);
   d_out1_reg_3_inst : DFF_X1 port map( D => n2954, CK => n640, Q => d_out1(3),
                           QN => net108132);
   d_out1_reg_2_inst : DFF_X1 port map( D => n2953, CK => n640, Q => d_out1(2),
                           QN => net108131);
   d_out1_reg_1_inst : DFF_X1 port map( D => n2952, CK => n640, Q => d_out1(1),
                           QN => net108130);
   d_out1_reg_0_inst : DFF_X1 port map( D => n2951, CK => n640, Q => d_out1(0),
                           QN => net108129);
   U3 : INV_X2 port map( A => clk, ZN => n640);
   U2064 : NOR3_X2 port map( A1 => rd2_addr(1), A2 => rd2_addr(2), A3 => n5594,
                           ZN => n4427);
   U2070 : NOR3_X2 port map( A1 => n4441, A2 => rd2_addr(1), A3 => n5593, ZN =>
                           n4425);
   U2105 : NOR3_X2 port map( A1 => rd2_addr(0), A2 => rd2_addr(4), A3 => n4461,
                           ZN => n4430);
   U3388 : NOR3_X2 port map( A1 => n5087, A2 => rd1_addr(3), A3 => n5096, ZN =>
                           n5081);
   U3406 : NOR2_X2 port map( A1 => n5090, A2 => rd1_addr(2), ZN => n5078);
   U3409 : NOR3_X2 port map( A1 => rd1_addr(0), A2 => rd1_addr(3), A3 => n5096,
                           ZN => n5088);
   U3430 : NAND3_X1 port map( A1 => n4433, A2 => n4434, A3 => n4425, ZN => 
                           n2749);
   U3431 : NAND3_X1 port map( A1 => n4438, A2 => n4439, A3 => n4440, ZN => 
                           n4414);
   U3432 : NAND3_X1 port map( A1 => n4442, A2 => n4439, A3 => n4440, ZN => 
                           n2750);
   U3433 : NAND3_X1 port map( A1 => n4426, A2 => n4443, A3 => n4440, ZN => 
                           n2755);
   U3435 : NAND3_X1 port map( A1 => n4458, A2 => n4441, A3 => n4442, ZN => 
                           n2726);
   U3436 : NAND3_X1 port map( A1 => n4433, A2 => n4434, A3 => n4443, ZN => 
                           n2731);
   U3437 : NAND3_X1 port map( A1 => rd2_en, A2 => en, A3 => n6156, ZN => n2752)
                           ;
   U3438 : NAND3_X1 port map( A1 => n5067, A2 => n5505, A3 => n5079, ZN => 
                           n4481);
   U3439 : NAND3_X1 port map( A1 => n5078, A2 => n5505, A3 => n5069, ZN => 
                           n4480);
   U3440 : NAND3_X1 port map( A1 => n5086, A2 => n5087, A3 => n5080, ZN => 
                           n4486);
   U3441 : NAND3_X1 port map( A1 => n5081, A2 => n5504, A3 => n5067, ZN => 
                           n4501);
   U3442 : NAND3_X1 port map( A1 => n5078, A2 => n5506, A3 => n5088, ZN => 
                           n4504);
   U3443 : NAND3_X1 port map( A1 => n5081, A2 => n5504, A3 => n5078, ZN => 
                           n4506);
   U3446 : NAND3_X1 port map( A1 => n5078, A2 => n5505, A3 => n5070, ZN => 
                           n4517);
   U4 : NOR3_X1 port map( A1 => rd1_addr(0), A2 => rd1_addr(4), A3 => n5097, ZN
                           => n5084);
   U5 : NOR3_X1 port map( A1 => n5087, A2 => rd1_addr(4), A3 => n5097, ZN => 
                           n5070);
   U6 : NOR3_X1 port map( A1 => n4434, A2 => rd2_addr(3), A3 => n4459, ZN => 
                           n4429);
   U7 : NOR2_X1 port map( A1 => wr_addr(0), A2 => wr_addr(1), ZN => n1803);
   U8 : NOR2_X1 port map( A1 => n5095, A2 => n5090, ZN => n5067);
   U9 : NOR2_X1 port map( A1 => n4458, A2 => rd2_addr(2), ZN => n4439);
   U10 : NOR3_X1 port map( A1 => rd2_addr(0), A2 => rd2_addr(3), A3 => n4459, 
                           ZN => n4428);
   U11 : NOR2_X1 port map( A1 => n2699, A2 => wr_addr(0), ZN => n1730);
   U12 : NOR2_X1 port map( A1 => n2664, A2 => wr_addr(1), ZN => n1694);
   U13 : AND2_X1 port map( A1 => n1765, A2 => n1695, ZN => n2050);
   U14 : BUF_X1 port map( A => n5798, Z => n5378);
   U15 : BUF_X1 port map( A => n5798, Z => n5379);
   U16 : BUF_X1 port map( A => n5798, Z => n5380);
   U17 : BUF_X1 port map( A => n5834, Z => n5390);
   U18 : BUF_X1 port map( A => n5924, Z => n5420);
   U19 : BUF_X1 port map( A => n5835, Z => n5391);
   U20 : BUF_X1 port map( A => n5925, Z => n5421);
   U21 : BUF_X1 port map( A => n5852, Z => n5397);
   U22 : BUF_X1 port map( A => n5852, Z => n5396);
   U23 : BUF_X1 port map( A => n5898, Z => n5411);
   U24 : BUF_X1 port map( A => n5898, Z => n5412);
   U25 : BUF_X1 port map( A => n5699, Z => n5345);
   U26 : BUF_X1 port map( A => n5699, Z => n5346);
   U27 : BUF_X1 port map( A => n5708, Z => n5348);
   U28 : BUF_X1 port map( A => n5708, Z => n5349);
   U29 : BUF_X1 port map( A => n5717, Z => n5351);
   U30 : BUF_X1 port map( A => n5717, Z => n5352);
   U31 : BUF_X1 port map( A => n5726, Z => n5354);
   U32 : BUF_X1 port map( A => n5726, Z => n5355);
   U33 : BUF_X1 port map( A => n5736, Z => n5357);
   U34 : BUF_X1 port map( A => n5736, Z => n5358);
   U35 : BUF_X1 port map( A => n5744, Z => n5360);
   U36 : BUF_X1 port map( A => n5744, Z => n5361);
   U37 : BUF_X1 port map( A => n5753, Z => n5363);
   U38 : BUF_X1 port map( A => n5753, Z => n5364);
   U39 : BUF_X1 port map( A => n5762, Z => n5366);
   U40 : BUF_X1 port map( A => n5762, Z => n5367);
   U41 : BUF_X1 port map( A => n5771, Z => n5369);
   U42 : BUF_X1 port map( A => n5771, Z => n5370);
   U43 : BUF_X1 port map( A => n5780, Z => n5372);
   U44 : BUF_X1 port map( A => n5780, Z => n5373);
   U45 : BUF_X1 port map( A => n5789, Z => n5375);
   U46 : BUF_X1 port map( A => n5789, Z => n5376);
   U47 : BUF_X1 port map( A => n5808, Z => n5381);
   U48 : BUF_X1 port map( A => n5808, Z => n5382);
   U49 : BUF_X1 port map( A => n5817, Z => n5384);
   U50 : BUF_X1 port map( A => n5817, Z => n5385);
   U51 : BUF_X1 port map( A => n5825, Z => n5387);
   U52 : BUF_X1 port map( A => n5825, Z => n5388);
   U53 : BUF_X1 port map( A => n5844, Z => n5393);
   U54 : BUF_X1 port map( A => n5844, Z => n5394);
   U55 : BUF_X1 port map( A => n5862, Z => n5399);
   U56 : BUF_X1 port map( A => n5862, Z => n5400);
   U57 : BUF_X1 port map( A => n5870, Z => n5402);
   U58 : BUF_X1 port map( A => n5870, Z => n5403);
   U59 : BUF_X1 port map( A => n5880, Z => n5405);
   U60 : BUF_X1 port map( A => n5880, Z => n5406);
   U61 : BUF_X1 port map( A => n5888, Z => n5408);
   U62 : BUF_X1 port map( A => n5888, Z => n5409);
   U63 : BUF_X1 port map( A => n5907, Z => n5414);
   U64 : BUF_X1 port map( A => n5907, Z => n5415);
   U65 : BUF_X1 port map( A => n5916, Z => n5417);
   U66 : BUF_X1 port map( A => n5916, Z => n5418);
   U67 : BUF_X1 port map( A => n5933, Z => n5423);
   U68 : BUF_X1 port map( A => n5933, Z => n5424);
   U69 : INV_X1 port map( A => n5952, ZN => n5942);
   U70 : INV_X1 port map( A => n5952, ZN => n5943);
   U71 : BUF_X1 port map( A => n5897, Z => n5413);
   U72 : BUF_X1 port map( A => n5853, Z => n5398);
   U73 : BUF_X1 port map( A => n5700, Z => n5347);
   U74 : BUF_X1 port map( A => n5709, Z => n5350);
   U75 : BUF_X1 port map( A => n5718, Z => n5353);
   U76 : BUF_X1 port map( A => n5726, Z => n5356);
   U77 : BUF_X1 port map( A => n5735, Z => n5359);
   U78 : BUF_X1 port map( A => n5745, Z => n5362);
   U79 : BUF_X1 port map( A => n5754, Z => n5365);
   U80 : BUF_X1 port map( A => n5762, Z => n5368);
   U81 : BUF_X1 port map( A => n5772, Z => n5371);
   U82 : BUF_X1 port map( A => n5781, Z => n5374);
   U83 : BUF_X1 port map( A => n5790, Z => n5377);
   U84 : BUF_X1 port map( A => n5807, Z => n5383);
   U85 : BUF_X1 port map( A => n5816, Z => n5386);
   U86 : BUF_X1 port map( A => n5826, Z => n5389);
   U87 : BUF_X1 port map( A => n5843, Z => n5395);
   U88 : BUF_X1 port map( A => n5861, Z => n5401);
   U89 : BUF_X1 port map( A => n5871, Z => n5404);
   U90 : BUF_X1 port map( A => n5879, Z => n5407);
   U91 : BUF_X1 port map( A => n5889, Z => n5410);
   U92 : BUF_X1 port map( A => n5906, Z => n5416);
   U93 : BUF_X1 port map( A => n5915, Z => n5419);
   U94 : BUF_X1 port map( A => n5933, Z => n5425);
   U95 : BUF_X1 port map( A => n5835, Z => n5392);
   U96 : BUF_X1 port map( A => n5925, Z => n5422);
   U97 : BUF_X1 port map( A => n2050, Z => n5952);
   U98 : BUF_X1 port map( A => n5948, Z => n5951);
   U99 : BUF_X1 port map( A => n5949, Z => n5950);
   U100 : BUF_X1 port map( A => n2050, Z => n5949);
   U101 : BUF_X1 port map( A => n2050, Z => n5948);
   U102 : BUF_X1 port map( A => n2050, Z => n5947);
   U103 : BUF_X1 port map( A => n2050, Z => n5946);
   U104 : BUF_X1 port map( A => n2050, Z => n5945);
   U105 : BUF_X1 port map( A => n2050, Z => n5944);
   U106 : BUF_X1 port map( A => n6157, Z => n6156);
   U107 : INV_X1 port map( A => n5961, ZN => n5954);
   U108 : INV_X1 port map( A => n5961, ZN => n5953);
   U109 : INV_X1 port map( A => n6066, ZN => n6058);
   U110 : INV_X1 port map( A => n6066, ZN => n6059);
   U111 : BUF_X1 port map( A => n2751, Z => n5595);
   U112 : BUF_X1 port map( A => n2751, Z => n5596);
   U113 : BUF_X1 port map( A => n4479, Z => n5590);
   U114 : BUF_X1 port map( A => n4479, Z => n5591);
   U115 : INV_X1 port map( A => n5594, ZN => n4440);
   U116 : BUF_X1 port map( A => n2751, Z => n5597);
   U117 : BUF_X1 port map( A => n4479, Z => n5592);
   U118 : INV_X1 port map( A => n2286, ZN => n5798);
   U119 : INV_X1 port map( A => n2286, ZN => n5799);
   U120 : BUF_X1 port map( A => n6067, Z => n6157);
   U121 : BUF_X1 port map( A => n6067, Z => n6158);
   U122 : BUF_X1 port map( A => n6068, Z => n6160);
   U123 : BUF_X1 port map( A => n6067, Z => n6159);
   U124 : BUF_X1 port map( A => n6068, Z => n6161);
   U125 : BUF_X1 port map( A => n6068, Z => n6162);
   U126 : BUF_X1 port map( A => n6069, Z => n6163);
   U127 : BUF_X1 port map( A => n6069, Z => n6165);
   U128 : BUF_X1 port map( A => n6070, Z => n6168);
   U129 : BUF_X1 port map( A => n6069, Z => n6164);
   U130 : BUF_X1 port map( A => n6070, Z => n6166);
   U131 : BUF_X1 port map( A => n6070, Z => n6167);
   U132 : BUF_X1 port map( A => n6071, Z => n6169);
   U133 : BUF_X1 port map( A => n6071, Z => n6170);
   U134 : INV_X2 port map( A => n4410, ZN => n2709);
   U135 : INV_X2 port map( A => n4414, ZN => n2745);
   U136 : INV_X2 port map( A => n4412, ZN => n2741);
   U137 : NAND2_X1 port map( A1 => n4448, A2 => n4464, ZN => n5594);
   U138 : NAND2_X1 port map( A1 => n4448, A2 => n4464, ZN => n5593);
   U139 : NAND2_X1 port map( A1 => n4448, A2 => n4464, ZN => n2714);
   U140 : BUF_X1 port map( A => n4499, Z => n5535);
   U141 : BUF_X1 port map( A => n4503, Z => n5529);
   U142 : BUF_X1 port map( A => n4499, Z => n5536);
   U143 : BUF_X1 port map( A => n4503, Z => n5530);
   U144 : BUF_X1 port map( A => n2754, Z => n5660);
   U145 : BUF_X1 port map( A => n4511, Z => n5432);
   U146 : BUF_X1 port map( A => n4516, Z => n5426);
   U147 : BUF_X1 port map( A => n4511, Z => n5433);
   U148 : BUF_X1 port map( A => n4516, Z => n5427);
   U149 : BUF_X1 port map( A => n2754, Z => n5661);
   U150 : BUF_X1 port map( A => n4517, Z => n5429);
   U151 : BUF_X1 port map( A => n4517, Z => n5430);
   U152 : BUF_X1 port map( A => n2755, Z => n5478);
   U153 : BUF_X1 port map( A => n2755, Z => n5479);
   U154 : BUF_X1 port map( A => n4500, Z => n5538);
   U155 : BUF_X1 port map( A => n4500, Z => n5539);
   U156 : BUF_X1 port map( A => n4486, Z => n5453);
   U157 : BUF_X1 port map( A => n4486, Z => n5454);
   U158 : BUF_X1 port map( A => n4508, Z => n5512);
   U159 : BUF_X1 port map( A => n4508, Z => n5513);
   U160 : BUF_X1 port map( A => n4513, Z => n5507);
   U161 : BUF_X1 port map( A => n4513, Z => n5508);
   U162 : BUF_X1 port map( A => n4478, Z => n5587);
   U163 : BUF_X1 port map( A => n4478, Z => n5588);
   U164 : BUF_X1 port map( A => n4475, Z => n5584);
   U165 : BUF_X1 port map( A => n4475, Z => n5585);
   U166 : BUF_X1 port map( A => n2750, Z => n5481);
   U167 : BUF_X1 port map( A => n2750, Z => n5482);
   U168 : BUF_X1 port map( A => n4499, Z => n5537);
   U169 : BUF_X1 port map( A => n4503, Z => n5531);
   U170 : BUF_X1 port map( A => n2754, Z => n5662);
   U171 : BUF_X1 port map( A => n4507, Z => n5526);
   U172 : BUF_X1 port map( A => n4507, Z => n5527);
   U173 : BUF_X1 port map( A => n4511, Z => n5434);
   U174 : BUF_X1 port map( A => n4516, Z => n5428);
   U175 : BUF_X1 port map( A => n2715, Z => n5683);
   U176 : BUF_X1 port map( A => n2715, Z => n5684);
   U177 : BUF_X1 port map( A => n2755, Z => n5480);
   U178 : BUF_X1 port map( A => n4517, Z => n5431);
   U179 : BUF_X1 port map( A => n4500, Z => n5540);
   U180 : BUF_X1 port map( A => n4505, Z => n5435);
   U181 : BUF_X1 port map( A => n4505, Z => n5436);
   U182 : BUF_X1 port map( A => n2748, Z => n5665);
   U183 : BUF_X1 port map( A => n2748, Z => n5666);
   U184 : BUF_X1 port map( A => n4484, Z => n5581);
   U185 : BUF_X1 port map( A => n4484, Z => n5582);
   U186 : BUF_X1 port map( A => n4486, Z => n5455);
   U187 : NAND2_X1 port map( A1 => n2217, A2 => n1765, ZN => n2286);
   U188 : BUF_X1 port map( A => n4508, Z => n5514);
   U189 : BUF_X1 port map( A => n4513, Z => n5509);
   U190 : BUF_X1 port map( A => n4478, Z => n5589);
   U191 : BUF_X1 port map( A => n4475, Z => n5586);
   U192 : BUF_X1 port map( A => n2750, Z => n5483);
   U193 : BUF_X1 port map( A => n4507, Z => n5528);
   U194 : BUF_X1 port map( A => n2715, Z => n5685);
   U195 : BUF_X1 port map( A => n4505, Z => n5437);
   U196 : BUF_X1 port map( A => n2748, Z => n5667);
   U197 : BUF_X1 port map( A => n4484, Z => n5583);
   U198 : INV_X1 port map( A => n2743, ZN => n5668);
   U199 : INV_X1 port map( A => n2743, ZN => n5669);
   U200 : AND3_X1 port map( A1 => n5067, A2 => n5505, A3 => n5069, ZN => n4479)
                           ;
   U201 : AND3_X1 port map( A1 => n4438, A2 => n4443, A3 => n4440, ZN => n2751)
                           ;
   U202 : BUF_X1 port map( A => n5068, Z => n5504);
   U203 : INV_X1 port map( A => n1769, ZN => n5933);
   U204 : INV_X1 port map( A => n1769, ZN => n5934);
   U205 : BUF_X1 port map( A => n1628, Z => n6065);
   U206 : BUF_X1 port map( A => n1628, Z => n6064);
   U207 : BUF_X1 port map( A => n1628, Z => n6063);
   U208 : BUF_X1 port map( A => n1628, Z => n6062);
   U209 : BUF_X1 port map( A => n1628, Z => n6061);
   U210 : BUF_X1 port map( A => n1628, Z => n6060);
   U211 : BUF_X1 port map( A => n1698, Z => n5960);
   U212 : BUF_X1 port map( A => n1698, Z => n5959);
   U213 : BUF_X1 port map( A => n1698, Z => n5958);
   U214 : BUF_X1 port map( A => n1698, Z => n5957);
   U215 : BUF_X1 port map( A => n1698, Z => n5956);
   U216 : BUF_X1 port map( A => n1698, Z => n5955);
   U217 : BUF_X1 port map( A => n5068, Z => n5505);
   U218 : INV_X1 port map( A => n4491, ZN => n5543);
   U219 : INV_X1 port map( A => n1805, ZN => n5924);
   U220 : INV_X1 port map( A => n2081, ZN => n5852);
   U221 : INV_X1 port map( A => n2081, ZN => n5853);
   U222 : INV_X1 port map( A => n2665, ZN => n5699);
   U223 : INV_X1 port map( A => n2665, ZN => n5700);
   U224 : INV_X1 port map( A => n2630, ZN => n5708);
   U225 : INV_X1 port map( A => n2630, ZN => n5709);
   U226 : INV_X1 port map( A => n2527, ZN => n5735);
   U227 : INV_X1 port map( A => n2527, ZN => n5736);
   U228 : INV_X1 port map( A => n2493, ZN => n5744);
   U229 : INV_X1 port map( A => n2493, ZN => n5745);
   U230 : INV_X1 port map( A => n2390, ZN => n5771);
   U231 : INV_X1 port map( A => n2390, ZN => n5772);
   U232 : INV_X1 port map( A => n2356, ZN => n5780);
   U233 : INV_X1 port map( A => n2356, ZN => n5781);
   U234 : INV_X1 port map( A => n2252, ZN => n5807);
   U235 : INV_X1 port map( A => n2252, ZN => n5808);
   U236 : INV_X1 port map( A => n2218, ZN => n5816);
   U237 : INV_X1 port map( A => n2218, ZN => n5817);
   U238 : INV_X1 port map( A => n2113, ZN => n5843);
   U239 : INV_X1 port map( A => n2113, ZN => n5844);
   U240 : INV_X1 port map( A => n1976, ZN => n5879);
   U241 : INV_X1 port map( A => n1976, ZN => n5880);
   U242 : INV_X1 port map( A => n1942, ZN => n5888);
   U243 : INV_X1 port map( A => n1942, ZN => n5889);
   U244 : INV_X1 port map( A => n1839, ZN => n5915);
   U245 : INV_X1 port map( A => n1839, ZN => n5916);
   U246 : INV_X1 port map( A => n1805, ZN => n5925);
   U247 : INV_X1 port map( A => n2147, ZN => n5834);
   U248 : INV_X1 port map( A => n2561, ZN => n5726);
   U249 : INV_X1 port map( A => n2561, ZN => n5727);
   U250 : INV_X1 port map( A => n2424, ZN => n5762);
   U251 : INV_X1 port map( A => n2424, ZN => n5763);
   U252 : INV_X1 port map( A => n2147, ZN => n5835);
   U253 : INV_X1 port map( A => n2010, ZN => n5870);
   U254 : INV_X1 port map( A => n2010, ZN => n5871);
   U255 : INV_X1 port map( A => n1873, ZN => n5906);
   U256 : INV_X1 port map( A => n1873, ZN => n5907);
   U257 : BUF_X1 port map( A => n1628, Z => n6066);
   U258 : INV_X1 port map( A => n5681, ZN => n4423);
   U259 : INV_X1 port map( A => n1909, ZN => n5898);
   U260 : INV_X1 port map( A => n1909, ZN => n5897);
   U261 : INV_X1 port map( A => n2595, ZN => n5717);
   U262 : INV_X1 port map( A => n2595, ZN => n5718);
   U263 : INV_X1 port map( A => n2458, ZN => n5753);
   U264 : INV_X1 port map( A => n2458, ZN => n5754);
   U265 : INV_X1 port map( A => n2321, ZN => n5789);
   U266 : INV_X1 port map( A => n2321, ZN => n5790);
   U267 : INV_X1 port map( A => n2183, ZN => n5825);
   U268 : INV_X1 port map( A => n2183, ZN => n5826);
   U269 : INV_X1 port map( A => n2044, ZN => n5861);
   U270 : INV_X1 port map( A => n2044, ZN => n5862);
   U271 : BUF_X1 port map( A => n1698, Z => n5961);
   U272 : BUF_X1 port map( A => n5563, Z => n5565);
   U273 : BUF_X1 port map( A => n5563, Z => n5566);
   U274 : BUF_X1 port map( A => n5563, Z => n5567);
   U275 : BUF_X1 port map( A => n5563, Z => n5568);
   U276 : BUF_X1 port map( A => n5564, Z => n5569);
   U277 : BUF_X1 port map( A => n5564, Z => n5570);
   U278 : BUF_X1 port map( A => n5564, Z => n5571);
   U279 : BUF_X1 port map( A => n5564, Z => n5572);
   U280 : BUF_X1 port map( A => n5068, Z => n5503);
   U281 : BUF_X1 port map( A => n5068, Z => n5506);
   U282 : BUF_X1 port map( A => n4488, Z => n5573);
   U283 : BUF_X1 port map( A => n4488, Z => n5574);
   U284 : BUF_X1 port map( A => n4488, Z => n5575);
   U285 : BUF_X1 port map( A => n4488, Z => n5576);
   U286 : BUF_X1 port map( A => n2733, Z => n5637);
   U287 : BUF_X1 port map( A => n2733, Z => n5638);
   U288 : BUF_X1 port map( A => n2724, Z => n5657);
   U289 : BUF_X1 port map( A => n2724, Z => n5658);
   U290 : BUF_X1 port map( A => n2733, Z => n5639);
   U291 : BUF_X1 port map( A => n2724, Z => n5659);
   U292 : INV_X1 port map( A => n5466, ZN => n4448);
   U293 : BUF_X1 port map( A => n6073, Z => n6067);
   U294 : BUF_X1 port map( A => n2731, Z => n5469);
   U295 : BUF_X1 port map( A => n2731, Z => n5470);
   U296 : BUF_X1 port map( A => n2726, Z => n5472);
   U297 : BUF_X1 port map( A => n2726, Z => n5473);
   U298 : BUF_X1 port map( A => n2721, Z => n5475);
   U299 : BUF_X1 port map( A => n2721, Z => n5476);
   U300 : BUF_X1 port map( A => n2731, Z => n5471);
   U301 : BUF_X1 port map( A => n2726, Z => n5474);
   U302 : BUF_X1 port map( A => n2721, Z => n5477);
   U303 : INV_X1 port map( A => n2730, ZN => n5629);
   U304 : INV_X1 port map( A => n2735, ZN => n5598);
   U305 : BUF_X1 port map( A => n5606, Z => n5607);
   U306 : BUF_X1 port map( A => n5606, Z => n5608);
   U307 : BUF_X1 port map( A => n5648, Z => n5649);
   U308 : BUF_X1 port map( A => n5648, Z => n5650);
   U309 : BUF_X1 port map( A => n5606, Z => n5609);
   U310 : BUF_X1 port map( A => n2736, Z => n5610);
   U311 : BUF_X1 port map( A => n2736, Z => n5611);
   U312 : BUF_X1 port map( A => n2736, Z => n5612);
   U313 : BUF_X1 port map( A => n5648, Z => n5651);
   U314 : BUF_X1 port map( A => n2720, Z => n5652);
   U315 : BUF_X1 port map( A => n2720, Z => n5653);
   U316 : BUF_X1 port map( A => n2720, Z => n5654);
   U317 : BUF_X1 port map( A => n6072, Z => n6069);
   U318 : BUF_X1 port map( A => n6072, Z => n6070);
   U319 : BUF_X1 port map( A => n6073, Z => n6068);
   U320 : BUF_X1 port map( A => n6072, Z => n6071);
   U321 : NOR2_X1 port map( A1 => n2699, A2 => n2664, ZN => n1765);
   U322 : INV_X2 port map( A => n4418, ZN => n2700);
   U323 : NAND2_X1 port map( A1 => n4425, A2 => n4430, ZN => n5682);
   U324 : NAND2_X1 port map( A1 => n4425, A2 => n4430, ZN => n5681);
   U325 : NAND2_X1 port map( A1 => n4425, A2 => n4430, ZN => n2744);
   U326 : NAND2_X1 port map( A1 => n4427, A2 => n4428, ZN => n5687);
   U327 : NAND2_X1 port map( A1 => n4427, A2 => n4428, ZN => n5686);
   U328 : NAND2_X1 port map( A1 => n4427, A2 => n4428, ZN => n2712);
   U329 : NAND2_X1 port map( A1 => n5080, A2 => n5088, ZN => n5561);
   U330 : NAND2_X1 port map( A1 => n5080, A2 => n5088, ZN => n5562);
   U331 : NAND2_X1 port map( A1 => n5083, A2 => n5070, ZN => n5541);
   U332 : NAND2_X1 port map( A1 => n5083, A2 => n5070, ZN => n5542);
   U333 : AND2_X1 port map( A1 => n4427, A2 => n4430, ZN => n5678);
   U334 : AND2_X1 port map( A1 => n4427, A2 => n4430, ZN => n5677);
   U335 : AND3_X1 port map( A1 => n4442, A2 => n4443, A3 => n4440, ZN => n2746)
                           ;
   U336 : AND3_X1 port map( A1 => n4442, A2 => n4443, A3 => n4440, ZN => n5663)
                           ;
   U337 : AND2_X1 port map( A1 => n4427, A2 => n4426, ZN => n5680);
   U338 : AND2_X1 port map( A1 => n4427, A2 => n4426, ZN => n5679);
   U339 : AND2_X1 port map( A1 => n5083, A2 => n5088, ZN => n5510);
   U340 : AND2_X1 port map( A1 => n5083, A2 => n5088, ZN => n5511);
   U341 : AND2_X1 port map( A1 => n5083, A2 => n5081, ZN => n5551);
   U342 : AND2_X1 port map( A1 => n5080, A2 => n5081, ZN => n5579);
   U343 : AND2_X1 port map( A1 => n5083, A2 => n5081, ZN => n5552);
   U344 : AND2_X1 port map( A1 => n5080, A2 => n5081, ZN => n5580);
   U345 : OAI222_X1 port map( A1 => n5238, A2 => n5684, B1 => n2154, B2 => 
                           n5686, C1 => n2479, C2 => n4410, ZN => n4424);
   U346 : OAI222_X1 port map( A1 => n5215, A2 => n5666, B1 => n2121, B2 => 
                           n5486, C1 => n2455, C2 => n5482, ZN => n4413);
   U347 : OAI222_X1 port map( A1 => n5216, A2 => n5665, B1 => n2122, B2 => 
                           n5488, C1 => n2456, C2 => n5481, ZN => n4392);
   U348 : OAI222_X1 port map( A1 => n5217, A2 => n5667, B1 => n2123, B2 => 
                           n5487, C1 => n2457, C2 => n5481, ZN => n4373);
   U349 : OAI222_X1 port map( A1 => n5218, A2 => n5665, B1 => n2124, B2 => 
                           n5487, C1 => n2459, C2 => n5483, ZN => n4354);
   U350 : OAI222_X1 port map( A1 => n5219, A2 => n5666, B1 => n2125, B2 => 
                           n5486, C1 => n2460, C2 => n5482, ZN => n4335);
   U351 : OAI222_X1 port map( A1 => n5220, A2 => n5666, B1 => n2126, B2 => 
                           n5488, C1 => n2461, C2 => n5482, ZN => n4316);
   U352 : OAI222_X1 port map( A1 => n5221, A2 => n5667, B1 => n2127, B2 => 
                           n5488, C1 => n2462, C2 => n5481, ZN => n4297);
   U353 : OAI222_X1 port map( A1 => n5222, A2 => n5667, B1 => n2140, B2 => 
                           n5487, C1 => n2463, C2 => n5483, ZN => n4278);
   U354 : OAI222_X1 port map( A1 => n5223, A2 => n5665, B1 => n2128, B2 => 
                           n5486, C1 => n2464, C2 => n5483, ZN => n4259);
   U355 : OAI222_X1 port map( A1 => n5224, A2 => n5666, B1 => n2129, B2 => 
                           n5486, C1 => n2465, C2 => n5482, ZN => n4240);
   U356 : OAI222_X1 port map( A1 => n5225, A2 => n5665, B1 => n2130, B2 => 
                           n5488, C1 => n2466, C2 => n5481, ZN => n4221);
   U357 : OAI222_X1 port map( A1 => n5226, A2 => n5667, B1 => n2131, B2 => 
                           n5487, C1 => n2467, C2 => n5481, ZN => n4202);
   U358 : OAI222_X1 port map( A1 => n5227, A2 => n5665, B1 => n2132, B2 => 
                           n5487, C1 => n2468, C2 => n5483, ZN => n4183);
   U359 : OAI222_X1 port map( A1 => n5228, A2 => n5666, B1 => n2133, B2 => 
                           n5486, C1 => n2469, C2 => n5482, ZN => n4164);
   U360 : OAI222_X1 port map( A1 => n5229, A2 => n5666, B1 => n2134, B2 => 
                           n5488, C1 => n2470, C2 => n5482, ZN => n4145);
   U361 : OAI222_X1 port map( A1 => n5230, A2 => n5667, B1 => n2135, B2 => 
                           n5488, C1 => n2471, C2 => n5481, ZN => n4126);
   U362 : OAI222_X1 port map( A1 => n5231, A2 => n5667, B1 => n2150, B2 => 
                           n5487, C1 => n2472, C2 => n5483, ZN => n4107);
   U363 : OAI222_X1 port map( A1 => n5232, A2 => n5665, B1 => n2136, B2 => 
                           n5486, C1 => n2473, C2 => n5483, ZN => n4088);
   U364 : OAI222_X1 port map( A1 => n5233, A2 => n5666, B1 => n2137, B2 => 
                           n5486, C1 => n2474, C2 => n5482, ZN => n4069);
   U365 : OAI222_X1 port map( A1 => n5234, A2 => n5665, B1 => n2141, B2 => 
                           n5488, C1 => n2475, C2 => n5481, ZN => n4050);
   U366 : OAI222_X1 port map( A1 => n5235, A2 => n5667, B1 => n2142, B2 => 
                           n5487, C1 => n2476, C2 => n5481, ZN => n4031);
   U367 : OAI222_X1 port map( A1 => n5236, A2 => n5665, B1 => n2143, B2 => 
                           n5487, C1 => n2477, C2 => n5483, ZN => n4012);
   U368 : OAI222_X1 port map( A1 => n5237, A2 => n5666, B1 => n2144, B2 => 
                           n5486, C1 => n2478, C2 => n5482, ZN => n2906);
   U369 : OAI222_X1 port map( A1 => n5239, A2 => n5666, B1 => n2145, B2 => 
                           n5488, C1 => n2480, C2 => n5482, ZN => n2887);
   U370 : OAI222_X1 port map( A1 => n5240, A2 => n5667, B1 => n2146, B2 => 
                           n5488, C1 => n2481, C2 => n5481, ZN => n2868);
   U371 : OAI222_X1 port map( A1 => n5241, A2 => n5667, B1 => n2151, B2 => 
                           n5487, C1 => n2482, C2 => n5483, ZN => n2849);
   U372 : OAI222_X1 port map( A1 => n5242, A2 => n5665, B1 => n2148, B2 => 
                           n5486, C1 => n2483, C2 => n5483, ZN => n2830);
   U373 : OAI222_X1 port map( A1 => n5243, A2 => n5666, B1 => n2149, B2 => 
                           n5486, C1 => n2484, C2 => n5482, ZN => n2811);
   U374 : OAI222_X1 port map( A1 => n5244, A2 => n5665, B1 => n2152, B2 => 
                           n5488, C1 => n2485, C2 => n5481, ZN => n2792);
   U375 : OAI222_X1 port map( A1 => n5245, A2 => n5667, B1 => n2138, B2 => 
                           n5487, C1 => n2486, C2 => n5481, ZN => n2773);
   U376 : OAI222_X1 port map( A1 => n5246, A2 => n5665, B1 => n2139, B2 => 
                           n5487, C1 => n2487, C2 => n5483, ZN => n2747);
   U377 : OAI222_X1 port map( A1 => n5247, A2 => n5436, B1 => n2389, B2 => 
                           n5441, C1 => n2153, C2 => n5527, ZN => n5091);
   U378 : OAI222_X1 port map( A1 => n5248, A2 => n5437, B1 => n2391, B2 => 
                           n5442, C1 => n2051, C2 => n5528, ZN => n5052);
   U379 : OAI222_X1 port map( A1 => n5249, A2 => n5435, B1 => n2392, B2 => 
                           n5440, C1 => n2052, C2 => n5526, ZN => n5034);
   U380 : OAI222_X1 port map( A1 => n5250, A2 => n5435, B1 => n2393, B2 => 
                           n5440, C1 => n2053, C2 => n5526, ZN => n5016);
   U381 : OAI222_X1 port map( A1 => n5251, A2 => n5436, B1 => n2394, B2 => 
                           n5441, C1 => n2054, C2 => n5527, ZN => n4998);
   U382 : OAI222_X1 port map( A1 => n5252, A2 => n5436, B1 => n2395, B2 => 
                           n5441, C1 => n2055, C2 => n5527, ZN => n4980);
   U383 : OAI222_X1 port map( A1 => n5253, A2 => n5437, B1 => n2396, B2 => 
                           n5442, C1 => n2056, C2 => n5528, ZN => n4962);
   U384 : OAI222_X1 port map( A1 => n5254, A2 => n5435, B1 => n2397, B2 => 
                           n5440, C1 => n2057, C2 => n5526, ZN => n4944);
   U385 : OAI222_X1 port map( A1 => n5255, A2 => n5437, B1 => n2398, B2 => 
                           n5442, C1 => n2058, C2 => n5528, ZN => n4926);
   U386 : OAI222_X1 port map( A1 => n5256, A2 => n5436, B1 => n2399, B2 => 
                           n5441, C1 => n2059, C2 => n5527, ZN => n4908);
   U387 : OAI222_X1 port map( A1 => n5257, A2 => n5437, B1 => n2400, B2 => 
                           n5442, C1 => n2060, C2 => n5528, ZN => n4890);
   U388 : OAI222_X1 port map( A1 => n5258, A2 => n5435, B1 => n2401, B2 => 
                           n5440, C1 => n2061, C2 => n5526, ZN => n4872);
   U389 : OAI222_X1 port map( A1 => n5259, A2 => n5435, B1 => n2402, B2 => 
                           n5440, C1 => n2062, C2 => n5526, ZN => n4854);
   U390 : OAI222_X1 port map( A1 => n5260, A2 => n5436, B1 => n2403, B2 => 
                           n5441, C1 => n2063, C2 => n5527, ZN => n4836);
   U391 : OAI222_X1 port map( A1 => n5261, A2 => n5436, B1 => n2404, B2 => 
                           n5441, C1 => n2064, C2 => n5527, ZN => n4818);
   U392 : OAI222_X1 port map( A1 => n5262, A2 => n5437, B1 => n2405, B2 => 
                           n5442, C1 => n2065, C2 => n5528, ZN => n4800);
   U393 : OAI222_X1 port map( A1 => n5263, A2 => n5435, B1 => n2406, B2 => 
                           n5440, C1 => n2066, C2 => n5526, ZN => n4782);
   U394 : OAI222_X1 port map( A1 => n5264, A2 => n5437, B1 => n2407, B2 => 
                           n5442, C1 => n2067, C2 => n5528, ZN => n4764);
   U395 : OAI222_X1 port map( A1 => n5265, A2 => n5436, B1 => n2408, B2 => 
                           n5441, C1 => n2068, C2 => n5527, ZN => n4746);
   U396 : OAI222_X1 port map( A1 => n5266, A2 => n5437, B1 => n2409, B2 => 
                           n5442, C1 => n2069, C2 => n5528, ZN => n4728);
   U397 : OAI222_X1 port map( A1 => n5267, A2 => n5435, B1 => n2410, B2 => 
                           n5440, C1 => n2070, C2 => n5526, ZN => n4710);
   U398 : OAI222_X1 port map( A1 => n5268, A2 => n5435, B1 => n2411, B2 => 
                           n5440, C1 => n2071, C2 => n5526, ZN => n4692);
   U399 : OAI222_X1 port map( A1 => n5269, A2 => n5436, B1 => n2412, B2 => 
                           n5441, C1 => n2072, C2 => n5527, ZN => n4674);
   U400 : OAI222_X1 port map( A1 => n5270, A2 => n5436, B1 => n2413, B2 => 
                           n5441, C1 => n2073, C2 => n5527, ZN => n4656);
   U401 : OAI222_X1 port map( A1 => n5271, A2 => n5437, B1 => n2414, B2 => 
                           n5442, C1 => n2074, C2 => n5528, ZN => n4638);
   U402 : OAI222_X1 port map( A1 => n5272, A2 => n5435, B1 => n2415, B2 => 
                           n5440, C1 => n2075, C2 => n5526, ZN => n4620);
   U403 : OAI222_X1 port map( A1 => n5273, A2 => n5437, B1 => n2416, B2 => 
                           n5442, C1 => n2076, C2 => n5528, ZN => n4602);
   U404 : OAI222_X1 port map( A1 => n5274, A2 => n5436, B1 => n2417, B2 => 
                           n5441, C1 => n2077, C2 => n5527, ZN => n4584);
   U405 : OAI222_X1 port map( A1 => n5275, A2 => n5437, B1 => n2418, B2 => 
                           n5442, C1 => n2080, C2 => n5528, ZN => n4566);
   U406 : OAI222_X1 port map( A1 => n5276, A2 => n5435, B1 => n2419, B2 => 
                           n5440, C1 => n2112, C2 => n5526, ZN => n4548);
   U407 : OAI222_X1 port map( A1 => n5277, A2 => n5435, B1 => n2420, B2 => 
                           n5440, C1 => n2114, C2 => n5526, ZN => n4530);
   U408 : OAI222_X1 port map( A1 => n5278, A2 => n5436, B1 => n2421, B2 => 
                           n5441, C1 => n2115, C2 => n5527, ZN => n4495);
   U409 : AND2_X1 port map( A1 => n5083, A2 => n5084, ZN => n5577);
   U410 : AND2_X1 port map( A1 => n5083, A2 => n5084, ZN => n5578);
   U411 : NAND2_X1 port map( A1 => n5080, A2 => n5088, ZN => n4485);
   U412 : NAND2_X1 port map( A1 => n5083, A2 => n5070, ZN => n4490);
   U413 : AND2_X1 port map( A1 => n4427, A2 => n4430, ZN => n2740);
   U414 : NAND4_X1 port map( A1 => n5071, A2 => n5072, A3 => n5491, A4 => n5073
                           , ZN => n4475);
   U415 : NOR4_X1 port map( A1 => n2182, A2 => n5074, A3 => n5075, A4 => n5076,
                           ZN => n5073);
   U416 : NAND4_X1 port map( A1 => n4446, A2 => n4447, A3 => n4448, A4 => n4449
                           , ZN => n2754);
   U417 : NOR4_X1 port map( A1 => n2182, A2 => n4450, A3 => n4451, A4 => n4452,
                           ZN => n4449);
   U418 : AND3_X1 port map( A1 => n4442, A2 => n4443, A3 => n4440, ZN => n5664)
                           ;
   U419 : AND2_X1 port map( A1 => n4427, A2 => n4426, ZN => n2710);
   U420 : AND2_X1 port map( A1 => n5083, A2 => n5088, ZN => n4514);
   U421 : AND2_X1 port map( A1 => n5083, A2 => n5081, ZN => n4493);
   U422 : AND2_X1 port map( A1 => n5080, A2 => n5081, ZN => n4483);
   U423 : AND2_X1 port map( A1 => n5083, A2 => n5084, ZN => n4489);
   U424 : NAND3_X1 port map( A1 => n5088, A2 => n5504, A3 => n5067, ZN => n4505
                           );
   U425 : NAND2_X1 port map( A1 => n4425, A2 => n4435, ZN => n2743);
   U426 : AND3_X1 port map( A1 => n5090, A2 => n5095, A3 => n5506, ZN => n5083)
                           ;
   U427 : NAND4_X1 port map( A1 => n5069, A2 => n5505, A3 => n5090, A4 => n5095
                           , ZN => n4503);
   U428 : NAND4_X1 port map( A1 => n5079, A2 => n5504, A3 => n5090, A4 => n5095
                           , ZN => n4500);
   U429 : NAND2_X1 port map( A1 => n4425, A2 => n4429, ZN => n2748);
   U430 : NAND4_X1 port map( A1 => n5086, A2 => n5067, A3 => n5504, A4 => n5087
                           , ZN => n4499);
   U431 : OAI22_X1 port map( A1 => n2523, A2 => n5670, B1 => n2288, B2 => n5682
                           , ZN => n4411);
   U432 : OAI22_X1 port map( A1 => n2526, A2 => n5675, B1 => n2291, B2 => n5682
                           , ZN => n4353);
   U433 : OAI22_X1 port map( A1 => n2530, A2 => n5673, B1 => n2294, B2 => n5682
                           , ZN => n4296);
   U434 : OAI22_X1 port map( A1 => n2533, A2 => n5674, B1 => n2297, B2 => n5682
                           , ZN => n4239);
   U435 : OAI22_X1 port map( A1 => n2536, A2 => n5672, B1 => n2300, B2 => n5682
                           , ZN => n4182);
   U436 : OAI22_X1 port map( A1 => n2539, A2 => n5673, B1 => n2303, B2 => n5682
                           , ZN => n4125);
   U437 : OAI22_X1 port map( A1 => n2542, A2 => n5674, B1 => n2306, B2 => n5682
                           , ZN => n4068);
   U438 : OAI22_X1 port map( A1 => n2546, A2 => n5670, B1 => n2318, B2 => n5682
                           , ZN => n2742);
   U439 : OAI22_X1 port map( A1 => n2525, A2 => n5674, B1 => n2290, B2 => n5681
                           , ZN => n4372);
   U440 : OAI22_X1 port map( A1 => n2529, A2 => n5672, B1 => n2293, B2 => n5681
                           , ZN => n4315);
   U441 : OAI22_X1 port map( A1 => n2532, A2 => n5673, B1 => n2296, B2 => n5681
                           , ZN => n4258);
   U442 : OAI22_X1 port map( A1 => n2535, A2 => n5671, B1 => n2299, B2 => n5681
                           , ZN => n4201);
   U443 : OAI22_X1 port map( A1 => n2538, A2 => n5673, B1 => n2302, B2 => n5681
                           , ZN => n4144);
   U444 : OAI22_X1 port map( A1 => n2541, A2 => n5672, B1 => n2305, B2 => n5681
                           , ZN => n4087);
   U445 : OAI22_X1 port map( A1 => n2544, A2 => n5674, B1 => n2308, B2 => n5681
                           , ZN => n4030);
   U446 : OAI22_X1 port map( A1 => n2545, A2 => n5670, B1 => n2317, B2 => n5681
                           , ZN => n2772);
   U447 : NAND2_X1 port map( A1 => n4425, A2 => n4428, ZN => n4412);
   U448 : NAND2_X1 port map( A1 => n4425, A2 => n4426, ZN => n4410);
   U449 : OAI22_X1 port map( A1 => n2524, A2 => n5670, B1 => n2289, B2 => n2744
                           , ZN => n4391);
   U450 : OAI22_X1 port map( A1 => n2528, A2 => n5671, B1 => n2292, B2 => n2744
                           , ZN => n4334);
   U451 : OAI22_X1 port map( A1 => n2531, A2 => n5672, B1 => n2295, B2 => n2744
                           , ZN => n4277);
   U452 : OAI22_X1 port map( A1 => n2534, A2 => n5672, B1 => n2298, B2 => n2744
                           , ZN => n4220);
   U453 : OAI22_X1 port map( A1 => n2537, A2 => n5673, B1 => n2301, B2 => n2744
                           , ZN => n4163);
   U454 : OAI22_X1 port map( A1 => n2540, A2 => n5671, B1 => n2304, B2 => n2744
                           , ZN => n4106);
   U455 : OAI22_X1 port map( A1 => n2543, A2 => n5671, B1 => n2307, B2 => n2744
                           , ZN => n4049);
   U456 : NAND3_X1 port map( A1 => n5078, A2 => n5503, A3 => n5084, ZN => n4516
                           );
   U457 : NAND2_X1 port map( A1 => n4427, A2 => n4429, ZN => n2715);
   U458 : NAND3_X1 port map( A1 => n5067, A2 => n5503, A3 => n5084, ZN => n4511
                           );
   U459 : OAI22_X1 port map( A1 => n2511, A2 => n5486, B1 => n2224, B2 => n4412
                           , ZN => n4432);
   U460 : OAI22_X1 port map( A1 => n2227, A2 => n5536, B1 => n2512, B2 => n5539
                           , ZN => n5094);
   U461 : OAI22_X1 port map( A1 => n2258, A2 => n5537, B1 => n2488, B2 => n5540
                           , ZN => n5055);
   U462 : OAI22_X1 port map( A1 => n2259, A2 => n5535, B1 => n2513, B2 => n5538
                           , ZN => n5037);
   U463 : OAI22_X1 port map( A1 => n2260, A2 => n5535, B1 => n2489, B2 => n5538
                           , ZN => n5019);
   U464 : OAI22_X1 port map( A1 => n2261, A2 => n5536, B1 => n2490, B2 => n5539
                           , ZN => n5001);
   U465 : OAI22_X1 port map( A1 => n2262, A2 => n5536, B1 => n2514, B2 => n5539
                           , ZN => n4983);
   U466 : OAI22_X1 port map( A1 => n2263, A2 => n5537, B1 => n2491, B2 => n5540
                           , ZN => n4965);
   U467 : OAI22_X1 port map( A1 => n2264, A2 => n5535, B1 => n2494, B2 => n5538
                           , ZN => n4947);
   U468 : OAI22_X1 port map( A1 => n2265, A2 => n5537, B1 => n2515, B2 => n5540
                           , ZN => n4929);
   U469 : OAI22_X1 port map( A1 => n2266, A2 => n5536, B1 => n2495, B2 => n5539
                           , ZN => n4911);
   U470 : OAI22_X1 port map( A1 => n2267, A2 => n5537, B1 => n2496, B2 => n5540
                           , ZN => n4893);
   U471 : OAI22_X1 port map( A1 => n2268, A2 => n5535, B1 => n2516, B2 => n5538
                           , ZN => n4875);
   U472 : OAI22_X1 port map( A1 => n2269, A2 => n5535, B1 => n2497, B2 => n5538
                           , ZN => n4857);
   U473 : OAI22_X1 port map( A1 => n2270, A2 => n5536, B1 => n2498, B2 => n5539
                           , ZN => n4839);
   U474 : OAI22_X1 port map( A1 => n2271, A2 => n5536, B1 => n2517, B2 => n5539
                           , ZN => n4821);
   U475 : OAI22_X1 port map( A1 => n2272, A2 => n5537, B1 => n2499, B2 => n5540
                           , ZN => n4803);
   U476 : OAI22_X1 port map( A1 => n2273, A2 => n5535, B1 => n2500, B2 => n5538
                           , ZN => n4785);
   U477 : OAI22_X1 port map( A1 => n2274, A2 => n5537, B1 => n2518, B2 => n5540
                           , ZN => n4767);
   U478 : OAI22_X1 port map( A1 => n2275, A2 => n5536, B1 => n2501, B2 => n5539
                           , ZN => n4749);
   U479 : OAI22_X1 port map( A1 => n2276, A2 => n5537, B1 => n2502, B2 => n5540
                           , ZN => n4731);
   U480 : OAI22_X1 port map( A1 => n2277, A2 => n5535, B1 => n2519, B2 => n5538
                           , ZN => n4713);
   U481 : OAI22_X1 port map( A1 => n2278, A2 => n5535, B1 => n2503, B2 => n5538
                           , ZN => n4695);
   U482 : OAI22_X1 port map( A1 => n2279, A2 => n5536, B1 => n2504, B2 => n5539
                           , ZN => n4677);
   U483 : OAI22_X1 port map( A1 => n2280, A2 => n5536, B1 => n2520, B2 => n5539
                           , ZN => n4659);
   U484 : OAI22_X1 port map( A1 => n2281, A2 => n5537, B1 => n2505, B2 => n5540
                           , ZN => n4641);
   U485 : OAI22_X1 port map( A1 => n2282, A2 => n5535, B1 => n2506, B2 => n5538
                           , ZN => n4623);
   U486 : OAI22_X1 port map( A1 => n2119, A2 => n5537, B1 => n2521, B2 => n5540
                           , ZN => n4605);
   U487 : OAI22_X1 port map( A1 => n2120, A2 => n5536, B1 => n2507, B2 => n5539
                           , ZN => n4587);
   U488 : OAI22_X1 port map( A1 => n2283, A2 => n5537, B1 => n2508, B2 => n5540
                           , ZN => n4569);
   U489 : OAI22_X1 port map( A1 => n2284, A2 => n5535, B1 => n2522, B2 => n5538
                           , ZN => n4551);
   U490 : OAI22_X1 port map( A1 => n2285, A2 => n5535, B1 => n2509, B2 => n5538
                           , ZN => n4533);
   U491 : OAI22_X1 port map( A1 => n2287, A2 => n5536, B1 => n2510, B2 => n5539
                           , ZN => n4498);
   U492 : OAI22_X1 port map( A1 => n2223, A2 => n5451, B1 => n2614, B2 => n5533
                           , ZN => n5093);
   U493 : OAI22_X1 port map( A1 => n2155, A2 => n5452, B1 => n2615, B2 => n5534
                           , ZN => n5054);
   U494 : OAI22_X1 port map( A1 => n2176, A2 => n5450, B1 => n2616, B2 => n5532
                           , ZN => n5036);
   U495 : OAI22_X1 port map( A1 => n2156, A2 => n5450, B1 => n2617, B2 => n5532
                           , ZN => n5018);
   U496 : OAI22_X1 port map( A1 => n2157, A2 => n5451, B1 => n2618, B2 => n5533
                           , ZN => n5000);
   U497 : OAI22_X1 port map( A1 => n2177, A2 => n5451, B1 => n2619, B2 => n5533
                           , ZN => n4982);
   U498 : OAI22_X1 port map( A1 => n2158, A2 => n5452, B1 => n2620, B2 => n5534
                           , ZN => n4964);
   U499 : OAI22_X1 port map( A1 => n2159, A2 => n5450, B1 => n2621, B2 => n5532
                           , ZN => n4946);
   U500 : OAI22_X1 port map( A1 => n2178, A2 => n5452, B1 => n2622, B2 => n5534
                           , ZN => n4928);
   U501 : OAI22_X1 port map( A1 => n2160, A2 => n5451, B1 => n2623, B2 => n5533
                           , ZN => n4910);
   U502 : OAI22_X1 port map( A1 => n2161, A2 => n5452, B1 => n2624, B2 => n5534
                           , ZN => n4892);
   U503 : OAI22_X1 port map( A1 => n2179, A2 => n5450, B1 => n2625, B2 => n5532
                           , ZN => n4874);
   U504 : OAI22_X1 port map( A1 => n2162, A2 => n5450, B1 => n2626, B2 => n5532
                           , ZN => n4856);
   U505 : OAI22_X1 port map( A1 => n2163, A2 => n5451, B1 => n2627, B2 => n5533
                           , ZN => n4838);
   U506 : OAI22_X1 port map( A1 => n2184, A2 => n5451, B1 => n2628, B2 => n5533
                           , ZN => n4820);
   U507 : OAI22_X1 port map( A1 => n2164, A2 => n5452, B1 => n2631, B2 => n5534
                           , ZN => n4802);
   U508 : OAI22_X1 port map( A1 => n2165, A2 => n5450, B1 => n2632, B2 => n5532
                           , ZN => n4784);
   U509 : OAI22_X1 port map( A1 => n2185, A2 => n5452, B1 => n2633, B2 => n5534
                           , ZN => n4766);
   U510 : OAI22_X1 port map( A1 => n2166, A2 => n5451, B1 => n2634, B2 => n5533
                           , ZN => n4748);
   U511 : OAI22_X1 port map( A1 => n2167, A2 => n5452, B1 => n2635, B2 => n5534
                           , ZN => n4730);
   U512 : OAI22_X1 port map( A1 => n2186, A2 => n5450, B1 => n2636, B2 => n5532
                           , ZN => n4712);
   U513 : OAI22_X1 port map( A1 => n2168, A2 => n5450, B1 => n2637, B2 => n5532
                           , ZN => n4694);
   U514 : OAI22_X1 port map( A1 => n2169, A2 => n5451, B1 => n2638, B2 => n5533
                           , ZN => n4676);
   U515 : OAI22_X1 port map( A1 => n2187, A2 => n5451, B1 => n2639, B2 => n5533
                           , ZN => n4658);
   U516 : OAI22_X1 port map( A1 => n2170, A2 => n5452, B1 => n2640, B2 => n5534
                           , ZN => n4640);
   U517 : OAI22_X1 port map( A1 => n2171, A2 => n5450, B1 => n2641, B2 => n5532
                           , ZN => n4622);
   U518 : OAI22_X1 port map( A1 => n2188, A2 => n5452, B1 => n2642, B2 => n5534
                           , ZN => n4604);
   U519 : OAI22_X1 port map( A1 => n2172, A2 => n5451, B1 => n2643, B2 => n5533
                           , ZN => n4586);
   U520 : OAI22_X1 port map( A1 => n2173, A2 => n5452, B1 => n2644, B2 => n5534
                           , ZN => n4568);
   U521 : OAI22_X1 port map( A1 => n2189, A2 => n5450, B1 => n2645, B2 => n5532
                           , ZN => n4550);
   U522 : OAI22_X1 port map( A1 => n2174, A2 => n5450, B1 => n2646, B2 => n5532
                           , ZN => n4532);
   U523 : OAI22_X1 port map( A1 => n2175, A2 => n5451, B1 => n2647, B2 => n5533
                           , ZN => n4497);
   U524 : OAI22_X1 port map( A1 => n2319, A2 => n5433, B1 => n2654, B2 => n5524
                           , ZN => n5098);
   U525 : OAI22_X1 port map( A1 => n2226, A2 => n5427, B1 => n2680, B2 => n5430
                           , ZN => n5099);
   U526 : OAI22_X1 port map( A1 => n2322, A2 => n5434, B1 => n2655, B2 => n5525
                           , ZN => n5056);
   U527 : OAI22_X1 port map( A1 => n2228, A2 => n5428, B1 => n2681, B2 => n5431
                           , ZN => n5057);
   U528 : OAI22_X1 port map( A1 => n2323, A2 => n5432, B1 => n2656, B2 => n5523
                           , ZN => n5038);
   U529 : OAI22_X1 port map( A1 => n2248, A2 => n5426, B1 => n2682, B2 => n5429
                           , ZN => n5039);
   U530 : OAI22_X1 port map( A1 => n2324, A2 => n5432, B1 => n2657, B2 => n5523
                           , ZN => n5020);
   U531 : OAI22_X1 port map( A1 => n2229, A2 => n5426, B1 => n2683, B2 => n5429
                           , ZN => n5021);
   U532 : OAI22_X1 port map( A1 => n2325, A2 => n5433, B1 => n2658, B2 => n5524
                           , ZN => n5002);
   U533 : OAI22_X1 port map( A1 => n2230, A2 => n5427, B1 => n2684, B2 => n5430
                           , ZN => n5003);
   U534 : OAI22_X1 port map( A1 => n2326, A2 => n5433, B1 => n2659, B2 => n5524
                           , ZN => n4984);
   U535 : OAI22_X1 port map( A1 => n2249, A2 => n5427, B1 => n2685, B2 => n5430
                           , ZN => n4985);
   U536 : OAI22_X1 port map( A1 => n2327, A2 => n5434, B1 => n2660, B2 => n5525
                           , ZN => n4966);
   U537 : OAI22_X1 port map( A1 => n2231, A2 => n5428, B1 => n2686, B2 => n5431
                           , ZN => n4967);
   U538 : OAI22_X1 port map( A1 => n2328, A2 => n5432, B1 => n2661, B2 => n5523
                           , ZN => n4948);
   U539 : OAI22_X1 port map( A1 => n2232, A2 => n5426, B1 => n2687, B2 => n5429
                           , ZN => n4949);
   U540 : OAI22_X1 port map( A1 => n2329, A2 => n5434, B1 => n2662, B2 => n5525
                           , ZN => n4930);
   U541 : OAI22_X1 port map( A1 => n2250, A2 => n5428, B1 => n2688, B2 => n5431
                           , ZN => n4931);
   U542 : OAI22_X1 port map( A1 => n2330, A2 => n5433, B1 => n2663, B2 => n5524
                           , ZN => n4912);
   U543 : OAI22_X1 port map( A1 => n2233, A2 => n5427, B1 => n2689, B2 => n5430
                           , ZN => n4913);
   U544 : OAI22_X1 port map( A1 => n2331, A2 => n5434, B1 => n2666, B2 => n5525
                           , ZN => n4894);
   U545 : OAI22_X1 port map( A1 => n2234, A2 => n5428, B1 => n2690, B2 => n5431
                           , ZN => n4895);
   U546 : OAI22_X1 port map( A1 => n2332, A2 => n5432, B1 => n2667, B2 => n5523
                           , ZN => n4876);
   U547 : OAI22_X1 port map( A1 => n2251, A2 => n5426, B1 => n2691, B2 => n5429
                           , ZN => n4877);
   U548 : OAI22_X1 port map( A1 => n2333, A2 => n5432, B1 => n2668, B2 => n5523
                           , ZN => n4858);
   U549 : OAI22_X1 port map( A1 => n2235, A2 => n5426, B1 => n2692, B2 => n5429
                           , ZN => n4859);
   U550 : OAI22_X1 port map( A1 => n2334, A2 => n5433, B1 => n2669, B2 => n5524
                           , ZN => n4840);
   U551 : OAI22_X1 port map( A1 => n2236, A2 => n5427, B1 => n2693, B2 => n5430
                           , ZN => n4841);
   U552 : OAI22_X1 port map( A1 => n2335, A2 => n5433, B1 => n2670, B2 => n5524
                           , ZN => n4822);
   U553 : OAI22_X1 port map( A1 => n2253, A2 => n5427, B1 => n2694, B2 => n5430
                           , ZN => n4823);
   U554 : OAI22_X1 port map( A1 => n2336, A2 => n5434, B1 => n2671, B2 => n5525
                           , ZN => n4804);
   U555 : OAI22_X1 port map( A1 => n2237, A2 => n5428, B1 => n2695, B2 => n5431
                           , ZN => n4805);
   U556 : OAI22_X1 port map( A1 => n2337, A2 => n5432, B1 => n2672, B2 => n5523
                           , ZN => n4786);
   U557 : OAI22_X1 port map( A1 => n2238, A2 => n5426, B1 => n2696, B2 => n5429
                           , ZN => n4787);
   U558 : OAI22_X1 port map( A1 => n2338, A2 => n5434, B1 => n2673, B2 => n5525
                           , ZN => n4768);
   U559 : OAI22_X1 port map( A1 => n2254, A2 => n5428, B1 => n2697, B2 => n5431
                           , ZN => n4769);
   U560 : OAI22_X1 port map( A1 => n2339, A2 => n5433, B1 => n2674, B2 => n5524
                           , ZN => n4750);
   U561 : OAI22_X1 port map( A1 => n2239, A2 => n5427, B1 => n2698, B2 => n5430
                           , ZN => n4751);
   U562 : OAI22_X1 port map( A1 => n2340, A2 => n5434, B1 => n2675, B2 => n5525
                           , ZN => n4732);
   U563 : OAI22_X1 port map( A1 => n2240, A2 => n5428, B1 => n2701, B2 => n5431
                           , ZN => n4733);
   U564 : OAI22_X1 port map( A1 => n2341, A2 => n5432, B1 => n2676, B2 => n5523
                           , ZN => n4714);
   U565 : OAI22_X1 port map( A1 => n2255, A2 => n5426, B1 => n2756, B2 => n5429
                           , ZN => n4715);
   U566 : OAI22_X1 port map( A1 => n2342, A2 => n5432, B1 => n2677, B2 => n5523
                           , ZN => n4696);
   U567 : OAI22_X1 port map( A1 => n2241, A2 => n5426, B1 => n2775, B2 => n5429
                           , ZN => n4697);
   U568 : OAI22_X1 port map( A1 => n2343, A2 => n5433, B1 => n2678, B2 => n5524
                           , ZN => n4678);
   U569 : OAI22_X1 port map( A1 => n2242, A2 => n5427, B1 => n2794, B2 => n5430
                           , ZN => n4679);
   U570 : OAI22_X1 port map( A1 => n2344, A2 => n5433, B1 => n2679, B2 => n5524
                           , ZN => n4660);
   U571 : OAI22_X1 port map( A1 => n2256, A2 => n5427, B1 => n2813, B2 => n5430
                           , ZN => n4661);
   U572 : OAI22_X1 port map( A1 => n2345, A2 => n5434, B1 => n2832, B2 => n5525
                           , ZN => n4642);
   U573 : OAI22_X1 port map( A1 => n2243, A2 => n5428, B1 => n2922, B2 => n5431
                           , ZN => n4643);
   U574 : OAI22_X1 port map( A1 => n2346, A2 => n5432, B1 => n2851, B2 => n5523
                           , ZN => n4624);
   U575 : OAI22_X1 port map( A1 => n2244, A2 => n5426, B1 => n2923, B2 => n5429
                           , ZN => n4625);
   U576 : OAI22_X1 port map( A1 => n2347, A2 => n5434, B1 => n2870, B2 => n5525
                           , ZN => n4606);
   U577 : OAI22_X1 port map( A1 => n2118, A2 => n5428, B1 => n2924, B2 => n5431
                           , ZN => n4607);
   U578 : OAI22_X1 port map( A1 => n2348, A2 => n5433, B1 => n2889, B2 => n5524
                           , ZN => n4588);
   U579 : OAI22_X1 port map( A1 => n2117, A2 => n5427, B1 => n2925, B2 => n5430
                           , ZN => n4589);
   U580 : OAI22_X1 port map( A1 => n2349, A2 => n5434, B1 => n2908, B2 => n5525
                           , ZN => n4570);
   U581 : OAI22_X1 port map( A1 => n2245, A2 => n5428, B1 => n2926, B2 => n5431
                           , ZN => n4571);
   U582 : OAI22_X1 port map( A1 => n2350, A2 => n5432, B1 => n2919, B2 => n5523
                           , ZN => n4552);
   U583 : OAI22_X1 port map( A1 => n2257, A2 => n5426, B1 => n2927, B2 => n5429
                           , ZN => n4553);
   U584 : OAI22_X1 port map( A1 => n2351, A2 => n5432, B1 => n2920, B2 => n5523
                           , ZN => n4534);
   U585 : OAI22_X1 port map( A1 => n2246, A2 => n5426, B1 => n2928, B2 => n5429
                           , ZN => n4535);
   U586 : OAI22_X1 port map( A1 => n2352, A2 => n5433, B1 => n2921, B2 => n5524
                           , ZN => n4510);
   U587 : OAI22_X1 port map( A1 => n2247, A2 => n5427, B1 => n2929, B2 => n5430
                           , ZN => n4515);
   U588 : OAI22_X1 port map( A1 => n4445, A2 => n2714, B1 => n5962, B2 => n5661
                           , ZN => n4444);
   U589 : NOR4_X1 port map( A1 => n4453, A2 => n4454, A3 => n4455, A4 => n4456,
                           ZN => n4445);
   U590 : OAI221_X1 port map( B1 => n5122, B2 => n5599, C1 => n2226, C2 => 
                           n5607, A => n4463, ZN => n4453);
   U591 : OAI221_X1 port map( B1 => n5123, B2 => n5630, C1 => n2227, C2 => 
                           n5470, A => n4462, ZN => n4454);
   U592 : OAI22_X1 port map( A1 => n5965, A2 => n5661, B1 => n2588, B2 => n5479
                           , ZN => n4415);
   U593 : OAI22_X1 port map( A1 => n5968, A2 => n5660, B1 => n2589, B2 => n5478
                           , ZN => n4393);
   U594 : OAI22_X1 port map( A1 => n5971, A2 => n5660, B1 => n2590, B2 => n5478
                           , ZN => n4374);
   U595 : OAI22_X1 port map( A1 => n5974, A2 => n5662, B1 => n2591, B2 => n5480
                           , ZN => n4355);
   U596 : OAI22_X1 port map( A1 => n5977, A2 => n5661, B1 => n2592, B2 => n5479
                           , ZN => n4336);
   U597 : OAI22_X1 port map( A1 => n5980, A2 => n5661, B1 => n2593, B2 => n5479
                           , ZN => n4317);
   U598 : OAI22_X1 port map( A1 => n5983, A2 => n5660, B1 => n2594, B2 => n5478
                           , ZN => n4298);
   U599 : OAI22_X1 port map( A1 => n5986, A2 => n5662, B1 => n2596, B2 => n5480
                           , ZN => n4279);
   U600 : OAI22_X1 port map( A1 => n5989, A2 => n5662, B1 => n2597, B2 => n5480
                           , ZN => n4260);
   U601 : OAI22_X1 port map( A1 => n5992, A2 => n5661, B1 => n2598, B2 => n5479
                           , ZN => n4241);
   U602 : OAI22_X1 port map( A1 => n5995, A2 => n5660, B1 => n2599, B2 => n5478
                           , ZN => n4222);
   U603 : OAI22_X1 port map( A1 => n5998, A2 => n5660, B1 => n2600, B2 => n5478
                           , ZN => n4203);
   U604 : OAI22_X1 port map( A1 => n6001, A2 => n5662, B1 => n2601, B2 => n5480
                           , ZN => n4184);
   U605 : OAI22_X1 port map( A1 => n6004, A2 => n5661, B1 => n2602, B2 => n5479
                           , ZN => n4165);
   U606 : OAI22_X1 port map( A1 => n6007, A2 => n5661, B1 => n2603, B2 => n5479
                           , ZN => n4146);
   U607 : OAI22_X1 port map( A1 => n6010, A2 => n5660, B1 => n2604, B2 => n5478
                           , ZN => n4127);
   U608 : OAI22_X1 port map( A1 => n6013, A2 => n5662, B1 => n2605, B2 => n5480
                           , ZN => n4108);
   U609 : OAI22_X1 port map( A1 => n6016, A2 => n5662, B1 => n2606, B2 => n5480
                           , ZN => n4089);
   U610 : OAI22_X1 port map( A1 => n6019, A2 => n5661, B1 => n2607, B2 => n5479
                           , ZN => n4070);
   U611 : OAI22_X1 port map( A1 => n6022, A2 => n5660, B1 => n2608, B2 => n5478
                           , ZN => n4051);
   U612 : OAI22_X1 port map( A1 => n6025, A2 => n5660, B1 => n2609, B2 => n5478
                           , ZN => n4032);
   U613 : OAI22_X1 port map( A1 => n6028, A2 => n5662, B1 => n2610, B2 => n5480
                           , ZN => n4013);
   U614 : OAI22_X1 port map( A1 => n6031, A2 => n5661, B1 => n2611, B2 => n5479
                           , ZN => n2907);
   U615 : OAI22_X1 port map( A1 => n6034, A2 => n5661, B1 => n2612, B2 => n5479
                           , ZN => n2888);
   U616 : OAI22_X1 port map( A1 => n6037, A2 => n5660, B1 => n2613, B2 => n5478
                           , ZN => n2869);
   U617 : OAI22_X1 port map( A1 => n6040, A2 => n5662, B1 => n2648, B2 => n5480
                           , ZN => n2850);
   U618 : OAI22_X1 port map( A1 => n6043, A2 => n5662, B1 => n2649, B2 => n5480
                           , ZN => n2831);
   U619 : OAI22_X1 port map( A1 => n6046, A2 => n5661, B1 => n2650, B2 => n5479
                           , ZN => n2812);
   U620 : OAI22_X1 port map( A1 => n6049, A2 => n5660, B1 => n2651, B2 => n5478
                           , ZN => n2793);
   U621 : OAI22_X1 port map( A1 => n6052, A2 => n5660, B1 => n2652, B2 => n5478
                           , ZN => n2774);
   U622 : OAI22_X1 port map( A1 => n6055, A2 => n5662, B1 => n2653, B2 => n5480
                           , ZN => n2753);
   U623 : OAI22_X1 port map( A1 => n2555, A2 => n5530, B1 => n2225, B2 => n5446
                           , ZN => n5092);
   U624 : OAI22_X1 port map( A1 => n2556, A2 => n5531, B1 => n2190, B2 => n5447
                           , ZN => n5053);
   U625 : OAI22_X1 port map( A1 => n2557, A2 => n5529, B1 => n2191, B2 => n5445
                           , ZN => n5035);
   U626 : OAI22_X1 port map( A1 => n2558, A2 => n5529, B1 => n2192, B2 => n5445
                           , ZN => n5017);
   U627 : OAI22_X1 port map( A1 => n2559, A2 => n5530, B1 => n2193, B2 => n5446
                           , ZN => n4999);
   U628 : OAI22_X1 port map( A1 => n2560, A2 => n5530, B1 => n2194, B2 => n5446
                           , ZN => n4981);
   U629 : OAI22_X1 port map( A1 => n2562, A2 => n5531, B1 => n2195, B2 => n5447
                           , ZN => n4963);
   U630 : OAI22_X1 port map( A1 => n2563, A2 => n5529, B1 => n2196, B2 => n5445
                           , ZN => n4945);
   U631 : OAI22_X1 port map( A1 => n2564, A2 => n5531, B1 => n2197, B2 => n5447
                           , ZN => n4927);
   U632 : OAI22_X1 port map( A1 => n2565, A2 => n5530, B1 => n2198, B2 => n5446
                           , ZN => n4909);
   U633 : OAI22_X1 port map( A1 => n2566, A2 => n5531, B1 => n2199, B2 => n5447
                           , ZN => n4891);
   U634 : OAI22_X1 port map( A1 => n2567, A2 => n5529, B1 => n2200, B2 => n5445
                           , ZN => n4873);
   U635 : OAI22_X1 port map( A1 => n2568, A2 => n5529, B1 => n2201, B2 => n5445
                           , ZN => n4855);
   U636 : OAI22_X1 port map( A1 => n2569, A2 => n5530, B1 => n2202, B2 => n5446
                           , ZN => n4837);
   U637 : OAI22_X1 port map( A1 => n2570, A2 => n5530, B1 => n2203, B2 => n5446
                           , ZN => n4819);
   U638 : OAI22_X1 port map( A1 => n2571, A2 => n5531, B1 => n2204, B2 => n5447
                           , ZN => n4801);
   U639 : OAI22_X1 port map( A1 => n2572, A2 => n5529, B1 => n2205, B2 => n5445
                           , ZN => n4783);
   U640 : OAI22_X1 port map( A1 => n2573, A2 => n5531, B1 => n2206, B2 => n5447
                           , ZN => n4765);
   U641 : OAI22_X1 port map( A1 => n2574, A2 => n5530, B1 => n2207, B2 => n5446
                           , ZN => n4747);
   U642 : OAI22_X1 port map( A1 => n2575, A2 => n5531, B1 => n2208, B2 => n5447
                           , ZN => n4729);
   U643 : OAI22_X1 port map( A1 => n2576, A2 => n5529, B1 => n2209, B2 => n5445
                           , ZN => n4711);
   U644 : OAI22_X1 port map( A1 => n2577, A2 => n5529, B1 => n2210, B2 => n5445
                           , ZN => n4693);
   U645 : OAI22_X1 port map( A1 => n2578, A2 => n5530, B1 => n2211, B2 => n5446
                           , ZN => n4675);
   U646 : OAI22_X1 port map( A1 => n2579, A2 => n5530, B1 => n2212, B2 => n5446
                           , ZN => n4657);
   U647 : OAI22_X1 port map( A1 => n2580, A2 => n5531, B1 => n2213, B2 => n5447
                           , ZN => n4639);
   U648 : OAI22_X1 port map( A1 => n2581, A2 => n5529, B1 => n2214, B2 => n5445
                           , ZN => n4621);
   U649 : OAI22_X1 port map( A1 => n2582, A2 => n5531, B1 => n2215, B2 => n5447
                           , ZN => n4603);
   U650 : OAI22_X1 port map( A1 => n2583, A2 => n5530, B1 => n2216, B2 => n5446
                           , ZN => n4585);
   U651 : OAI22_X1 port map( A1 => n2584, A2 => n5531, B1 => n2219, B2 => n5447
                           , ZN => n4567);
   U652 : OAI22_X1 port map( A1 => n2585, A2 => n5529, B1 => n2220, B2 => n5445
                           , ZN => n4549);
   U653 : OAI22_X1 port map( A1 => n2586, A2 => n5529, B1 => n2221, B2 => n5445
                           , ZN => n4531);
   U654 : OAI22_X1 port map( A1 => n2587, A2 => n5530, B1 => n2222, B2 => n5446
                           , ZN => n4496);
   U655 : NAND4_X1 port map( A1 => n4447, A2 => n4465, A3 => n4446, A4 => n4466
                           , ZN => n4464);
   U656 : NOR3_X1 port map( A1 => n4451, A2 => n2182, A3 => n4450, ZN => n4466)
                           ;
   U657 : INV_X1 port map( A => n4452, ZN => n4465);
   U658 : NAND4_X1 port map( A1 => n5085, A2 => n5506, A3 => n5090, A4 => n5095
                           , ZN => n4507);
   U659 : BUF_X1 port map( A => n1692, Z => n5962);
   U660 : BUF_X1 port map( A => n1690, Z => n5965);
   U661 : BUF_X1 port map( A => n1688, Z => n5968);
   U662 : BUF_X1 port map( A => n1686, Z => n5971);
   U663 : BUF_X1 port map( A => n1684, Z => n5974);
   U664 : BUF_X1 port map( A => n1682, Z => n5977);
   U665 : BUF_X1 port map( A => n1680, Z => n5980);
   U666 : BUF_X1 port map( A => n1678, Z => n5983);
   U667 : BUF_X1 port map( A => n1676, Z => n5986);
   U668 : BUF_X1 port map( A => n1674, Z => n5989);
   U669 : BUF_X1 port map( A => n1672, Z => n5992);
   U670 : BUF_X1 port map( A => n1670, Z => n5995);
   U671 : BUF_X1 port map( A => n1668, Z => n5998);
   U672 : BUF_X1 port map( A => n1666, Z => n6001);
   U673 : BUF_X1 port map( A => n1664, Z => n6004);
   U674 : BUF_X1 port map( A => n1662, Z => n6007);
   U675 : BUF_X1 port map( A => n1660, Z => n6010);
   U676 : BUF_X1 port map( A => n1658, Z => n6013);
   U677 : BUF_X1 port map( A => n1656, Z => n6016);
   U678 : BUF_X1 port map( A => n1654, Z => n6019);
   U679 : BUF_X1 port map( A => n1652, Z => n6022);
   U680 : BUF_X1 port map( A => n1650, Z => n6025);
   U681 : BUF_X1 port map( A => n1648, Z => n6028);
   U682 : BUF_X1 port map( A => n1646, Z => n6031);
   U683 : BUF_X1 port map( A => n1644, Z => n6034);
   U684 : BUF_X1 port map( A => n1642, Z => n6037);
   U685 : BUF_X1 port map( A => n1640, Z => n6040);
   U686 : BUF_X1 port map( A => n1638, Z => n6043);
   U687 : BUF_X1 port map( A => n1636, Z => n6046);
   U688 : BUF_X1 port map( A => n1634, Z => n6049);
   U689 : BUF_X1 port map( A => n1632, Z => n6052);
   U690 : BUF_X1 port map( A => n1629, Z => n6055);
   U691 : BUF_X1 port map( A => n1692, Z => n5963);
   U692 : BUF_X1 port map( A => n1690, Z => n5966);
   U693 : BUF_X1 port map( A => n1688, Z => n5969);
   U694 : BUF_X1 port map( A => n1686, Z => n5972);
   U695 : BUF_X1 port map( A => n1684, Z => n5975);
   U696 : BUF_X1 port map( A => n1682, Z => n5978);
   U697 : BUF_X1 port map( A => n1680, Z => n5981);
   U698 : BUF_X1 port map( A => n1678, Z => n5984);
   U699 : BUF_X1 port map( A => n1676, Z => n5987);
   U700 : BUF_X1 port map( A => n1674, Z => n5990);
   U701 : BUF_X1 port map( A => n1672, Z => n5993);
   U702 : BUF_X1 port map( A => n1670, Z => n5996);
   U703 : BUF_X1 port map( A => n1668, Z => n5999);
   U704 : BUF_X1 port map( A => n1666, Z => n6002);
   U705 : BUF_X1 port map( A => n1664, Z => n6005);
   U706 : BUF_X1 port map( A => n1662, Z => n6008);
   U707 : BUF_X1 port map( A => n1660, Z => n6011);
   U708 : BUF_X1 port map( A => n1658, Z => n6014);
   U709 : BUF_X1 port map( A => n1656, Z => n6017);
   U710 : BUF_X1 port map( A => n1654, Z => n6020);
   U711 : BUF_X1 port map( A => n1652, Z => n6023);
   U712 : BUF_X1 port map( A => n1650, Z => n6026);
   U713 : BUF_X1 port map( A => n1648, Z => n6029);
   U714 : BUF_X1 port map( A => n1646, Z => n6032);
   U715 : BUF_X1 port map( A => n1644, Z => n6035);
   U716 : BUF_X1 port map( A => n1642, Z => n6038);
   U717 : BUF_X1 port map( A => n1640, Z => n6041);
   U718 : BUF_X1 port map( A => n1638, Z => n6044);
   U719 : BUF_X1 port map( A => n1636, Z => n6047);
   U720 : BUF_X1 port map( A => n1634, Z => n6050);
   U721 : BUF_X1 port map( A => n1632, Z => n6053);
   U722 : BUF_X1 port map( A => n1629, Z => n6056);
   U723 : NAND2_X1 port map( A1 => n1730, A2 => n1695, ZN => n1698);
   U724 : NAND2_X1 port map( A1 => n1694, A2 => n1695, ZN => n1628);
   U725 : NAND2_X1 port map( A1 => n1803, A2 => n1804, ZN => n1769);
   U726 : OAI22_X1 port map( A1 => n5966, A2 => n5837, B1 => n5390, B2 => n2588
                           , ZN => n3528);
   U727 : OAI22_X1 port map( A1 => n5969, A2 => n5842, B1 => n5390, B2 => n2589
                           , ZN => n3529);
   U728 : OAI22_X1 port map( A1 => n5972, A2 => n5836, B1 => n5390, B2 => n2590
                           , ZN => n3530);
   U729 : OAI22_X1 port map( A1 => n5975, A2 => n5837, B1 => n5390, B2 => n2591
                           , ZN => n3531);
   U730 : OAI22_X1 port map( A1 => n5978, A2 => n5841, B1 => n5390, B2 => n2592
                           , ZN => n3532);
   U731 : OAI22_X1 port map( A1 => n5981, A2 => n5839, B1 => n5390, B2 => n2593
                           , ZN => n3533);
   U732 : OAI22_X1 port map( A1 => n5984, A2 => n5838, B1 => n5390, B2 => n2594
                           , ZN => n3534);
   U733 : OAI22_X1 port map( A1 => n5987, A2 => n5838, B1 => n5390, B2 => n2596
                           , ZN => n3535);
   U734 : OAI22_X1 port map( A1 => n5990, A2 => n5838, B1 => n5390, B2 => n2597
                           , ZN => n3536);
   U735 : OAI22_X1 port map( A1 => n5993, A2 => n5837, B1 => n5390, B2 => n2598
                           , ZN => n3537);
   U736 : OAI22_X1 port map( A1 => n5996, A2 => n5839, B1 => n5390, B2 => n2599
                           , ZN => n3538);
   U737 : OAI22_X1 port map( A1 => n5999, A2 => n5838, B1 => n5390, B2 => n2600
                           , ZN => n3539);
   U738 : OAI22_X1 port map( A1 => n5967, A2 => n5927, B1 => n5420, B2 => n2523
                           , ZN => n3848);
   U739 : OAI22_X1 port map( A1 => n5970, A2 => n5931, B1 => n5420, B2 => n2524
                           , ZN => n3849);
   U740 : OAI22_X1 port map( A1 => n5973, A2 => n5926, B1 => n5420, B2 => n2525
                           , ZN => n3850);
   U741 : OAI22_X1 port map( A1 => n5976, A2 => n5927, B1 => n5420, B2 => n2526
                           , ZN => n3851);
   U742 : OAI22_X1 port map( A1 => n5979, A2 => n5931, B1 => n5420, B2 => n2528
                           , ZN => n3852);
   U743 : OAI22_X1 port map( A1 => n5982, A2 => n5929, B1 => n5420, B2 => n2529
                           , ZN => n3853);
   U744 : OAI22_X1 port map( A1 => n5985, A2 => n5927, B1 => n5420, B2 => n2530
                           , ZN => n3854);
   U745 : OAI22_X1 port map( A1 => n5988, A2 => n5928, B1 => n5420, B2 => n2531
                           , ZN => n3855);
   U746 : OAI22_X1 port map( A1 => n5991, A2 => n5928, B1 => n5420, B2 => n2532
                           , ZN => n3856);
   U747 : OAI22_X1 port map( A1 => n5994, A2 => n5927, B1 => n5420, B2 => n2533
                           , ZN => n3857);
   U748 : OAI22_X1 port map( A1 => n5997, A2 => n5929, B1 => n5420, B2 => n2534
                           , ZN => n3858);
   U749 : OAI22_X1 port map( A1 => n6000, A2 => n5927, B1 => n5420, B2 => n2535
                           , ZN => n3859);
   U750 : OAI22_X1 port map( A1 => n6002, A2 => n5838, B1 => n5391, B2 => n2601
                           , ZN => n3540);
   U751 : OAI22_X1 port map( A1 => n6005, A2 => n5838, B1 => n5391, B2 => n2602
                           , ZN => n3541);
   U752 : OAI22_X1 port map( A1 => n6008, A2 => n5840, B1 => n5391, B2 => n2603
                           , ZN => n3542);
   U753 : OAI22_X1 port map( A1 => n6011, A2 => n5839, B1 => n5391, B2 => n2604
                           , ZN => n3543);
   U754 : OAI22_X1 port map( A1 => n6014, A2 => n5840, B1 => n5391, B2 => n2605
                           , ZN => n3544);
   U755 : OAI22_X1 port map( A1 => n6017, A2 => n5840, B1 => n5391, B2 => n2606
                           , ZN => n3545);
   U756 : OAI22_X1 port map( A1 => n6020, A2 => n5837, B1 => n5391, B2 => n2607
                           , ZN => n3546);
   U757 : OAI22_X1 port map( A1 => n6023, A2 => n5836, B1 => n5391, B2 => n2608
                           , ZN => n3547);
   U758 : OAI22_X1 port map( A1 => n6026, A2 => n5840, B1 => n5391, B2 => n2609
                           , ZN => n3548);
   U759 : OAI22_X1 port map( A1 => n6029, A2 => n5839, B1 => n5391, B2 => n2610
                           , ZN => n3549);
   U760 : OAI22_X1 port map( A1 => n6032, A2 => n5842, B1 => n5391, B2 => n2611
                           , ZN => n3550);
   U761 : OAI22_X1 port map( A1 => n6035, A2 => n5841, B1 => n5391, B2 => n2612
                           , ZN => n3551);
   U762 : OAI22_X1 port map( A1 => n6038, A2 => n5842, B1 => n5391, B2 => n2613
                           , ZN => n3552);
   U763 : OAI22_X1 port map( A1 => n6003, A2 => n5928, B1 => n5421, B2 => n2536
                           , ZN => n3860);
   U764 : OAI22_X1 port map( A1 => n6006, A2 => n5927, B1 => n5421, B2 => n2537
                           , ZN => n3861);
   U765 : OAI22_X1 port map( A1 => n6009, A2 => n5930, B1 => n5421, B2 => n2538
                           , ZN => n3862);
   U766 : OAI22_X1 port map( A1 => n6012, A2 => n5929, B1 => n5421, B2 => n2539
                           , ZN => n3863);
   U767 : OAI22_X1 port map( A1 => n6015, A2 => n5930, B1 => n5421, B2 => n2540
                           , ZN => n3864);
   U768 : OAI22_X1 port map( A1 => n6018, A2 => n5929, B1 => n5421, B2 => n2541
                           , ZN => n3865);
   U769 : OAI22_X1 port map( A1 => n6021, A2 => n5927, B1 => n5421, B2 => n2542
                           , ZN => n3866);
   U770 : OAI22_X1 port map( A1 => n6024, A2 => n5926, B1 => n5421, B2 => n2543
                           , ZN => n3867);
   U771 : OAI22_X1 port map( A1 => n6027, A2 => n5930, B1 => n5421, B2 => n2544
                           , ZN => n3868);
   U772 : OAI22_X1 port map( A1 => n6030, A2 => n5930, B1 => n5421, B2 => n2547
                           , ZN => n3869);
   U773 : OAI22_X1 port map( A1 => n6033, A2 => n5932, B1 => n5421, B2 => n2548
                           , ZN => n3870);
   U774 : OAI22_X1 port map( A1 => n6036, A2 => n5931, B1 => n5421, B2 => n2549
                           , ZN => n3871);
   U775 : OAI22_X1 port map( A1 => n6039, A2 => n5932, B1 => n5421, B2 => n2550
                           , ZN => n3872);
   U776 : OAI22_X1 port map( A1 => n5962, A2 => n5703, B1 => n5345, B2 => n5312
                           , ZN => n3047);
   U777 : OAI22_X1 port map( A1 => n5965, A2 => n5701, B1 => n5345, B2 => n5280
                           , ZN => n3048);
   U778 : OAI22_X1 port map( A1 => n5968, A2 => n5703, B1 => n5345, B2 => n5281
                           , ZN => n3049);
   U779 : OAI22_X1 port map( A1 => n5971, A2 => n5702, B1 => n5345, B2 => n5282
                           , ZN => n3050);
   U780 : OAI22_X1 port map( A1 => n5974, A2 => n5701, B1 => n5345, B2 => n5283
                           , ZN => n3051);
   U781 : OAI22_X1 port map( A1 => n5977, A2 => n5706, B1 => n5345, B2 => n5284
                           , ZN => n3052);
   U782 : OAI22_X1 port map( A1 => n5980, A2 => n5702, B1 => n5345, B2 => n5285
                           , ZN => n3053);
   U783 : OAI22_X1 port map( A1 => n5983, A2 => n5703, B1 => n5345, B2 => n5286
                           , ZN => n3054);
   U784 : OAI22_X1 port map( A1 => n5986, A2 => n5703, B1 => n5345, B2 => n5299
                           , ZN => n3055);
   U785 : OAI22_X1 port map( A1 => n5989, A2 => n5706, B1 => n5345, B2 => n5287
                           , ZN => n3056);
   U786 : OAI22_X1 port map( A1 => n5992, A2 => n5704, B1 => n5345, B2 => n5288
                           , ZN => n3057);
   U787 : OAI22_X1 port map( A1 => n5995, A2 => n5705, B1 => n5345, B2 => n5289
                           , ZN => n3058);
   U788 : OAI22_X1 port map( A1 => n5998, A2 => n5702, B1 => n5346, B2 => n5290
                           , ZN => n3059);
   U789 : OAI22_X1 port map( A1 => n6001, A2 => n5703, B1 => n5346, B2 => n5291
                           , ZN => n3060);
   U790 : OAI22_X1 port map( A1 => n6004, A2 => n5702, B1 => n5346, B2 => n5292
                           , ZN => n3061);
   U791 : OAI22_X1 port map( A1 => n6007, A2 => n5707, B1 => n5346, B2 => n5293
                           , ZN => n3062);
   U792 : OAI22_X1 port map( A1 => n6010, A2 => n5704, B1 => n5346, B2 => n5294
                           , ZN => n3063);
   U793 : OAI22_X1 port map( A1 => n6013, A2 => n5705, B1 => n5346, B2 => n5308
                           , ZN => n3064);
   U794 : OAI22_X1 port map( A1 => n6016, A2 => n5705, B1 => n5346, B2 => n5295
                           , ZN => n3065);
   U795 : OAI22_X1 port map( A1 => n6019, A2 => n5701, B1 => n5346, B2 => n5296
                           , ZN => n3066);
   U796 : OAI22_X1 port map( A1 => n6022, A2 => n5704, B1 => n5346, B2 => n5300
                           , ZN => n3067);
   U797 : OAI22_X1 port map( A1 => n6025, A2 => n5707, B1 => n5346, B2 => n5301
                           , ZN => n3068);
   U798 : OAI22_X1 port map( A1 => n6028, A2 => n5706, B1 => n5346, B2 => n5302
                           , ZN => n3069);
   U799 : OAI22_X1 port map( A1 => n6031, A2 => n5707, B1 => n5346, B2 => n5303
                           , ZN => n3070);
   U800 : OAI22_X1 port map( A1 => n5962, A2 => n5712, B1 => n5348, B2 => n2654
                           , ZN => n3079);
   U801 : OAI22_X1 port map( A1 => n5965, A2 => n5710, B1 => n5348, B2 => n2655
                           , ZN => n3080);
   U802 : OAI22_X1 port map( A1 => n5968, A2 => n5712, B1 => n5348, B2 => n2656
                           , ZN => n3081);
   U803 : OAI22_X1 port map( A1 => n5971, A2 => n5711, B1 => n5348, B2 => n2657
                           , ZN => n3082);
   U804 : OAI22_X1 port map( A1 => n5974, A2 => n5710, B1 => n5348, B2 => n2658
                           , ZN => n3083);
   U805 : OAI22_X1 port map( A1 => n5977, A2 => n5715, B1 => n5348, B2 => n2659
                           , ZN => n3084);
   U806 : OAI22_X1 port map( A1 => n5980, A2 => n5711, B1 => n5348, B2 => n2660
                           , ZN => n3085);
   U807 : OAI22_X1 port map( A1 => n5983, A2 => n5712, B1 => n5348, B2 => n2661
                           , ZN => n3086);
   U808 : OAI22_X1 port map( A1 => n5986, A2 => n5712, B1 => n5348, B2 => n2662
                           , ZN => n3087);
   U809 : OAI22_X1 port map( A1 => n5989, A2 => n5715, B1 => n5348, B2 => n2663
                           , ZN => n3088);
   U810 : OAI22_X1 port map( A1 => n5992, A2 => n5713, B1 => n5348, B2 => n2666
                           , ZN => n3089);
   U811 : OAI22_X1 port map( A1 => n5995, A2 => n5714, B1 => n5348, B2 => n2667
                           , ZN => n3090);
   U812 : OAI22_X1 port map( A1 => n5998, A2 => n5711, B1 => n5349, B2 => n2668
                           , ZN => n3091);
   U813 : OAI22_X1 port map( A1 => n6001, A2 => n5712, B1 => n5349, B2 => n2669
                           , ZN => n3092);
   U814 : OAI22_X1 port map( A1 => n6004, A2 => n5711, B1 => n5349, B2 => n2670
                           , ZN => n3093);
   U815 : OAI22_X1 port map( A1 => n6007, A2 => n5716, B1 => n5349, B2 => n2671
                           , ZN => n3094);
   U816 : OAI22_X1 port map( A1 => n6010, A2 => n5713, B1 => n5349, B2 => n2672
                           , ZN => n3095);
   U817 : OAI22_X1 port map( A1 => n6013, A2 => n5714, B1 => n5349, B2 => n2673
                           , ZN => n3096);
   U818 : OAI22_X1 port map( A1 => n6016, A2 => n5714, B1 => n5349, B2 => n2674
                           , ZN => n3097);
   U819 : OAI22_X1 port map( A1 => n6019, A2 => n5710, B1 => n5349, B2 => n2675
                           , ZN => n3098);
   U820 : OAI22_X1 port map( A1 => n6022, A2 => n5713, B1 => n5349, B2 => n2676
                           , ZN => n3099);
   U821 : OAI22_X1 port map( A1 => n6025, A2 => n5716, B1 => n5349, B2 => n2677
                           , ZN => n3100);
   U822 : OAI22_X1 port map( A1 => n6028, A2 => n5715, B1 => n5349, B2 => n2678
                           , ZN => n3101);
   U823 : OAI22_X1 port map( A1 => n6031, A2 => n5716, B1 => n5349, B2 => n2679
                           , ZN => n3102);
   U824 : OAI22_X1 port map( A1 => n5962, A2 => n5721, B1 => n5351, B2 => n2614
                           , ZN => n3111);
   U825 : OAI22_X1 port map( A1 => n5965, A2 => n5719, B1 => n5351, B2 => n2615
                           , ZN => n3112);
   U826 : OAI22_X1 port map( A1 => n5968, A2 => n5721, B1 => n5351, B2 => n2616
                           , ZN => n3113);
   U827 : OAI22_X1 port map( A1 => n5971, A2 => n5720, B1 => n5351, B2 => n2617
                           , ZN => n3114);
   U828 : OAI22_X1 port map( A1 => n5974, A2 => n5719, B1 => n5351, B2 => n2618
                           , ZN => n3115);
   U829 : OAI22_X1 port map( A1 => n5977, A2 => n5724, B1 => n5351, B2 => n2619
                           , ZN => n3116);
   U830 : OAI22_X1 port map( A1 => n5980, A2 => n5720, B1 => n5351, B2 => n2620
                           , ZN => n3117);
   U831 : OAI22_X1 port map( A1 => n5983, A2 => n5721, B1 => n5351, B2 => n2621
                           , ZN => n3118);
   U832 : OAI22_X1 port map( A1 => n5986, A2 => n5721, B1 => n5351, B2 => n2622
                           , ZN => n3119);
   U833 : OAI22_X1 port map( A1 => n5989, A2 => n5724, B1 => n5351, B2 => n2623
                           , ZN => n3120);
   U834 : OAI22_X1 port map( A1 => n5992, A2 => n5722, B1 => n5351, B2 => n2624
                           , ZN => n3121);
   U835 : OAI22_X1 port map( A1 => n5995, A2 => n5723, B1 => n5351, B2 => n2625
                           , ZN => n3122);
   U836 : OAI22_X1 port map( A1 => n5998, A2 => n5720, B1 => n5352, B2 => n2626
                           , ZN => n3123);
   U837 : OAI22_X1 port map( A1 => n6001, A2 => n5721, B1 => n5352, B2 => n2627
                           , ZN => n3124);
   U838 : OAI22_X1 port map( A1 => n6004, A2 => n5720, B1 => n5352, B2 => n2628
                           , ZN => n3125);
   U839 : OAI22_X1 port map( A1 => n6007, A2 => n5725, B1 => n5352, B2 => n2631
                           , ZN => n3126);
   U840 : OAI22_X1 port map( A1 => n6010, A2 => n5722, B1 => n5352, B2 => n2632
                           , ZN => n3127);
   U841 : OAI22_X1 port map( A1 => n6013, A2 => n5723, B1 => n5352, B2 => n2633
                           , ZN => n3128);
   U842 : OAI22_X1 port map( A1 => n6016, A2 => n5723, B1 => n5352, B2 => n2634
                           , ZN => n3129);
   U843 : OAI22_X1 port map( A1 => n6019, A2 => n5719, B1 => n5352, B2 => n2635
                           , ZN => n3130);
   U844 : OAI22_X1 port map( A1 => n6022, A2 => n5722, B1 => n5352, B2 => n2636
                           , ZN => n3131);
   U845 : OAI22_X1 port map( A1 => n6025, A2 => n5725, B1 => n5352, B2 => n2637
                           , ZN => n3132);
   U846 : OAI22_X1 port map( A1 => n6028, A2 => n5724, B1 => n5352, B2 => n2638
                           , ZN => n3133);
   U847 : OAI22_X1 port map( A1 => n6031, A2 => n5725, B1 => n5352, B2 => n2639
                           , ZN => n3134);
   U848 : OAI22_X1 port map( A1 => n5962, A2 => n5729, B1 => n5354, B2 => n2116
                           , ZN => n3143);
   U849 : OAI22_X1 port map( A1 => n5965, A2 => n5728, B1 => n5354, B2 => n2353
                           , ZN => n3144);
   U850 : OAI22_X1 port map( A1 => n5968, A2 => n5729, B1 => n5354, B2 => n2354
                           , ZN => n3145);
   U851 : OAI22_X1 port map( A1 => n5971, A2 => n5731, B1 => n5354, B2 => n2357
                           , ZN => n3146);
   U852 : OAI22_X1 port map( A1 => n5974, A2 => n5729, B1 => n5354, B2 => n2358
                           , ZN => n3147);
   U853 : OAI22_X1 port map( A1 => n5977, A2 => n5734, B1 => n5354, B2 => n2359
                           , ZN => n3148);
   U854 : OAI22_X1 port map( A1 => n5980, A2 => n5730, B1 => n5354, B2 => n2360
                           , ZN => n3149);
   U855 : OAI22_X1 port map( A1 => n5983, A2 => n5731, B1 => n5354, B2 => n2361
                           , ZN => n3150);
   U856 : OAI22_X1 port map( A1 => n5986, A2 => n5731, B1 => n5354, B2 => n2374
                           , ZN => n3151);
   U857 : OAI22_X1 port map( A1 => n5989, A2 => n5733, B1 => n5354, B2 => n2362
                           , ZN => n3152);
   U858 : OAI22_X1 port map( A1 => n5992, A2 => n5733, B1 => n5354, B2 => n2363
                           , ZN => n3153);
   U859 : OAI22_X1 port map( A1 => n5995, A2 => n5732, B1 => n5354, B2 => n2364
                           , ZN => n3154);
   U860 : OAI22_X1 port map( A1 => n5998, A2 => n5730, B1 => n5355, B2 => n2365
                           , ZN => n3155);
   U861 : OAI22_X1 port map( A1 => n6001, A2 => n5731, B1 => n5355, B2 => n2366
                           , ZN => n3156);
   U862 : OAI22_X1 port map( A1 => n6004, A2 => n5730, B1 => n5355, B2 => n2367
                           , ZN => n3157);
   U863 : OAI22_X1 port map( A1 => n6007, A2 => n5732, B1 => n5355, B2 => n2368
                           , ZN => n3158);
   U864 : OAI22_X1 port map( A1 => n6010, A2 => n5732, B1 => n5355, B2 => n2369
                           , ZN => n3159);
   U865 : OAI22_X1 port map( A1 => n6013, A2 => n5732, B1 => n5355, B2 => n2383
                           , ZN => n3160);
   U866 : OAI22_X1 port map( A1 => n6016, A2 => n5733, B1 => n5355, B2 => n2370
                           , ZN => n3161);
   U867 : OAI22_X1 port map( A1 => n6019, A2 => n5729, B1 => n5355, B2 => n2371
                           , ZN => n3162);
   U868 : OAI22_X1 port map( A1 => n6022, A2 => n5733, B1 => n5355, B2 => n2375
                           , ZN => n3163);
   U869 : OAI22_X1 port map( A1 => n6025, A2 => n5732, B1 => n5355, B2 => n2376
                           , ZN => n3164);
   U870 : OAI22_X1 port map( A1 => n6028, A2 => n5733, B1 => n5355, B2 => n2377
                           , ZN => n3165);
   U871 : OAI22_X1 port map( A1 => n6031, A2 => n5734, B1 => n5355, B2 => n2378
                           , ZN => n3166);
   U872 : OAI22_X1 port map( A1 => n5963, A2 => n5738, B1 => n5357, B2 => n5279
                           , ZN => n3175);
   U873 : OAI22_X1 port map( A1 => n5966, A2 => n5737, B1 => n5357, B2 => n2455
                           , ZN => n3176);
   U874 : OAI22_X1 port map( A1 => n5969, A2 => n5738, B1 => n5357, B2 => n2456
                           , ZN => n3177);
   U875 : OAI22_X1 port map( A1 => n5972, A2 => n5740, B1 => n5357, B2 => n2457
                           , ZN => n3178);
   U876 : OAI22_X1 port map( A1 => n5975, A2 => n5738, B1 => n5357, B2 => n2459
                           , ZN => n3179);
   U877 : OAI22_X1 port map( A1 => n5978, A2 => n5743, B1 => n5357, B2 => n2460
                           , ZN => n3180);
   U878 : OAI22_X1 port map( A1 => n5981, A2 => n5739, B1 => n5357, B2 => n2461
                           , ZN => n3181);
   U879 : OAI22_X1 port map( A1 => n5984, A2 => n5740, B1 => n5357, B2 => n2462
                           , ZN => n3182);
   U880 : OAI22_X1 port map( A1 => n5987, A2 => n5740, B1 => n5357, B2 => n2463
                           , ZN => n3183);
   U881 : OAI22_X1 port map( A1 => n5990, A2 => n5742, B1 => n5357, B2 => n2464
                           , ZN => n3184);
   U882 : OAI22_X1 port map( A1 => n5993, A2 => n5742, B1 => n5357, B2 => n2465
                           , ZN => n3185);
   U883 : OAI22_X1 port map( A1 => n5996, A2 => n5741, B1 => n5357, B2 => n2466
                           , ZN => n3186);
   U884 : OAI22_X1 port map( A1 => n5999, A2 => n5739, B1 => n5358, B2 => n2467
                           , ZN => n3187);
   U885 : OAI22_X1 port map( A1 => n6002, A2 => n5740, B1 => n5358, B2 => n2468
                           , ZN => n3188);
   U886 : OAI22_X1 port map( A1 => n6005, A2 => n5739, B1 => n5358, B2 => n2469
                           , ZN => n3189);
   U887 : OAI22_X1 port map( A1 => n6008, A2 => n5741, B1 => n5358, B2 => n2470
                           , ZN => n3190);
   U888 : OAI22_X1 port map( A1 => n6011, A2 => n5741, B1 => n5358, B2 => n2471
                           , ZN => n3191);
   U889 : OAI22_X1 port map( A1 => n6014, A2 => n5741, B1 => n5358, B2 => n2472
                           , ZN => n3192);
   U890 : OAI22_X1 port map( A1 => n6017, A2 => n5742, B1 => n5358, B2 => n2473
                           , ZN => n3193);
   U891 : OAI22_X1 port map( A1 => n6020, A2 => n5738, B1 => n5358, B2 => n2474
                           , ZN => n3194);
   U892 : OAI22_X1 port map( A1 => n6023, A2 => n5742, B1 => n5358, B2 => n2475
                           , ZN => n3195);
   U893 : OAI22_X1 port map( A1 => n6026, A2 => n5741, B1 => n5358, B2 => n2476
                           , ZN => n3196);
   U894 : OAI22_X1 port map( A1 => n6029, A2 => n5742, B1 => n5358, B2 => n2477
                           , ZN => n3197);
   U895 : OAI22_X1 port map( A1 => n6032, A2 => n5743, B1 => n5358, B2 => n2478
                           , ZN => n3198);
   U896 : OAI22_X1 port map( A1 => n5962, A2 => n5748, B1 => n5360, B2 => n2555
                           , ZN => n3207);
   U897 : OAI22_X1 port map( A1 => n5965, A2 => n5746, B1 => n5360, B2 => n2556
                           , ZN => n3208);
   U898 : OAI22_X1 port map( A1 => n5968, A2 => n5748, B1 => n5360, B2 => n2557
                           , ZN => n3209);
   U899 : OAI22_X1 port map( A1 => n5971, A2 => n5747, B1 => n5360, B2 => n2558
                           , ZN => n3210);
   U900 : OAI22_X1 port map( A1 => n5974, A2 => n5746, B1 => n5360, B2 => n2559
                           , ZN => n3211);
   U901 : OAI22_X1 port map( A1 => n5977, A2 => n5751, B1 => n5360, B2 => n2560
                           , ZN => n3212);
   U902 : OAI22_X1 port map( A1 => n5980, A2 => n5747, B1 => n5360, B2 => n2562
                           , ZN => n3213);
   U903 : OAI22_X1 port map( A1 => n5983, A2 => n5748, B1 => n5360, B2 => n2563
                           , ZN => n3214);
   U904 : OAI22_X1 port map( A1 => n5986, A2 => n5748, B1 => n5360, B2 => n2564
                           , ZN => n3215);
   U905 : OAI22_X1 port map( A1 => n5989, A2 => n5751, B1 => n5360, B2 => n2565
                           , ZN => n3216);
   U906 : OAI22_X1 port map( A1 => n5992, A2 => n5749, B1 => n5360, B2 => n2566
                           , ZN => n3217);
   U907 : OAI22_X1 port map( A1 => n5995, A2 => n5750, B1 => n5360, B2 => n2567
                           , ZN => n3218);
   U908 : OAI22_X1 port map( A1 => n5998, A2 => n5747, B1 => n5361, B2 => n2568
                           , ZN => n3219);
   U909 : OAI22_X1 port map( A1 => n6001, A2 => n5748, B1 => n5361, B2 => n2569
                           , ZN => n3220);
   U910 : OAI22_X1 port map( A1 => n6004, A2 => n5747, B1 => n5361, B2 => n2570
                           , ZN => n3221);
   U911 : OAI22_X1 port map( A1 => n6007, A2 => n5752, B1 => n5361, B2 => n2571
                           , ZN => n3222);
   U912 : OAI22_X1 port map( A1 => n6010, A2 => n5749, B1 => n5361, B2 => n2572
                           , ZN => n3223);
   U913 : OAI22_X1 port map( A1 => n6013, A2 => n5750, B1 => n5361, B2 => n2573
                           , ZN => n3224);
   U914 : OAI22_X1 port map( A1 => n6016, A2 => n5750, B1 => n5361, B2 => n2574
                           , ZN => n3225);
   U915 : OAI22_X1 port map( A1 => n6019, A2 => n5746, B1 => n5361, B2 => n2575
                           , ZN => n3226);
   U916 : OAI22_X1 port map( A1 => n6022, A2 => n5749, B1 => n5361, B2 => n2576
                           , ZN => n3227);
   U917 : OAI22_X1 port map( A1 => n6025, A2 => n5752, B1 => n5361, B2 => n2577
                           , ZN => n3228);
   U918 : OAI22_X1 port map( A1 => n6028, A2 => n5751, B1 => n5361, B2 => n2578
                           , ZN => n3229);
   U919 : OAI22_X1 port map( A1 => n6031, A2 => n5752, B1 => n5361, B2 => n2579
                           , ZN => n3230);
   U920 : OAI22_X1 port map( A1 => n5962, A2 => n5757, B1 => n5363, B2 => n2512
                           , ZN => n3239);
   U921 : OAI22_X1 port map( A1 => n5965, A2 => n5755, B1 => n5363, B2 => n2488
                           , ZN => n3240);
   U922 : OAI22_X1 port map( A1 => n5968, A2 => n5757, B1 => n5363, B2 => n2513
                           , ZN => n3241);
   U923 : OAI22_X1 port map( A1 => n5971, A2 => n5756, B1 => n5363, B2 => n2489
                           , ZN => n3242);
   U924 : OAI22_X1 port map( A1 => n5974, A2 => n5755, B1 => n5363, B2 => n2490
                           , ZN => n3243);
   U925 : OAI22_X1 port map( A1 => n5977, A2 => n5760, B1 => n5363, B2 => n2514
                           , ZN => n3244);
   U926 : OAI22_X1 port map( A1 => n5980, A2 => n5756, B1 => n5363, B2 => n2491
                           , ZN => n3245);
   U927 : OAI22_X1 port map( A1 => n5983, A2 => n5757, B1 => n5363, B2 => n2494
                           , ZN => n3246);
   U928 : OAI22_X1 port map( A1 => n5986, A2 => n5757, B1 => n5363, B2 => n2515
                           , ZN => n3247);
   U929 : OAI22_X1 port map( A1 => n5989, A2 => n5760, B1 => n5363, B2 => n2495
                           , ZN => n3248);
   U930 : OAI22_X1 port map( A1 => n5992, A2 => n5758, B1 => n5363, B2 => n2496
                           , ZN => n3249);
   U931 : OAI22_X1 port map( A1 => n5995, A2 => n5759, B1 => n5363, B2 => n2516
                           , ZN => n3250);
   U932 : OAI22_X1 port map( A1 => n5998, A2 => n5756, B1 => n5364, B2 => n2497
                           , ZN => n3251);
   U933 : OAI22_X1 port map( A1 => n6001, A2 => n5757, B1 => n5364, B2 => n2498
                           , ZN => n3252);
   U934 : OAI22_X1 port map( A1 => n6004, A2 => n5756, B1 => n5364, B2 => n2517
                           , ZN => n3253);
   U935 : OAI22_X1 port map( A1 => n6007, A2 => n5761, B1 => n5364, B2 => n2499
                           , ZN => n3254);
   U936 : OAI22_X1 port map( A1 => n6010, A2 => n5758, B1 => n5364, B2 => n2500
                           , ZN => n3255);
   U937 : OAI22_X1 port map( A1 => n6013, A2 => n5759, B1 => n5364, B2 => n2518
                           , ZN => n3256);
   U938 : OAI22_X1 port map( A1 => n6016, A2 => n5759, B1 => n5364, B2 => n2501
                           , ZN => n3257);
   U939 : OAI22_X1 port map( A1 => n6019, A2 => n5755, B1 => n5364, B2 => n2502
                           , ZN => n3258);
   U940 : OAI22_X1 port map( A1 => n6022, A2 => n5758, B1 => n5364, B2 => n2519
                           , ZN => n3259);
   U941 : OAI22_X1 port map( A1 => n6025, A2 => n5761, B1 => n5364, B2 => n2503
                           , ZN => n3260);
   U942 : OAI22_X1 port map( A1 => n6028, A2 => n5760, B1 => n5364, B2 => n2504
                           , ZN => n3261);
   U943 : OAI22_X1 port map( A1 => n6031, A2 => n5761, B1 => n5364, B2 => n2520
                           , ZN => n3262);
   U944 : OAI22_X1 port map( A1 => n5962, A2 => n5765, B1 => n5366, B2 => n2223
                           , ZN => n3271);
   U945 : OAI22_X1 port map( A1 => n5965, A2 => n5764, B1 => n5366, B2 => n2155
                           , ZN => n3272);
   U946 : OAI22_X1 port map( A1 => n5968, A2 => n5765, B1 => n5366, B2 => n2176
                           , ZN => n3273);
   U947 : OAI22_X1 port map( A1 => n5971, A2 => n5767, B1 => n5366, B2 => n2156
                           , ZN => n3274);
   U948 : OAI22_X1 port map( A1 => n5974, A2 => n5765, B1 => n5366, B2 => n2157
                           , ZN => n3275);
   U949 : OAI22_X1 port map( A1 => n5977, A2 => n5770, B1 => n5366, B2 => n2177
                           , ZN => n3276);
   U950 : OAI22_X1 port map( A1 => n5980, A2 => n5766, B1 => n5366, B2 => n2158
                           , ZN => n3277);
   U951 : OAI22_X1 port map( A1 => n5983, A2 => n5767, B1 => n5366, B2 => n2159
                           , ZN => n3278);
   U952 : OAI22_X1 port map( A1 => n5986, A2 => n5767, B1 => n5366, B2 => n2178
                           , ZN => n3279);
   U953 : OAI22_X1 port map( A1 => n5989, A2 => n5769, B1 => n5366, B2 => n2160
                           , ZN => n3280);
   U954 : OAI22_X1 port map( A1 => n5992, A2 => n5769, B1 => n5366, B2 => n2161
                           , ZN => n3281);
   U955 : OAI22_X1 port map( A1 => n5995, A2 => n5768, B1 => n5366, B2 => n2179
                           , ZN => n3282);
   U956 : OAI22_X1 port map( A1 => n5998, A2 => n5766, B1 => n5367, B2 => n2162
                           , ZN => n3283);
   U957 : OAI22_X1 port map( A1 => n6001, A2 => n5767, B1 => n5367, B2 => n2163
                           , ZN => n3284);
   U958 : OAI22_X1 port map( A1 => n6004, A2 => n5766, B1 => n5367, B2 => n2184
                           , ZN => n3285);
   U959 : OAI22_X1 port map( A1 => n6007, A2 => n5768, B1 => n5367, B2 => n2164
                           , ZN => n3286);
   U960 : OAI22_X1 port map( A1 => n6010, A2 => n5768, B1 => n5367, B2 => n2165
                           , ZN => n3287);
   U961 : OAI22_X1 port map( A1 => n6013, A2 => n5768, B1 => n5367, B2 => n2185
                           , ZN => n3288);
   U962 : OAI22_X1 port map( A1 => n6016, A2 => n5769, B1 => n5367, B2 => n2166
                           , ZN => n3289);
   U963 : OAI22_X1 port map( A1 => n6019, A2 => n5765, B1 => n5367, B2 => n2167
                           , ZN => n3290);
   U964 : OAI22_X1 port map( A1 => n6022, A2 => n5769, B1 => n5367, B2 => n2186
                           , ZN => n3291);
   U965 : OAI22_X1 port map( A1 => n6025, A2 => n5768, B1 => n5367, B2 => n2168
                           , ZN => n3292);
   U966 : OAI22_X1 port map( A1 => n6028, A2 => n5769, B1 => n5367, B2 => n2169
                           , ZN => n3293);
   U967 : OAI22_X1 port map( A1 => n6031, A2 => n5770, B1 => n5367, B2 => n2187
                           , ZN => n3294);
   U968 : OAI22_X1 port map( A1 => n5962, A2 => n5775, B1 => n5369, B2 => n5247
                           , ZN => n3303);
   U969 : OAI22_X1 port map( A1 => n5965, A2 => n5773, B1 => n5369, B2 => n5248
                           , ZN => n3304);
   U970 : OAI22_X1 port map( A1 => n5968, A2 => n5775, B1 => n5369, B2 => n5249
                           , ZN => n3305);
   U971 : OAI22_X1 port map( A1 => n5971, A2 => n5774, B1 => n5369, B2 => n5250
                           , ZN => n3306);
   U972 : OAI22_X1 port map( A1 => n5974, A2 => n5773, B1 => n5369, B2 => n5251
                           , ZN => n3307);
   U973 : OAI22_X1 port map( A1 => n5977, A2 => n5778, B1 => n5369, B2 => n5252
                           , ZN => n3308);
   U974 : OAI22_X1 port map( A1 => n5980, A2 => n5774, B1 => n5369, B2 => n5253
                           , ZN => n3309);
   U975 : OAI22_X1 port map( A1 => n5983, A2 => n5775, B1 => n5369, B2 => n5254
                           , ZN => n3310);
   U976 : OAI22_X1 port map( A1 => n5986, A2 => n5775, B1 => n5369, B2 => n5255
                           , ZN => n3311);
   U977 : OAI22_X1 port map( A1 => n5989, A2 => n5778, B1 => n5369, B2 => n5256
                           , ZN => n3312);
   U978 : OAI22_X1 port map( A1 => n5992, A2 => n5776, B1 => n5369, B2 => n5257
                           , ZN => n3313);
   U979 : OAI22_X1 port map( A1 => n5995, A2 => n5777, B1 => n5369, B2 => n5258
                           , ZN => n3314);
   U980 : OAI22_X1 port map( A1 => n5998, A2 => n5774, B1 => n5370, B2 => n5259
                           , ZN => n3315);
   U981 : OAI22_X1 port map( A1 => n6001, A2 => n5775, B1 => n5370, B2 => n5260
                           , ZN => n3316);
   U982 : OAI22_X1 port map( A1 => n6004, A2 => n5774, B1 => n5370, B2 => n5261
                           , ZN => n3317);
   U983 : OAI22_X1 port map( A1 => n6007, A2 => n5779, B1 => n5370, B2 => n5262
                           , ZN => n3318);
   U984 : OAI22_X1 port map( A1 => n6010, A2 => n5776, B1 => n5370, B2 => n5263
                           , ZN => n3319);
   U985 : OAI22_X1 port map( A1 => n6013, A2 => n5777, B1 => n5370, B2 => n5264
                           , ZN => n3320);
   U986 : OAI22_X1 port map( A1 => n6016, A2 => n5777, B1 => n5370, B2 => n5265
                           , ZN => n3321);
   U987 : OAI22_X1 port map( A1 => n6019, A2 => n5773, B1 => n5370, B2 => n5266
                           , ZN => n3322);
   U988 : OAI22_X1 port map( A1 => n6022, A2 => n5776, B1 => n5370, B2 => n5267
                           , ZN => n3323);
   U989 : OAI22_X1 port map( A1 => n6025, A2 => n5779, B1 => n5370, B2 => n5268
                           , ZN => n3324);
   U990 : OAI22_X1 port map( A1 => n6028, A2 => n5778, B1 => n5370, B2 => n5269
                           , ZN => n3325);
   U991 : OAI22_X1 port map( A1 => n6031, A2 => n5779, B1 => n5370, B2 => n5270
                           , ZN => n3326);
   U992 : OAI22_X1 port map( A1 => n5962, A2 => n5784, B1 => n5372, B2 => n2422
                           , ZN => n3335);
   U993 : OAI22_X1 port map( A1 => n5965, A2 => n5782, B1 => n5372, B2 => n5215
                           , ZN => n3336);
   U994 : OAI22_X1 port map( A1 => n5968, A2 => n5784, B1 => n5372, B2 => n5216
                           , ZN => n3337);
   U995 : OAI22_X1 port map( A1 => n5971, A2 => n5783, B1 => n5372, B2 => n5217
                           , ZN => n3338);
   U996 : OAI22_X1 port map( A1 => n5974, A2 => n5782, B1 => n5372, B2 => n5218
                           , ZN => n3339);
   U997 : OAI22_X1 port map( A1 => n5977, A2 => n5787, B1 => n5372, B2 => n5219
                           , ZN => n3340);
   U998 : OAI22_X1 port map( A1 => n5980, A2 => n5783, B1 => n5372, B2 => n5220
                           , ZN => n3341);
   U999 : OAI22_X1 port map( A1 => n5983, A2 => n5784, B1 => n5372, B2 => n5221
                           , ZN => n3342);
   U1000 : OAI22_X1 port map( A1 => n5986, A2 => n5784, B1 => n5372, B2 => 
                           n5222, ZN => n3343);
   U1001 : OAI22_X1 port map( A1 => n5989, A2 => n5787, B1 => n5372, B2 => 
                           n5223, ZN => n3344);
   U1002 : OAI22_X1 port map( A1 => n5992, A2 => n5785, B1 => n5372, B2 => 
                           n5224, ZN => n3345);
   U1003 : OAI22_X1 port map( A1 => n5995, A2 => n5786, B1 => n5372, B2 => 
                           n5225, ZN => n3346);
   U1004 : OAI22_X1 port map( A1 => n5998, A2 => n5783, B1 => n5373, B2 => 
                           n5226, ZN => n3347);
   U1005 : OAI22_X1 port map( A1 => n6001, A2 => n5784, B1 => n5373, B2 => 
                           n5227, ZN => n3348);
   U1006 : OAI22_X1 port map( A1 => n6004, A2 => n5783, B1 => n5373, B2 => 
                           n5228, ZN => n3349);
   U1007 : OAI22_X1 port map( A1 => n6007, A2 => n5788, B1 => n5373, B2 => 
                           n5229, ZN => n3350);
   U1008 : OAI22_X1 port map( A1 => n6010, A2 => n5785, B1 => n5373, B2 => 
                           n5230, ZN => n3351);
   U1009 : OAI22_X1 port map( A1 => n6013, A2 => n5786, B1 => n5373, B2 => 
                           n5231, ZN => n3352);
   U1010 : OAI22_X1 port map( A1 => n6016, A2 => n5786, B1 => n5373, B2 => 
                           n5232, ZN => n3353);
   U1011 : OAI22_X1 port map( A1 => n6019, A2 => n5782, B1 => n5373, B2 => 
                           n5233, ZN => n3354);
   U1012 : OAI22_X1 port map( A1 => n6022, A2 => n5785, B1 => n5373, B2 => 
                           n5234, ZN => n3355);
   U1013 : OAI22_X1 port map( A1 => n6025, A2 => n5788, B1 => n5373, B2 => 
                           n5235, ZN => n3356);
   U1014 : OAI22_X1 port map( A1 => n6028, A2 => n5787, B1 => n5373, B2 => 
                           n5236, ZN => n3357);
   U1015 : OAI22_X1 port map( A1 => n6031, A2 => n5788, B1 => n5373, B2 => 
                           n5237, ZN => n3358);
   U1016 : OAI22_X1 port map( A1 => n5963, A2 => n5793, B1 => n5375, B2 => 
                           n2224, ZN => n3367);
   U1017 : OAI22_X1 port map( A1 => n5966, A2 => n5791, B1 => n5375, B2 => 
                           n2930, ZN => n3368);
   U1018 : OAI22_X1 port map( A1 => n5969, A2 => n5793, B1 => n5375, B2 => 
                           n2931, ZN => n3369);
   U1019 : OAI22_X1 port map( A1 => n5972, A2 => n5792, B1 => n5375, B2 => 
                           n2932, ZN => n3370);
   U1020 : OAI22_X1 port map( A1 => n5975, A2 => n5791, B1 => n5375, B2 => 
                           n2933, ZN => n3371);
   U1021 : OAI22_X1 port map( A1 => n5978, A2 => n5796, B1 => n5375, B2 => 
                           n2934, ZN => n3372);
   U1022 : OAI22_X1 port map( A1 => n5981, A2 => n5792, B1 => n5375, B2 => 
                           n2935, ZN => n3373);
   U1023 : OAI22_X1 port map( A1 => n5984, A2 => n5793, B1 => n5375, B2 => 
                           n2936, ZN => n3374);
   U1024 : OAI22_X1 port map( A1 => n5987, A2 => n5793, B1 => n5375, B2 => 
                           n2949, ZN => n3375);
   U1025 : OAI22_X1 port map( A1 => n5990, A2 => n5796, B1 => n5375, B2 => 
                           n2937, ZN => n3376);
   U1026 : OAI22_X1 port map( A1 => n5993, A2 => n5794, B1 => n5375, B2 => 
                           n2938, ZN => n3377);
   U1027 : OAI22_X1 port map( A1 => n5996, A2 => n5795, B1 => n5375, B2 => 
                           n2939, ZN => n3378);
   U1028 : OAI22_X1 port map( A1 => n5999, A2 => n5792, B1 => n5376, B2 => 
                           n2940, ZN => n3379);
   U1029 : OAI22_X1 port map( A1 => n6002, A2 => n5793, B1 => n5376, B2 => 
                           n2941, ZN => n3380);
   U1030 : OAI22_X1 port map( A1 => n6005, A2 => n5792, B1 => n5376, B2 => 
                           n2942, ZN => n3381);
   U1031 : OAI22_X1 port map( A1 => n6008, A2 => n5797, B1 => n5376, B2 => 
                           n2943, ZN => n3382);
   U1032 : OAI22_X1 port map( A1 => n6011, A2 => n5794, B1 => n5376, B2 => 
                           n2944, ZN => n3383);
   U1033 : OAI22_X1 port map( A1 => n6014, A2 => n5795, B1 => n5376, B2 => 
                           n4166, ZN => n3384);
   U1034 : OAI22_X1 port map( A1 => n6017, A2 => n5795, B1 => n5376, B2 => 
                           n2945, ZN => n3385);
   U1035 : OAI22_X1 port map( A1 => n6020, A2 => n5791, B1 => n5376, B2 => 
                           n2946, ZN => n3386);
   U1036 : OAI22_X1 port map( A1 => n6023, A2 => n5794, B1 => n5376, B2 => 
                           n4014, ZN => n3387);
   U1037 : OAI22_X1 port map( A1 => n6026, A2 => n5797, B1 => n5376, B2 => 
                           n4033, ZN => n3388);
   U1038 : OAI22_X1 port map( A1 => n6029, A2 => n5796, B1 => n5376, B2 => 
                           n4052, ZN => n3389);
   U1039 : OAI22_X1 port map( A1 => n6032, A2 => n5797, B1 => n5376, B2 => 
                           n4071, ZN => n3390);
   U1040 : OAI22_X1 port map( A1 => n5963, A2 => n5801, B1 => n5378, B2 => 
                           n2389, ZN => n3399);
   U1041 : OAI22_X1 port map( A1 => n5966, A2 => n5800, B1 => n5378, B2 => 
                           n2391, ZN => n3400);
   U1042 : OAI22_X1 port map( A1 => n5969, A2 => n5801, B1 => n5378, B2 => 
                           n2392, ZN => n3401);
   U1043 : OAI22_X1 port map( A1 => n5972, A2 => n5803, B1 => n5378, B2 => 
                           n2393, ZN => n3402);
   U1044 : OAI22_X1 port map( A1 => n5975, A2 => n5801, B1 => n5378, B2 => 
                           n2394, ZN => n3403);
   U1045 : OAI22_X1 port map( A1 => n5978, A2 => n5806, B1 => n5378, B2 => 
                           n2395, ZN => n3404);
   U1046 : OAI22_X1 port map( A1 => n5981, A2 => n5802, B1 => n5378, B2 => 
                           n2396, ZN => n3405);
   U1047 : OAI22_X1 port map( A1 => n5984, A2 => n5803, B1 => n5378, B2 => 
                           n2397, ZN => n3406);
   U1048 : OAI22_X1 port map( A1 => n5987, A2 => n5803, B1 => n5378, B2 => 
                           n2398, ZN => n3407);
   U1049 : OAI22_X1 port map( A1 => n5990, A2 => n5805, B1 => n5378, B2 => 
                           n2399, ZN => n3408);
   U1050 : OAI22_X1 port map( A1 => n5993, A2 => n5805, B1 => n5378, B2 => 
                           n2400, ZN => n3409);
   U1051 : OAI22_X1 port map( A1 => n5996, A2 => n5804, B1 => n5378, B2 => 
                           n2401, ZN => n3410);
   U1052 : OAI22_X1 port map( A1 => n5999, A2 => n5802, B1 => n5379, B2 => 
                           n2402, ZN => n3411);
   U1053 : OAI22_X1 port map( A1 => n6002, A2 => n5803, B1 => n5379, B2 => 
                           n2403, ZN => n3412);
   U1054 : OAI22_X1 port map( A1 => n6005, A2 => n5802, B1 => n5379, B2 => 
                           n2404, ZN => n3413);
   U1055 : OAI22_X1 port map( A1 => n6008, A2 => n5804, B1 => n5379, B2 => 
                           n2405, ZN => n3414);
   U1056 : OAI22_X1 port map( A1 => n6011, A2 => n5804, B1 => n5379, B2 => 
                           n2406, ZN => n3415);
   U1057 : OAI22_X1 port map( A1 => n6014, A2 => n5804, B1 => n5379, B2 => 
                           n2407, ZN => n3416);
   U1058 : OAI22_X1 port map( A1 => n6017, A2 => n5805, B1 => n5379, B2 => 
                           n2408, ZN => n3417);
   U1059 : OAI22_X1 port map( A1 => n6020, A2 => n5801, B1 => n5379, B2 => 
                           n2409, ZN => n3418);
   U1060 : OAI22_X1 port map( A1 => n6023, A2 => n5805, B1 => n5379, B2 => 
                           n2410, ZN => n3419);
   U1061 : OAI22_X1 port map( A1 => n6026, A2 => n5804, B1 => n5379, B2 => 
                           n2411, ZN => n3420);
   U1062 : OAI22_X1 port map( A1 => n6029, A2 => n5805, B1 => n5379, B2 => 
                           n2412, ZN => n3421);
   U1063 : OAI22_X1 port map( A1 => n6032, A2 => n5806, B1 => n5379, B2 => 
                           n2413, ZN => n3422);
   U1064 : OAI22_X1 port map( A1 => n5963, A2 => n5810, B1 => n5381, B2 => 
                           n2225, ZN => n3431);
   U1065 : OAI22_X1 port map( A1 => n5966, A2 => n5809, B1 => n5381, B2 => 
                           n2190, ZN => n3432);
   U1066 : OAI22_X1 port map( A1 => n5969, A2 => n5810, B1 => n5381, B2 => 
                           n2191, ZN => n3433);
   U1067 : OAI22_X1 port map( A1 => n5972, A2 => n5812, B1 => n5381, B2 => 
                           n2192, ZN => n3434);
   U1068 : OAI22_X1 port map( A1 => n5975, A2 => n5810, B1 => n5381, B2 => 
                           n2193, ZN => n3435);
   U1069 : OAI22_X1 port map( A1 => n5978, A2 => n5815, B1 => n5381, B2 => 
                           n2194, ZN => n3436);
   U1070 : OAI22_X1 port map( A1 => n5981, A2 => n5811, B1 => n5381, B2 => 
                           n2195, ZN => n3437);
   U1071 : OAI22_X1 port map( A1 => n5984, A2 => n5812, B1 => n5381, B2 => 
                           n2196, ZN => n3438);
   U1072 : OAI22_X1 port map( A1 => n5987, A2 => n5812, B1 => n5381, B2 => 
                           n2197, ZN => n3439);
   U1073 : OAI22_X1 port map( A1 => n5990, A2 => n5814, B1 => n5381, B2 => 
                           n2198, ZN => n3440);
   U1074 : OAI22_X1 port map( A1 => n5993, A2 => n5814, B1 => n5381, B2 => 
                           n2199, ZN => n3441);
   U1075 : OAI22_X1 port map( A1 => n5996, A2 => n5813, B1 => n5381, B2 => 
                           n2200, ZN => n3442);
   U1076 : OAI22_X1 port map( A1 => n5999, A2 => n5811, B1 => n5382, B2 => 
                           n2201, ZN => n3443);
   U1077 : OAI22_X1 port map( A1 => n6002, A2 => n5812, B1 => n5382, B2 => 
                           n2202, ZN => n3444);
   U1078 : OAI22_X1 port map( A1 => n6005, A2 => n5811, B1 => n5382, B2 => 
                           n2203, ZN => n3445);
   U1079 : OAI22_X1 port map( A1 => n6008, A2 => n5813, B1 => n5382, B2 => 
                           n2204, ZN => n3446);
   U1080 : OAI22_X1 port map( A1 => n6011, A2 => n5813, B1 => n5382, B2 => 
                           n2205, ZN => n3447);
   U1081 : OAI22_X1 port map( A1 => n6014, A2 => n5813, B1 => n5382, B2 => 
                           n2206, ZN => n3448);
   U1082 : OAI22_X1 port map( A1 => n6017, A2 => n5814, B1 => n5382, B2 => 
                           n2207, ZN => n3449);
   U1083 : OAI22_X1 port map( A1 => n6020, A2 => n5810, B1 => n5382, B2 => 
                           n2208, ZN => n3450);
   U1084 : OAI22_X1 port map( A1 => n6023, A2 => n5814, B1 => n5382, B2 => 
                           n2209, ZN => n3451);
   U1085 : OAI22_X1 port map( A1 => n6026, A2 => n5813, B1 => n5382, B2 => 
                           n2210, ZN => n3452);
   U1086 : OAI22_X1 port map( A1 => n6029, A2 => n5814, B1 => n5382, B2 => 
                           n2211, ZN => n3453);
   U1087 : OAI22_X1 port map( A1 => n6032, A2 => n5815, B1 => n5382, B2 => 
                           n2212, ZN => n3454);
   U1088 : OAI22_X1 port map( A1 => n5963, A2 => n5819, B1 => n5384, B2 => 
                           n5238, ZN => n3463);
   U1089 : OAI22_X1 port map( A1 => n5966, A2 => n5818, B1 => n5384, B2 => 
                           n2423, ZN => n3464);
   U1090 : OAI22_X1 port map( A1 => n5969, A2 => n5819, B1 => n5384, B2 => 
                           n2445, ZN => n3465);
   U1091 : OAI22_X1 port map( A1 => n5972, A2 => n5821, B1 => n5384, B2 => 
                           n2425, ZN => n3466);
   U1092 : OAI22_X1 port map( A1 => n5975, A2 => n5819, B1 => n5384, B2 => 
                           n2426, ZN => n3467);
   U1093 : OAI22_X1 port map( A1 => n5978, A2 => n5824, B1 => n5384, B2 => 
                           n2446, ZN => n3468);
   U1094 : OAI22_X1 port map( A1 => n5981, A2 => n5820, B1 => n5384, B2 => 
                           n2427, ZN => n3469);
   U1095 : OAI22_X1 port map( A1 => n5984, A2 => n5821, B1 => n5384, B2 => 
                           n2428, ZN => n3470);
   U1096 : OAI22_X1 port map( A1 => n5987, A2 => n5821, B1 => n5384, B2 => 
                           n2447, ZN => n3471);
   U1097 : OAI22_X1 port map( A1 => n5990, A2 => n5823, B1 => n5384, B2 => 
                           n2429, ZN => n3472);
   U1098 : OAI22_X1 port map( A1 => n5993, A2 => n5823, B1 => n5384, B2 => 
                           n2430, ZN => n3473);
   U1099 : OAI22_X1 port map( A1 => n5996, A2 => n5822, B1 => n5384, B2 => 
                           n2448, ZN => n3474);
   U1100 : OAI22_X1 port map( A1 => n5999, A2 => n5820, B1 => n5385, B2 => 
                           n2431, ZN => n3475);
   U1101 : OAI22_X1 port map( A1 => n6002, A2 => n5821, B1 => n5385, B2 => 
                           n2432, ZN => n3476);
   U1102 : OAI22_X1 port map( A1 => n6005, A2 => n5820, B1 => n5385, B2 => 
                           n2449, ZN => n3477);
   U1103 : OAI22_X1 port map( A1 => n6008, A2 => n5822, B1 => n5385, B2 => 
                           n2433, ZN => n3478);
   U1104 : OAI22_X1 port map( A1 => n6011, A2 => n5822, B1 => n5385, B2 => 
                           n2434, ZN => n3479);
   U1105 : OAI22_X1 port map( A1 => n6014, A2 => n5822, B1 => n5385, B2 => 
                           n2450, ZN => n3480);
   U1106 : OAI22_X1 port map( A1 => n6017, A2 => n5823, B1 => n5385, B2 => 
                           n2435, ZN => n3481);
   U1107 : OAI22_X1 port map( A1 => n6020, A2 => n5819, B1 => n5385, B2 => 
                           n2436, ZN => n3482);
   U1108 : OAI22_X1 port map( A1 => n6023, A2 => n5823, B1 => n5385, B2 => 
                           n2451, ZN => n3483);
   U1109 : OAI22_X1 port map( A1 => n6026, A2 => n5822, B1 => n5385, B2 => 
                           n2437, ZN => n3484);
   U1110 : OAI22_X1 port map( A1 => n6029, A2 => n5823, B1 => n5385, B2 => 
                           n2438, ZN => n3485);
   U1111 : OAI22_X1 port map( A1 => n6032, A2 => n5824, B1 => n5385, B2 => 
                           n2452, ZN => n3486);
   U1112 : OAI22_X1 port map( A1 => n5963, A2 => n5829, B1 => n5387, B2 => 
                           n2154, ZN => n3495);
   U1113 : OAI22_X1 port map( A1 => n5966, A2 => n5827, B1 => n5387, B2 => 
                           n5184, ZN => n3496);
   U1114 : OAI22_X1 port map( A1 => n5969, A2 => n5829, B1 => n5387, B2 => 
                           n5205, ZN => n3497);
   U1115 : OAI22_X1 port map( A1 => n5972, A2 => n5828, B1 => n5387, B2 => 
                           n5185, ZN => n3498);
   U1116 : OAI22_X1 port map( A1 => n5975, A2 => n5827, B1 => n5387, B2 => 
                           n5186, ZN => n3499);
   U1117 : OAI22_X1 port map( A1 => n5978, A2 => n5832, B1 => n5387, B2 => 
                           n5206, ZN => n3500);
   U1118 : OAI22_X1 port map( A1 => n5981, A2 => n5828, B1 => n5387, B2 => 
                           n5187, ZN => n3501);
   U1119 : OAI22_X1 port map( A1 => n5984, A2 => n5829, B1 => n5387, B2 => 
                           n5188, ZN => n3502);
   U1120 : OAI22_X1 port map( A1 => n5987, A2 => n5829, B1 => n5387, B2 => 
                           n5207, ZN => n3503);
   U1121 : OAI22_X1 port map( A1 => n5990, A2 => n5832, B1 => n5387, B2 => 
                           n5189, ZN => n3504);
   U1122 : OAI22_X1 port map( A1 => n5993, A2 => n5830, B1 => n5387, B2 => 
                           n5190, ZN => n3505);
   U1123 : OAI22_X1 port map( A1 => n5996, A2 => n5831, B1 => n5387, B2 => 
                           n5208, ZN => n3506);
   U1124 : OAI22_X1 port map( A1 => n5999, A2 => n5828, B1 => n5388, B2 => 
                           n5191, ZN => n3507);
   U1125 : OAI22_X1 port map( A1 => n6002, A2 => n5829, B1 => n5388, B2 => 
                           n5192, ZN => n3508);
   U1126 : OAI22_X1 port map( A1 => n6005, A2 => n5828, B1 => n5388, B2 => 
                           n5209, ZN => n3509);
   U1127 : OAI22_X1 port map( A1 => n6008, A2 => n5833, B1 => n5388, B2 => 
                           n5193, ZN => n3510);
   U1128 : OAI22_X1 port map( A1 => n6011, A2 => n5830, B1 => n5388, B2 => 
                           n5194, ZN => n3511);
   U1129 : OAI22_X1 port map( A1 => n6014, A2 => n5831, B1 => n5388, B2 => 
                           n5210, ZN => n3512);
   U1130 : OAI22_X1 port map( A1 => n6017, A2 => n5831, B1 => n5388, B2 => 
                           n5195, ZN => n3513);
   U1131 : OAI22_X1 port map( A1 => n6020, A2 => n5827, B1 => n5388, B2 => 
                           n5196, ZN => n3514);
   U1132 : OAI22_X1 port map( A1 => n6023, A2 => n5830, B1 => n5388, B2 => 
                           n5211, ZN => n3515);
   U1133 : OAI22_X1 port map( A1 => n6026, A2 => n5833, B1 => n5388, B2 => 
                           n5197, ZN => n3516);
   U1134 : OAI22_X1 port map( A1 => n6029, A2 => n5832, B1 => n5388, B2 => 
                           n5198, ZN => n3517);
   U1135 : OAI22_X1 port map( A1 => n6032, A2 => n5833, B1 => n5388, B2 => 
                           n5212, ZN => n3518);
   U1136 : OAI22_X1 port map( A1 => n5963, A2 => n5846, B1 => n5393, B2 => 
                           n2319, ZN => n3559);
   U1137 : OAI22_X1 port map( A1 => n5966, A2 => n5845, B1 => n5393, B2 => 
                           n2322, ZN => n3560);
   U1138 : OAI22_X1 port map( A1 => n5969, A2 => n5846, B1 => n5393, B2 => 
                           n2323, ZN => n3561);
   U1139 : OAI22_X1 port map( A1 => n5972, A2 => n5848, B1 => n5393, B2 => 
                           n2324, ZN => n3562);
   U1140 : OAI22_X1 port map( A1 => n5975, A2 => n5846, B1 => n5393, B2 => 
                           n2325, ZN => n3563);
   U1141 : OAI22_X1 port map( A1 => n5978, A2 => n5851, B1 => n5393, B2 => 
                           n2326, ZN => n3564);
   U1142 : OAI22_X1 port map( A1 => n5981, A2 => n5847, B1 => n5393, B2 => 
                           n2327, ZN => n3565);
   U1143 : OAI22_X1 port map( A1 => n5984, A2 => n5848, B1 => n5393, B2 => 
                           n2328, ZN => n3566);
   U1144 : OAI22_X1 port map( A1 => n5987, A2 => n5848, B1 => n5393, B2 => 
                           n2329, ZN => n3567);
   U1145 : OAI22_X1 port map( A1 => n5990, A2 => n5850, B1 => n5393, B2 => 
                           n2330, ZN => n3568);
   U1146 : OAI22_X1 port map( A1 => n5993, A2 => n5850, B1 => n5393, B2 => 
                           n2331, ZN => n3569);
   U1147 : OAI22_X1 port map( A1 => n5996, A2 => n5849, B1 => n5393, B2 => 
                           n2332, ZN => n3570);
   U1148 : OAI22_X1 port map( A1 => n5999, A2 => n5847, B1 => n5394, B2 => 
                           n2333, ZN => n3571);
   U1149 : OAI22_X1 port map( A1 => n6002, A2 => n5848, B1 => n5394, B2 => 
                           n2334, ZN => n3572);
   U1150 : OAI22_X1 port map( A1 => n6005, A2 => n5847, B1 => n5394, B2 => 
                           n2335, ZN => n3573);
   U1151 : OAI22_X1 port map( A1 => n6008, A2 => n5849, B1 => n5394, B2 => 
                           n2336, ZN => n3574);
   U1152 : OAI22_X1 port map( A1 => n6011, A2 => n5849, B1 => n5394, B2 => 
                           n2337, ZN => n3575);
   U1153 : OAI22_X1 port map( A1 => n6014, A2 => n5849, B1 => n5394, B2 => 
                           n2338, ZN => n3576);
   U1154 : OAI22_X1 port map( A1 => n6017, A2 => n5850, B1 => n5394, B2 => 
                           n2339, ZN => n3577);
   U1155 : OAI22_X1 port map( A1 => n6020, A2 => n5846, B1 => n5394, B2 => 
                           n2340, ZN => n3578);
   U1156 : OAI22_X1 port map( A1 => n6023, A2 => n5850, B1 => n5394, B2 => 
                           n2341, ZN => n3579);
   U1157 : OAI22_X1 port map( A1 => n6026, A2 => n5849, B1 => n5394, B2 => 
                           n2342, ZN => n3580);
   U1158 : OAI22_X1 port map( A1 => n6029, A2 => n5850, B1 => n5394, B2 => 
                           n2343, ZN => n3581);
   U1159 : OAI22_X1 port map( A1 => n6032, A2 => n5851, B1 => n5394, B2 => 
                           n2344, ZN => n3582);
   U1160 : OAI22_X1 port map( A1 => n5963, A2 => n5864, B1 => n5399, B2 => 
                           n5311, ZN => n3623);
   U1161 : OAI22_X1 port map( A1 => n5966, A2 => n5863, B1 => n5399, B2 => 
                           n2288, ZN => n3624);
   U1162 : OAI22_X1 port map( A1 => n5969, A2 => n5864, B1 => n5399, B2 => 
                           n2289, ZN => n3625);
   U1163 : OAI22_X1 port map( A1 => n5972, A2 => n5866, B1 => n5399, B2 => 
                           n2290, ZN => n3626);
   U1164 : OAI22_X1 port map( A1 => n5975, A2 => n5864, B1 => n5399, B2 => 
                           n2291, ZN => n3627);
   U1165 : OAI22_X1 port map( A1 => n5978, A2 => n5869, B1 => n5399, B2 => 
                           n2292, ZN => n3628);
   U1166 : OAI22_X1 port map( A1 => n5981, A2 => n5865, B1 => n5399, B2 => 
                           n2293, ZN => n3629);
   U1167 : OAI22_X1 port map( A1 => n5984, A2 => n5866, B1 => n5399, B2 => 
                           n2294, ZN => n3630);
   U1168 : OAI22_X1 port map( A1 => n5987, A2 => n5866, B1 => n5399, B2 => 
                           n2295, ZN => n3631);
   U1169 : OAI22_X1 port map( A1 => n5990, A2 => n5868, B1 => n5399, B2 => 
                           n2296, ZN => n3632);
   U1170 : OAI22_X1 port map( A1 => n5993, A2 => n5868, B1 => n5399, B2 => 
                           n2297, ZN => n3633);
   U1171 : OAI22_X1 port map( A1 => n5996, A2 => n5867, B1 => n5399, B2 => 
                           n2298, ZN => n3634);
   U1172 : OAI22_X1 port map( A1 => n5999, A2 => n5865, B1 => n5400, B2 => 
                           n2299, ZN => n3635);
   U1173 : OAI22_X1 port map( A1 => n6002, A2 => n5866, B1 => n5400, B2 => 
                           n2300, ZN => n3636);
   U1174 : OAI22_X1 port map( A1 => n6005, A2 => n5865, B1 => n5400, B2 => 
                           n2301, ZN => n3637);
   U1175 : OAI22_X1 port map( A1 => n6008, A2 => n5867, B1 => n5400, B2 => 
                           n2302, ZN => n3638);
   U1176 : OAI22_X1 port map( A1 => n6011, A2 => n5867, B1 => n5400, B2 => 
                           n2303, ZN => n3639);
   U1177 : OAI22_X1 port map( A1 => n6014, A2 => n5867, B1 => n5400, B2 => 
                           n2304, ZN => n3640);
   U1178 : OAI22_X1 port map( A1 => n6017, A2 => n5868, B1 => n5400, B2 => 
                           n2305, ZN => n3641);
   U1179 : OAI22_X1 port map( A1 => n6020, A2 => n5864, B1 => n5400, B2 => 
                           n2306, ZN => n3642);
   U1180 : OAI22_X1 port map( A1 => n6023, A2 => n5868, B1 => n5400, B2 => 
                           n2307, ZN => n3643);
   U1181 : OAI22_X1 port map( A1 => n6026, A2 => n5867, B1 => n5400, B2 => 
                           n2308, ZN => n3644);
   U1182 : OAI22_X1 port map( A1 => n6029, A2 => n5868, B1 => n5400, B2 => 
                           n2309, ZN => n3645);
   U1183 : OAI22_X1 port map( A1 => n6032, A2 => n5869, B1 => n5400, B2 => 
                           n2310, ZN => n3646);
   U1184 : OAI22_X1 port map( A1 => n5963, A2 => n5872, B1 => n5402, B2 => 
                           n2680, ZN => n3655);
   U1185 : OAI22_X1 port map( A1 => n5966, A2 => n5872, B1 => n5402, B2 => 
                           n2681, ZN => n3656);
   U1186 : OAI22_X1 port map( A1 => n5969, A2 => n5874, B1 => n5402, B2 => 
                           n2682, ZN => n3657);
   U1187 : OAI22_X1 port map( A1 => n5972, A2 => n5873, B1 => n5402, B2 => 
                           n2683, ZN => n3658);
   U1188 : OAI22_X1 port map( A1 => n5975, A2 => n5872, B1 => n5402, B2 => 
                           n2684, ZN => n3659);
   U1189 : OAI22_X1 port map( A1 => n5978, A2 => n5877, B1 => n5402, B2 => 
                           n2685, ZN => n3660);
   U1190 : OAI22_X1 port map( A1 => n5981, A2 => n5873, B1 => n5402, B2 => 
                           n2686, ZN => n3661);
   U1191 : OAI22_X1 port map( A1 => n5984, A2 => n5874, B1 => n5402, B2 => 
                           n2687, ZN => n3662);
   U1192 : OAI22_X1 port map( A1 => n5987, A2 => n5874, B1 => n5402, B2 => 
                           n2688, ZN => n3663);
   U1193 : OAI22_X1 port map( A1 => n5990, A2 => n5877, B1 => n5402, B2 => 
                           n2689, ZN => n3664);
   U1194 : OAI22_X1 port map( A1 => n5993, A2 => n5875, B1 => n5402, B2 => 
                           n2690, ZN => n3665);
   U1195 : OAI22_X1 port map( A1 => n5996, A2 => n5876, B1 => n5402, B2 => 
                           n2691, ZN => n3666);
   U1196 : OAI22_X1 port map( A1 => n5999, A2 => n5873, B1 => n5403, B2 => 
                           n2692, ZN => n3667);
   U1197 : OAI22_X1 port map( A1 => n6002, A2 => n5874, B1 => n5403, B2 => 
                           n2693, ZN => n3668);
   U1198 : OAI22_X1 port map( A1 => n6005, A2 => n5873, B1 => n5403, B2 => 
                           n2694, ZN => n3669);
   U1199 : OAI22_X1 port map( A1 => n6008, A2 => n5878, B1 => n5403, B2 => 
                           n2695, ZN => n3670);
   U1200 : OAI22_X1 port map( A1 => n6011, A2 => n5875, B1 => n5403, B2 => 
                           n2696, ZN => n3671);
   U1201 : OAI22_X1 port map( A1 => n6014, A2 => n5876, B1 => n5403, B2 => 
                           n2697, ZN => n3672);
   U1202 : OAI22_X1 port map( A1 => n6017, A2 => n5876, B1 => n5403, B2 => 
                           n2698, ZN => n3673);
   U1203 : OAI22_X1 port map( A1 => n6020, A2 => n5872, B1 => n5403, B2 => 
                           n2701, ZN => n3674);
   U1204 : OAI22_X1 port map( A1 => n6023, A2 => n5875, B1 => n5403, B2 => 
                           n2756, ZN => n3675);
   U1205 : OAI22_X1 port map( A1 => n6026, A2 => n5878, B1 => n5403, B2 => 
                           n2775, ZN => n3676);
   U1206 : OAI22_X1 port map( A1 => n6029, A2 => n5877, B1 => n5403, B2 => 
                           n2794, ZN => n3677);
   U1207 : OAI22_X1 port map( A1 => n6032, A2 => n5878, B1 => n5403, B2 => 
                           n2813, ZN => n3678);
   U1208 : OAI22_X1 port map( A1 => n5963, A2 => n5881, B1 => n5405, B2 => 
                           n2226, ZN => n3687);
   U1209 : OAI22_X1 port map( A1 => n5966, A2 => n5882, B1 => n5405, B2 => 
                           n2228, ZN => n3688);
   U1210 : OAI22_X1 port map( A1 => n5969, A2 => n5886, B1 => n5405, B2 => 
                           n2248, ZN => n3689);
   U1211 : OAI22_X1 port map( A1 => n5972, A2 => n5885, B1 => n5405, B2 => 
                           n2229, ZN => n3690);
   U1212 : OAI22_X1 port map( A1 => n5975, A2 => n5882, B1 => n5405, B2 => 
                           n2230, ZN => n3691);
   U1213 : OAI22_X1 port map( A1 => n5978, A2 => n5883, B1 => n5405, B2 => 
                           n2249, ZN => n3692);
   U1214 : OAI22_X1 port map( A1 => n5981, A2 => n5883, B1 => n5405, B2 => 
                           n2231, ZN => n3693);
   U1215 : OAI22_X1 port map( A1 => n5984, A2 => n5883, B1 => n5405, B2 => 
                           n2232, ZN => n3694);
   U1216 : OAI22_X1 port map( A1 => n5987, A2 => n5882, B1 => n5405, B2 => 
                           n2250, ZN => n3695);
   U1217 : OAI22_X1 port map( A1 => n5990, A2 => n5882, B1 => n5405, B2 => 
                           n2233, ZN => n3696);
   U1218 : OAI22_X1 port map( A1 => n5993, A2 => n5884, B1 => n5405, B2 => 
                           n2234, ZN => n3697);
   U1219 : OAI22_X1 port map( A1 => n5996, A2 => n5885, B1 => n5405, B2 => 
                           n2251, ZN => n3698);
   U1220 : OAI22_X1 port map( A1 => n5999, A2 => n5883, B1 => n5406, B2 => 
                           n2235, ZN => n3699);
   U1221 : OAI22_X1 port map( A1 => n6002, A2 => n5883, B1 => n5406, B2 => 
                           n2236, ZN => n3700);
   U1222 : OAI22_X1 port map( A1 => n6005, A2 => n5884, B1 => n5406, B2 => 
                           n2253, ZN => n3701);
   U1223 : OAI22_X1 port map( A1 => n6008, A2 => n5881, B1 => n5406, B2 => 
                           n2237, ZN => n3702);
   U1224 : OAI22_X1 port map( A1 => n6011, A2 => n5884, B1 => n5406, B2 => 
                           n2238, ZN => n3703);
   U1225 : OAI22_X1 port map( A1 => n6014, A2 => n5885, B1 => n5406, B2 => 
                           n2254, ZN => n3704);
   U1226 : OAI22_X1 port map( A1 => n6017, A2 => n5885, B1 => n5406, B2 => 
                           n2239, ZN => n3705);
   U1227 : OAI22_X1 port map( A1 => n6020, A2 => n5882, B1 => n5406, B2 => 
                           n2240, ZN => n3706);
   U1228 : OAI22_X1 port map( A1 => n6023, A2 => n5884, B1 => n5406, B2 => 
                           n2255, ZN => n3707);
   U1229 : OAI22_X1 port map( A1 => n6026, A2 => n5887, B1 => n5406, B2 => 
                           n2241, ZN => n3708);
   U1230 : OAI22_X1 port map( A1 => n6029, A2 => n5886, B1 => n5406, B2 => 
                           n2242, ZN => n3709);
   U1231 : OAI22_X1 port map( A1 => n6032, A2 => n5887, B1 => n5406, B2 => 
                           n2256, ZN => n3710);
   U1232 : OAI22_X1 port map( A1 => n5963, A2 => n5892, B1 => n5408, B2 => 
                           n2387, ZN => n3719);
   U1233 : OAI22_X1 port map( A1 => n5966, A2 => n5890, B1 => n5408, B2 => 
                           n4223, ZN => n3720);
   U1234 : OAI22_X1 port map( A1 => n5969, A2 => n5892, B1 => n5408, B2 => 
                           n4242, ZN => n3721);
   U1235 : OAI22_X1 port map( A1 => n5972, A2 => n5891, B1 => n5408, B2 => 
                           n4261, ZN => n3722);
   U1236 : OAI22_X1 port map( A1 => n5975, A2 => n5890, B1 => n5408, B2 => 
                           n4280, ZN => n3723);
   U1237 : OAI22_X1 port map( A1 => n5978, A2 => n5895, B1 => n5408, B2 => 
                           n4299, ZN => n3724);
   U1238 : OAI22_X1 port map( A1 => n5981, A2 => n5891, B1 => n5408, B2 => 
                           n4318, ZN => n3725);
   U1239 : OAI22_X1 port map( A1 => n5984, A2 => n5892, B1 => n5408, B2 => 
                           n4337, ZN => n3726);
   U1240 : OAI22_X1 port map( A1 => n5987, A2 => n5892, B1 => n5408, B2 => 
                           n4356, ZN => n3727);
   U1241 : OAI22_X1 port map( A1 => n5990, A2 => n5895, B1 => n5408, B2 => 
                           n4375, ZN => n3728);
   U1242 : OAI22_X1 port map( A1 => n5993, A2 => n5893, B1 => n5408, B2 => 
                           n4394, ZN => n3729);
   U1243 : OAI22_X1 port map( A1 => n5996, A2 => n5894, B1 => n5408, B2 => 
                           n4416, ZN => n3730);
   U1244 : OAI22_X1 port map( A1 => n5999, A2 => n5891, B1 => n5409, B2 => 
                           n4431, ZN => n3731);
   U1245 : OAI22_X1 port map( A1 => n6002, A2 => n5892, B1 => n5409, B2 => 
                           n5103, ZN => n3732);
   U1246 : OAI22_X1 port map( A1 => n6005, A2 => n5891, B1 => n5409, B2 => 
                           n5104, ZN => n3733);
   U1247 : OAI22_X1 port map( A1 => n6008, A2 => n5896, B1 => n5409, B2 => 
                           n5105, ZN => n3734);
   U1248 : OAI22_X1 port map( A1 => n6011, A2 => n5893, B1 => n5409, B2 => 
                           n5106, ZN => n3735);
   U1249 : OAI22_X1 port map( A1 => n6014, A2 => n5894, B1 => n5409, B2 => 
                           n5107, ZN => n3736);
   U1250 : OAI22_X1 port map( A1 => n6017, A2 => n5894, B1 => n5409, B2 => 
                           n5108, ZN => n3737);
   U1251 : OAI22_X1 port map( A1 => n6020, A2 => n5890, B1 => n5409, B2 => 
                           n5109, ZN => n3738);
   U1252 : OAI22_X1 port map( A1 => n6023, A2 => n5893, B1 => n5409, B2 => 
                           n5110, ZN => n3739);
   U1253 : OAI22_X1 port map( A1 => n6026, A2 => n5896, B1 => n5409, B2 => 
                           n5111, ZN => n3740);
   U1254 : OAI22_X1 port map( A1 => n6029, A2 => n5895, B1 => n5409, B2 => 
                           n5112, ZN => n3741);
   U1255 : OAI22_X1 port map( A1 => n6032, A2 => n5896, B1 => n5409, B2 => 
                           n5113, ZN => n3742);
   U1256 : OAI22_X1 port map( A1 => n5963, A2 => n5908, B1 => n5414, B2 => 
                           n5122, ZN => n3783);
   U1257 : OAI22_X1 port map( A1 => n5966, A2 => n5909, B1 => n5414, B2 => 
                           n5124, ZN => n3784);
   U1258 : OAI22_X1 port map( A1 => n5969, A2 => n5913, B1 => n5414, B2 => 
                           n5145, ZN => n3785);
   U1259 : OAI22_X1 port map( A1 => n5972, A2 => n5912, B1 => n5414, B2 => 
                           n5125, ZN => n3786);
   U1260 : OAI22_X1 port map( A1 => n5975, A2 => n5909, B1 => n5414, B2 => 
                           n5126, ZN => n3787);
   U1261 : OAI22_X1 port map( A1 => n5978, A2 => n5910, B1 => n5414, B2 => 
                           n5146, ZN => n3788);
   U1262 : OAI22_X1 port map( A1 => n5981, A2 => n5910, B1 => n5414, B2 => 
                           n5127, ZN => n3789);
   U1263 : OAI22_X1 port map( A1 => n5984, A2 => n5910, B1 => n5414, B2 => 
                           n5128, ZN => n3790);
   U1264 : OAI22_X1 port map( A1 => n5987, A2 => n5909, B1 => n5414, B2 => 
                           n5147, ZN => n3791);
   U1265 : OAI22_X1 port map( A1 => n5990, A2 => n5909, B1 => n5414, B2 => 
                           n5129, ZN => n3792);
   U1266 : OAI22_X1 port map( A1 => n5993, A2 => n5911, B1 => n5414, B2 => 
                           n5130, ZN => n3793);
   U1267 : OAI22_X1 port map( A1 => n5996, A2 => n5912, B1 => n5414, B2 => 
                           n5148, ZN => n3794);
   U1268 : OAI22_X1 port map( A1 => n5999, A2 => n5910, B1 => n5415, B2 => 
                           n5131, ZN => n3795);
   U1269 : OAI22_X1 port map( A1 => n6002, A2 => n5910, B1 => n5415, B2 => 
                           n5132, ZN => n3796);
   U1270 : OAI22_X1 port map( A1 => n6005, A2 => n5911, B1 => n5415, B2 => 
                           n5149, ZN => n3797);
   U1271 : OAI22_X1 port map( A1 => n6008, A2 => n5908, B1 => n5415, B2 => 
                           n5133, ZN => n3798);
   U1272 : OAI22_X1 port map( A1 => n6011, A2 => n5911, B1 => n5415, B2 => 
                           n5134, ZN => n3799);
   U1273 : OAI22_X1 port map( A1 => n6014, A2 => n5912, B1 => n5415, B2 => 
                           n5150, ZN => n3800);
   U1274 : OAI22_X1 port map( A1 => n6017, A2 => n5912, B1 => n5415, B2 => 
                           n5135, ZN => n3801);
   U1275 : OAI22_X1 port map( A1 => n6020, A2 => n5909, B1 => n5415, B2 => 
                           n5136, ZN => n3802);
   U1276 : OAI22_X1 port map( A1 => n6023, A2 => n5911, B1 => n5415, B2 => 
                           n5151, ZN => n3803);
   U1277 : OAI22_X1 port map( A1 => n6026, A2 => n5914, B1 => n5415, B2 => 
                           n5137, ZN => n3804);
   U1278 : OAI22_X1 port map( A1 => n6029, A2 => n5913, B1 => n5415, B2 => 
                           n5138, ZN => n3805);
   U1279 : OAI22_X1 port map( A1 => n6032, A2 => n5914, B1 => n5415, B2 => 
                           n5152, ZN => n3806);
   U1280 : OAI22_X1 port map( A1 => n5964, A2 => n5917, B1 => n5417, B2 => 
                           n2227, ZN => n3815);
   U1281 : OAI22_X1 port map( A1 => n5967, A2 => n5918, B1 => n5417, B2 => 
                           n2258, ZN => n3816);
   U1282 : OAI22_X1 port map( A1 => n5970, A2 => n5922, B1 => n5417, B2 => 
                           n2259, ZN => n3817);
   U1283 : OAI22_X1 port map( A1 => n5973, A2 => n5921, B1 => n5417, B2 => 
                           n2260, ZN => n3818);
   U1284 : OAI22_X1 port map( A1 => n5976, A2 => n5918, B1 => n5417, B2 => 
                           n2261, ZN => n3819);
   U1285 : OAI22_X1 port map( A1 => n5979, A2 => n5919, B1 => n5417, B2 => 
                           n2262, ZN => n3820);
   U1286 : OAI22_X1 port map( A1 => n5982, A2 => n5919, B1 => n5417, B2 => 
                           n2263, ZN => n3821);
   U1287 : OAI22_X1 port map( A1 => n5985, A2 => n5919, B1 => n5417, B2 => 
                           n2264, ZN => n3822);
   U1288 : OAI22_X1 port map( A1 => n5988, A2 => n5918, B1 => n5417, B2 => 
                           n2265, ZN => n3823);
   U1289 : OAI22_X1 port map( A1 => n5991, A2 => n5918, B1 => n5417, B2 => 
                           n2266, ZN => n3824);
   U1290 : OAI22_X1 port map( A1 => n5994, A2 => n5920, B1 => n5417, B2 => 
                           n2267, ZN => n3825);
   U1291 : OAI22_X1 port map( A1 => n5997, A2 => n5921, B1 => n5417, B2 => 
                           n2268, ZN => n3826);
   U1292 : OAI22_X1 port map( A1 => n6000, A2 => n5919, B1 => n5418, B2 => 
                           n2269, ZN => n3827);
   U1293 : OAI22_X1 port map( A1 => n6003, A2 => n5919, B1 => n5418, B2 => 
                           n2270, ZN => n3828);
   U1294 : OAI22_X1 port map( A1 => n6006, A2 => n5920, B1 => n5418, B2 => 
                           n2271, ZN => n3829);
   U1295 : OAI22_X1 port map( A1 => n6009, A2 => n5917, B1 => n5418, B2 => 
                           n2272, ZN => n3830);
   U1296 : OAI22_X1 port map( A1 => n6012, A2 => n5920, B1 => n5418, B2 => 
                           n2273, ZN => n3831);
   U1297 : OAI22_X1 port map( A1 => n6015, A2 => n5921, B1 => n5418, B2 => 
                           n2274, ZN => n3832);
   U1298 : OAI22_X1 port map( A1 => n6018, A2 => n5921, B1 => n5418, B2 => 
                           n2275, ZN => n3833);
   U1299 : OAI22_X1 port map( A1 => n6021, A2 => n5918, B1 => n5418, B2 => 
                           n2276, ZN => n3834);
   U1300 : OAI22_X1 port map( A1 => n6024, A2 => n5920, B1 => n5418, B2 => 
                           n2277, ZN => n3835);
   U1301 : OAI22_X1 port map( A1 => n6027, A2 => n5923, B1 => n5418, B2 => 
                           n2278, ZN => n3836);
   U1302 : OAI22_X1 port map( A1 => n6030, A2 => n5922, B1 => n5418, B2 => 
                           n2279, ZN => n3837);
   U1303 : OAI22_X1 port map( A1 => n6033, A2 => n5922, B1 => n5418, B2 => 
                           n2280, ZN => n3838);
   U1304 : OAI22_X1 port map( A1 => n5964, A2 => n5936, B1 => n5423, B2 => 
                           n2511, ZN => n3879);
   U1305 : OAI22_X1 port map( A1 => n5967, A2 => n5935, B1 => n5423, B2 => 
                           n2121, ZN => n3880);
   U1306 : OAI22_X1 port map( A1 => n5970, A2 => n5936, B1 => n5423, B2 => 
                           n2122, ZN => n3881);
   U1307 : OAI22_X1 port map( A1 => n5973, A2 => n5938, B1 => n5423, B2 => 
                           n2123, ZN => n3882);
   U1308 : OAI22_X1 port map( A1 => n5976, A2 => n5936, B1 => n5423, B2 => 
                           n2124, ZN => n3883);
   U1309 : OAI22_X1 port map( A1 => n5979, A2 => n5941, B1 => n5423, B2 => 
                           n2125, ZN => n3884);
   U1310 : OAI22_X1 port map( A1 => n5982, A2 => n5937, B1 => n5423, B2 => 
                           n2126, ZN => n3885);
   U1311 : OAI22_X1 port map( A1 => n5985, A2 => n5938, B1 => n5423, B2 => 
                           n2127, ZN => n3886);
   U1312 : OAI22_X1 port map( A1 => n5988, A2 => n5938, B1 => n5423, B2 => 
                           n2140, ZN => n3887);
   U1313 : OAI22_X1 port map( A1 => n5991, A2 => n5940, B1 => n5423, B2 => 
                           n2128, ZN => n3888);
   U1314 : OAI22_X1 port map( A1 => n5994, A2 => n5940, B1 => n5423, B2 => 
                           n2129, ZN => n3889);
   U1315 : OAI22_X1 port map( A1 => n5997, A2 => n5939, B1 => n5423, B2 => 
                           n2130, ZN => n3890);
   U1316 : OAI22_X1 port map( A1 => n6000, A2 => n5937, B1 => n5424, B2 => 
                           n2131, ZN => n3891);
   U1317 : OAI22_X1 port map( A1 => n6003, A2 => n5938, B1 => n5424, B2 => 
                           n2132, ZN => n3892);
   U1318 : OAI22_X1 port map( A1 => n6006, A2 => n5937, B1 => n5424, B2 => 
                           n2133, ZN => n3893);
   U1319 : OAI22_X1 port map( A1 => n6009, A2 => n5939, B1 => n5424, B2 => 
                           n2134, ZN => n3894);
   U1320 : OAI22_X1 port map( A1 => n6012, A2 => n5939, B1 => n5424, B2 => 
                           n2135, ZN => n3895);
   U1321 : OAI22_X1 port map( A1 => n6015, A2 => n5939, B1 => n5424, B2 => 
                           n2150, ZN => n3896);
   U1322 : OAI22_X1 port map( A1 => n6018, A2 => n5940, B1 => n5424, B2 => 
                           n2136, ZN => n3897);
   U1323 : OAI22_X1 port map( A1 => n6021, A2 => n5936, B1 => n5424, B2 => 
                           n2137, ZN => n3898);
   U1324 : OAI22_X1 port map( A1 => n6024, A2 => n5940, B1 => n5424, B2 => 
                           n2141, ZN => n3899);
   U1325 : OAI22_X1 port map( A1 => n6027, A2 => n5939, B1 => n5424, B2 => 
                           n2142, ZN => n3900);
   U1326 : OAI22_X1 port map( A1 => n6030, A2 => n5940, B1 => n5424, B2 => 
                           n2143, ZN => n3901);
   U1327 : OAI22_X1 port map( A1 => n6033, A2 => n5941, B1 => n5424, B2 => 
                           n2144, ZN => n3902);
   U1328 : BUF_X1 port map( A => n5448, Z => n5450);
   U1329 : BUF_X1 port map( A => n5449, Z => n5451);
   U1330 : BUF_X1 port map( A => n4502, Z => n5532);
   U1331 : BUF_X1 port map( A => n4512, Z => n5523);
   U1332 : BUF_X1 port map( A => n4502, Z => n5533);
   U1333 : BUF_X1 port map( A => n4512, Z => n5524);
   U1334 : OAI22_X1 port map( A1 => n6061, A2 => n6034, B1 => n6058, B2 => 
                           n2074, ZN => n3999);
   U1335 : OAI22_X1 port map( A1 => n6061, A2 => n6037, B1 => n6059, B2 => 
                           n2075, ZN => n4000);
   U1336 : OAI22_X1 port map( A1 => n6061, A2 => n6040, B1 => n6058, B2 => 
                           n2076, ZN => n4001);
   U1337 : OAI22_X1 port map( A1 => n6060, A2 => n6043, B1 => n6059, B2 => 
                           n2077, ZN => n4002);
   U1338 : OAI22_X1 port map( A1 => n6060, A2 => n6046, B1 => n6058, B2 => 
                           n2080, ZN => n4003);
   U1339 : OAI22_X1 port map( A1 => n6060, A2 => n6049, B1 => n6059, B2 => 
                           n2112, ZN => n4004);
   U1340 : OAI22_X1 port map( A1 => n6060, A2 => n6052, B1 => n6058, B2 => 
                           n2114, ZN => n4005);
   U1341 : OAI22_X1 port map( A1 => n6060, A2 => n6055, B1 => n6059, B2 => 
                           n2115, ZN => n4006);
   U1342 : BUF_X1 port map( A => n5443, Z => n5445);
   U1343 : BUF_X1 port map( A => n5444, Z => n5446);
   U1344 : BUF_X1 port map( A => n5461, Z => n5463);
   U1345 : BUF_X1 port map( A => n5462, Z => n5464);
   U1346 : OAI22_X1 port map( A1 => n5963, A2 => n5854, B1 => n5398, B2 => 
                           n2479, ZN => n3591);
   U1347 : OAI22_X1 port map( A1 => n6034, A2 => n5706, B1 => n5347, B2 => 
                           n5304, ZN => n3071);
   U1348 : OAI22_X1 port map( A1 => n6037, A2 => n5706, B1 => n5347, B2 => 
                           n5305, ZN => n3072);
   U1349 : OAI22_X1 port map( A1 => n6040, A2 => n5707, B1 => n5347, B2 => 
                           n5309, ZN => n3073);
   U1350 : OAI22_X1 port map( A1 => n6043, A2 => n5707, B1 => n5347, B2 => 
                           n5306, ZN => n3074);
   U1351 : OAI22_X1 port map( A1 => n6046, A2 => n5702, B1 => n5347, B2 => 
                           n5307, ZN => n3075);
   U1352 : OAI22_X1 port map( A1 => n6049, A2 => n5702, B1 => n5347, B2 => 
                           n5310, ZN => n3076);
   U1353 : OAI22_X1 port map( A1 => n6052, A2 => n5705, B1 => n5347, B2 => 
                           n5297, ZN => n3077);
   U1354 : OAI22_X1 port map( A1 => n6055, A2 => n5704, B1 => n5347, B2 => 
                           n5298, ZN => n3078);
   U1355 : OAI22_X1 port map( A1 => n6034, A2 => n5715, B1 => n5350, B2 => 
                           n2832, ZN => n3103);
   U1356 : OAI22_X1 port map( A1 => n6037, A2 => n5715, B1 => n5350, B2 => 
                           n2851, ZN => n3104);
   U1357 : OAI22_X1 port map( A1 => n6040, A2 => n5716, B1 => n5350, B2 => 
                           n2870, ZN => n3105);
   U1358 : OAI22_X1 port map( A1 => n6043, A2 => n5716, B1 => n5350, B2 => 
                           n2889, ZN => n3106);
   U1359 : OAI22_X1 port map( A1 => n6046, A2 => n5711, B1 => n5350, B2 => 
                           n2908, ZN => n3107);
   U1360 : OAI22_X1 port map( A1 => n6049, A2 => n5711, B1 => n5350, B2 => 
                           n2919, ZN => n3108);
   U1361 : OAI22_X1 port map( A1 => n6052, A2 => n5714, B1 => n5350, B2 => 
                           n2920, ZN => n3109);
   U1362 : OAI22_X1 port map( A1 => n6055, A2 => n5713, B1 => n5350, B2 => 
                           n2921, ZN => n3110);
   U1363 : OAI22_X1 port map( A1 => n6034, A2 => n5724, B1 => n5353, B2 => 
                           n2640, ZN => n3135);
   U1364 : OAI22_X1 port map( A1 => n6037, A2 => n5724, B1 => n5353, B2 => 
                           n2641, ZN => n3136);
   U1365 : OAI22_X1 port map( A1 => n6040, A2 => n5725, B1 => n5353, B2 => 
                           n2642, ZN => n3137);
   U1366 : OAI22_X1 port map( A1 => n6043, A2 => n5725, B1 => n5353, B2 => 
                           n2643, ZN => n3138);
   U1367 : OAI22_X1 port map( A1 => n6046, A2 => n5720, B1 => n5353, B2 => 
                           n2644, ZN => n3139);
   U1368 : OAI22_X1 port map( A1 => n6049, A2 => n5720, B1 => n5353, B2 => 
                           n2645, ZN => n3140);
   U1369 : OAI22_X1 port map( A1 => n6052, A2 => n5723, B1 => n5353, B2 => 
                           n2646, ZN => n3141);
   U1370 : OAI22_X1 port map( A1 => n6055, A2 => n5722, B1 => n5353, B2 => 
                           n2647, ZN => n3142);
   U1371 : OAI22_X1 port map( A1 => n6034, A2 => n5734, B1 => n5356, B2 => 
                           n2379, ZN => n3167);
   U1372 : OAI22_X1 port map( A1 => n6037, A2 => n5734, B1 => n5356, B2 => 
                           n2380, ZN => n3168);
   U1373 : OAI22_X1 port map( A1 => n6040, A2 => n5730, B1 => n5356, B2 => 
                           n2384, ZN => n3169);
   U1374 : OAI22_X1 port map( A1 => n6043, A2 => n5734, B1 => n5356, B2 => 
                           n2381, ZN => n3170);
   U1375 : OAI22_X1 port map( A1 => n6046, A2 => n5728, B1 => n5356, B2 => 
                           n2382, ZN => n3171);
   U1376 : OAI22_X1 port map( A1 => n6049, A2 => n5728, B1 => n5356, B2 => 
                           n2385, ZN => n3172);
   U1377 : OAI22_X1 port map( A1 => n6052, A2 => n5728, B1 => n5356, B2 => 
                           n2372, ZN => n3173);
   U1378 : OAI22_X1 port map( A1 => n6055, A2 => n5730, B1 => n5356, B2 => 
                           n2373, ZN => n3174);
   U1379 : OAI22_X1 port map( A1 => n6035, A2 => n5743, B1 => n5359, B2 => 
                           n2480, ZN => n3199);
   U1380 : OAI22_X1 port map( A1 => n6038, A2 => n5743, B1 => n5359, B2 => 
                           n2481, ZN => n3200);
   U1381 : OAI22_X1 port map( A1 => n6041, A2 => n5743, B1 => n5359, B2 => 
                           n2482, ZN => n3201);
   U1382 : OAI22_X1 port map( A1 => n6044, A2 => n5743, B1 => n5359, B2 => 
                           n2483, ZN => n3202);
   U1383 : OAI22_X1 port map( A1 => n6047, A2 => n5737, B1 => n5359, B2 => 
                           n2484, ZN => n3203);
   U1384 : OAI22_X1 port map( A1 => n6050, A2 => n5737, B1 => n5359, B2 => 
                           n2485, ZN => n3204);
   U1385 : OAI22_X1 port map( A1 => n6053, A2 => n5737, B1 => n5359, B2 => 
                           n2486, ZN => n3205);
   U1386 : OAI22_X1 port map( A1 => n6056, A2 => n5739, B1 => n5359, B2 => 
                           n2487, ZN => n3206);
   U1387 : OAI22_X1 port map( A1 => n6034, A2 => n5751, B1 => n5362, B2 => 
                           n2580, ZN => n3231);
   U1388 : OAI22_X1 port map( A1 => n6037, A2 => n5751, B1 => n5362, B2 => 
                           n2581, ZN => n3232);
   U1389 : OAI22_X1 port map( A1 => n6040, A2 => n5752, B1 => n5362, B2 => 
                           n2582, ZN => n3233);
   U1390 : OAI22_X1 port map( A1 => n6043, A2 => n5752, B1 => n5362, B2 => 
                           n2583, ZN => n3234);
   U1391 : OAI22_X1 port map( A1 => n6046, A2 => n5747, B1 => n5362, B2 => 
                           n2584, ZN => n3235);
   U1392 : OAI22_X1 port map( A1 => n6049, A2 => n5747, B1 => n5362, B2 => 
                           n2585, ZN => n3236);
   U1393 : OAI22_X1 port map( A1 => n6052, A2 => n5750, B1 => n5362, B2 => 
                           n2586, ZN => n3237);
   U1394 : OAI22_X1 port map( A1 => n6055, A2 => n5749, B1 => n5362, B2 => 
                           n2587, ZN => n3238);
   U1395 : OAI22_X1 port map( A1 => n6034, A2 => n5760, B1 => n5365, B2 => 
                           n2505, ZN => n3263);
   U1396 : OAI22_X1 port map( A1 => n6037, A2 => n5760, B1 => n5365, B2 => 
                           n2506, ZN => n3264);
   U1397 : OAI22_X1 port map( A1 => n6040, A2 => n5761, B1 => n5365, B2 => 
                           n2521, ZN => n3265);
   U1398 : OAI22_X1 port map( A1 => n6043, A2 => n5761, B1 => n5365, B2 => 
                           n2507, ZN => n3266);
   U1399 : OAI22_X1 port map( A1 => n6046, A2 => n5756, B1 => n5365, B2 => 
                           n2508, ZN => n3267);
   U1400 : OAI22_X1 port map( A1 => n6049, A2 => n5756, B1 => n5365, B2 => 
                           n2522, ZN => n3268);
   U1401 : OAI22_X1 port map( A1 => n6052, A2 => n5759, B1 => n5365, B2 => 
                           n2509, ZN => n3269);
   U1402 : OAI22_X1 port map( A1 => n6055, A2 => n5758, B1 => n5365, B2 => 
                           n2510, ZN => n3270);
   U1403 : OAI22_X1 port map( A1 => n6034, A2 => n5770, B1 => n5368, B2 => 
                           n2170, ZN => n3295);
   U1404 : OAI22_X1 port map( A1 => n6037, A2 => n5770, B1 => n5368, B2 => 
                           n2171, ZN => n3296);
   U1405 : OAI22_X1 port map( A1 => n6040, A2 => n5766, B1 => n5368, B2 => 
                           n2188, ZN => n3297);
   U1406 : OAI22_X1 port map( A1 => n6043, A2 => n5770, B1 => n5368, B2 => 
                           n2172, ZN => n3298);
   U1407 : OAI22_X1 port map( A1 => n6046, A2 => n5764, B1 => n5368, B2 => 
                           n2173, ZN => n3299);
   U1408 : OAI22_X1 port map( A1 => n6049, A2 => n5764, B1 => n5368, B2 => 
                           n2189, ZN => n3300);
   U1409 : OAI22_X1 port map( A1 => n6052, A2 => n5764, B1 => n5368, B2 => 
                           n2174, ZN => n3301);
   U1410 : OAI22_X1 port map( A1 => n6055, A2 => n5766, B1 => n5368, B2 => 
                           n2175, ZN => n3302);
   U1411 : OAI22_X1 port map( A1 => n6034, A2 => n5778, B1 => n5371, B2 => 
                           n5271, ZN => n3327);
   U1412 : OAI22_X1 port map( A1 => n6037, A2 => n5778, B1 => n5371, B2 => 
                           n5272, ZN => n3328);
   U1413 : OAI22_X1 port map( A1 => n6040, A2 => n5779, B1 => n5371, B2 => 
                           n5273, ZN => n3329);
   U1414 : OAI22_X1 port map( A1 => n6043, A2 => n5779, B1 => n5371, B2 => 
                           n5274, ZN => n3330);
   U1415 : OAI22_X1 port map( A1 => n6046, A2 => n5774, B1 => n5371, B2 => 
                           n5275, ZN => n3331);
   U1416 : OAI22_X1 port map( A1 => n6049, A2 => n5774, B1 => n5371, B2 => 
                           n5276, ZN => n3332);
   U1417 : OAI22_X1 port map( A1 => n6052, A2 => n5777, B1 => n5371, B2 => 
                           n5277, ZN => n3333);
   U1418 : OAI22_X1 port map( A1 => n6055, A2 => n5776, B1 => n5371, B2 => 
                           n5278, ZN => n3334);
   U1419 : OAI22_X1 port map( A1 => n6034, A2 => n5787, B1 => n5374, B2 => 
                           n5239, ZN => n3359);
   U1420 : OAI22_X1 port map( A1 => n6037, A2 => n5787, B1 => n5374, B2 => 
                           n5240, ZN => n3360);
   U1421 : OAI22_X1 port map( A1 => n6040, A2 => n5788, B1 => n5374, B2 => 
                           n5241, ZN => n3361);
   U1422 : OAI22_X1 port map( A1 => n6043, A2 => n5788, B1 => n5374, B2 => 
                           n5242, ZN => n3362);
   U1423 : OAI22_X1 port map( A1 => n6046, A2 => n5783, B1 => n5374, B2 => 
                           n5243, ZN => n3363);
   U1424 : OAI22_X1 port map( A1 => n6049, A2 => n5783, B1 => n5374, B2 => 
                           n5244, ZN => n3364);
   U1425 : OAI22_X1 port map( A1 => n6052, A2 => n5786, B1 => n5374, B2 => 
                           n5245, ZN => n3365);
   U1426 : OAI22_X1 port map( A1 => n6055, A2 => n5785, B1 => n5374, B2 => 
                           n5246, ZN => n3366);
   U1427 : OAI22_X1 port map( A1 => n6035, A2 => n5796, B1 => n5377, B2 => 
                           n4090, ZN => n3391);
   U1428 : OAI22_X1 port map( A1 => n6038, A2 => n5796, B1 => n5377, B2 => 
                           n4109, ZN => n3392);
   U1429 : OAI22_X1 port map( A1 => n6041, A2 => n5797, B1 => n5377, B2 => 
                           n4185, ZN => n3393);
   U1430 : OAI22_X1 port map( A1 => n6044, A2 => n5797, B1 => n5377, B2 => 
                           n4128, ZN => n3394);
   U1431 : OAI22_X1 port map( A1 => n6047, A2 => n5792, B1 => n5377, B2 => 
                           n4147, ZN => n3395);
   U1432 : OAI22_X1 port map( A1 => n6050, A2 => n5792, B1 => n5377, B2 => 
                           n4204, ZN => n3396);
   U1433 : OAI22_X1 port map( A1 => n6053, A2 => n5795, B1 => n5377, B2 => 
                           n2947, ZN => n3397);
   U1434 : OAI22_X1 port map( A1 => n6056, A2 => n5794, B1 => n5377, B2 => 
                           n2948, ZN => n3398);
   U1435 : OAI22_X1 port map( A1 => n6035, A2 => n5806, B1 => n5380, B2 => 
                           n2414, ZN => n3423);
   U1436 : OAI22_X1 port map( A1 => n6038, A2 => n5806, B1 => n5380, B2 => 
                           n2415, ZN => n3424);
   U1437 : OAI22_X1 port map( A1 => n6041, A2 => n5802, B1 => n5380, B2 => 
                           n2416, ZN => n3425);
   U1438 : OAI22_X1 port map( A1 => n6044, A2 => n5806, B1 => n5380, B2 => 
                           n2417, ZN => n3426);
   U1439 : OAI22_X1 port map( A1 => n6047, A2 => n5800, B1 => n5380, B2 => 
                           n2418, ZN => n3427);
   U1440 : OAI22_X1 port map( A1 => n6050, A2 => n5800, B1 => n5380, B2 => 
                           n2419, ZN => n3428);
   U1441 : OAI22_X1 port map( A1 => n6053, A2 => n5800, B1 => n5380, B2 => 
                           n2420, ZN => n3429);
   U1442 : OAI22_X1 port map( A1 => n6056, A2 => n5802, B1 => n5380, B2 => 
                           n2421, ZN => n3430);
   U1443 : OAI22_X1 port map( A1 => n6035, A2 => n5815, B1 => n5383, B2 => 
                           n2213, ZN => n3455);
   U1444 : OAI22_X1 port map( A1 => n6038, A2 => n5815, B1 => n5383, B2 => 
                           n2214, ZN => n3456);
   U1445 : OAI22_X1 port map( A1 => n6041, A2 => n5815, B1 => n5383, B2 => 
                           n2215, ZN => n3457);
   U1446 : OAI22_X1 port map( A1 => n6044, A2 => n5815, B1 => n5383, B2 => 
                           n2216, ZN => n3458);
   U1447 : OAI22_X1 port map( A1 => n6047, A2 => n5809, B1 => n5383, B2 => 
                           n2219, ZN => n3459);
   U1448 : OAI22_X1 port map( A1 => n6050, A2 => n5809, B1 => n5383, B2 => 
                           n2220, ZN => n3460);
   U1449 : OAI22_X1 port map( A1 => n6053, A2 => n5809, B1 => n5383, B2 => 
                           n2221, ZN => n3461);
   U1450 : OAI22_X1 port map( A1 => n6056, A2 => n5811, B1 => n5383, B2 => 
                           n2222, ZN => n3462);
   U1451 : OAI22_X1 port map( A1 => n6035, A2 => n5824, B1 => n5386, B2 => 
                           n2439, ZN => n3487);
   U1452 : OAI22_X1 port map( A1 => n6038, A2 => n5824, B1 => n5386, B2 => 
                           n2440, ZN => n3488);
   U1453 : OAI22_X1 port map( A1 => n6041, A2 => n5824, B1 => n5386, B2 => 
                           n2453, ZN => n3489);
   U1454 : OAI22_X1 port map( A1 => n6044, A2 => n5824, B1 => n5386, B2 => 
                           n2441, ZN => n3490);
   U1455 : OAI22_X1 port map( A1 => n6047, A2 => n5818, B1 => n5386, B2 => 
                           n2442, ZN => n3491);
   U1456 : OAI22_X1 port map( A1 => n6050, A2 => n5818, B1 => n5386, B2 => 
                           n2454, ZN => n3492);
   U1457 : OAI22_X1 port map( A1 => n6053, A2 => n5818, B1 => n5386, B2 => 
                           n2443, ZN => n3493);
   U1458 : OAI22_X1 port map( A1 => n6056, A2 => n5820, B1 => n5386, B2 => 
                           n2444, ZN => n3494);
   U1459 : OAI22_X1 port map( A1 => n6035, A2 => n5832, B1 => n5389, B2 => 
                           n5199, ZN => n3519);
   U1460 : OAI22_X1 port map( A1 => n6038, A2 => n5832, B1 => n5389, B2 => 
                           n5200, ZN => n3520);
   U1461 : OAI22_X1 port map( A1 => n6041, A2 => n5833, B1 => n5389, B2 => 
                           n5213, ZN => n3521);
   U1462 : OAI22_X1 port map( A1 => n6044, A2 => n5833, B1 => n5389, B2 => 
                           n5201, ZN => n3522);
   U1463 : OAI22_X1 port map( A1 => n6047, A2 => n5828, B1 => n5389, B2 => 
                           n5202, ZN => n3523);
   U1464 : OAI22_X1 port map( A1 => n6050, A2 => n5828, B1 => n5389, B2 => 
                           n5214, ZN => n3524);
   U1465 : OAI22_X1 port map( A1 => n6053, A2 => n5831, B1 => n5389, B2 => 
                           n5203, ZN => n3525);
   U1466 : OAI22_X1 port map( A1 => n6056, A2 => n5830, B1 => n5389, B2 => 
                           n5204, ZN => n3526);
   U1467 : OAI22_X1 port map( A1 => n6035, A2 => n5851, B1 => n5395, B2 => 
                           n2345, ZN => n3583);
   U1468 : OAI22_X1 port map( A1 => n6038, A2 => n5851, B1 => n5395, B2 => 
                           n2346, ZN => n3584);
   U1469 : OAI22_X1 port map( A1 => n6041, A2 => n5851, B1 => n5395, B2 => 
                           n2347, ZN => n3585);
   U1470 : OAI22_X1 port map( A1 => n6044, A2 => n5851, B1 => n5395, B2 => 
                           n2348, ZN => n3586);
   U1471 : OAI22_X1 port map( A1 => n6047, A2 => n5845, B1 => n5395, B2 => 
                           n2349, ZN => n3587);
   U1472 : OAI22_X1 port map( A1 => n6050, A2 => n5845, B1 => n5395, B2 => 
                           n2350, ZN => n3588);
   U1473 : OAI22_X1 port map( A1 => n6053, A2 => n5845, B1 => n5395, B2 => 
                           n2351, ZN => n3589);
   U1474 : OAI22_X1 port map( A1 => n6056, A2 => n5847, B1 => n5395, B2 => 
                           n2352, ZN => n3590);
   U1475 : OAI22_X1 port map( A1 => n6035, A2 => n5869, B1 => n5401, B2 => 
                           n2311, ZN => n3647);
   U1476 : OAI22_X1 port map( A1 => n6038, A2 => n5869, B1 => n5401, B2 => 
                           n2312, ZN => n3648);
   U1477 : OAI22_X1 port map( A1 => n6041, A2 => n5869, B1 => n5401, B2 => 
                           n2313, ZN => n3649);
   U1478 : OAI22_X1 port map( A1 => n6044, A2 => n5869, B1 => n5401, B2 => 
                           n2314, ZN => n3650);
   U1479 : OAI22_X1 port map( A1 => n6047, A2 => n5863, B1 => n5401, B2 => 
                           n2315, ZN => n3651);
   U1480 : OAI22_X1 port map( A1 => n6050, A2 => n5863, B1 => n5401, B2 => 
                           n2316, ZN => n3652);
   U1481 : OAI22_X1 port map( A1 => n6053, A2 => n5863, B1 => n5401, B2 => 
                           n2317, ZN => n3653);
   U1482 : OAI22_X1 port map( A1 => n6056, A2 => n5865, B1 => n5401, B2 => 
                           n2318, ZN => n3654);
   U1483 : OAI22_X1 port map( A1 => n6035, A2 => n5877, B1 => n5404, B2 => 
                           n2922, ZN => n3679);
   U1484 : OAI22_X1 port map( A1 => n6038, A2 => n5877, B1 => n5404, B2 => 
                           n2923, ZN => n3680);
   U1485 : OAI22_X1 port map( A1 => n6041, A2 => n5878, B1 => n5404, B2 => 
                           n2924, ZN => n3681);
   U1486 : OAI22_X1 port map( A1 => n6044, A2 => n5878, B1 => n5404, B2 => 
                           n2925, ZN => n3682);
   U1487 : OAI22_X1 port map( A1 => n6047, A2 => n5872, B1 => n5404, B2 => 
                           n2926, ZN => n3683);
   U1488 : OAI22_X1 port map( A1 => n6050, A2 => n5872, B1 => n5404, B2 => 
                           n2927, ZN => n3684);
   U1489 : OAI22_X1 port map( A1 => n6053, A2 => n5876, B1 => n5404, B2 => 
                           n2928, ZN => n3685);
   U1490 : OAI22_X1 port map( A1 => n6056, A2 => n5875, B1 => n5404, B2 => 
                           n2929, ZN => n3686);
   U1491 : OAI22_X1 port map( A1 => n6035, A2 => n5886, B1 => n5407, B2 => 
                           n2243, ZN => n3711);
   U1492 : OAI22_X1 port map( A1 => n6038, A2 => n5887, B1 => n5407, B2 => 
                           n2244, ZN => n3712);
   U1493 : OAI22_X1 port map( A1 => n6041, A2 => n5886, B1 => n5407, B2 => 
                           n2118, ZN => n3713);
   U1494 : OAI22_X1 port map( A1 => n6044, A2 => n5887, B1 => n5407, B2 => 
                           n2117, ZN => n3714);
   U1495 : OAI22_X1 port map( A1 => n6047, A2 => n5881, B1 => n5407, B2 => 
                           n2245, ZN => n3715);
   U1496 : OAI22_X1 port map( A1 => n6050, A2 => n5881, B1 => n5407, B2 => 
                           n2257, ZN => n3716);
   U1497 : OAI22_X1 port map( A1 => n6053, A2 => n5886, B1 => n5407, B2 => 
                           n2246, ZN => n3717);
   U1498 : OAI22_X1 port map( A1 => n6056, A2 => n5884, B1 => n5407, B2 => 
                           n2247, ZN => n3718);
   U1499 : OAI22_X1 port map( A1 => n6035, A2 => n5895, B1 => n5410, B2 => 
                           n5114, ZN => n3743);
   U1500 : OAI22_X1 port map( A1 => n6038, A2 => n5895, B1 => n5410, B2 => 
                           n5115, ZN => n3744);
   U1501 : OAI22_X1 port map( A1 => n6041, A2 => n5896, B1 => n5410, B2 => 
                           n5116, ZN => n3745);
   U1502 : OAI22_X1 port map( A1 => n6044, A2 => n5896, B1 => n5410, B2 => 
                           n5117, ZN => n3746);
   U1503 : OAI22_X1 port map( A1 => n6047, A2 => n5891, B1 => n5410, B2 => 
                           n5118, ZN => n3747);
   U1504 : OAI22_X1 port map( A1 => n6050, A2 => n5891, B1 => n5410, B2 => 
                           n5119, ZN => n3748);
   U1505 : OAI22_X1 port map( A1 => n6053, A2 => n5894, B1 => n5410, B2 => 
                           n5120, ZN => n3749);
   U1506 : OAI22_X1 port map( A1 => n6056, A2 => n5893, B1 => n5410, B2 => 
                           n5121, ZN => n3750);
   U1507 : OAI22_X1 port map( A1 => n6035, A2 => n5913, B1 => n5416, B2 => 
                           n5139, ZN => n3807);
   U1508 : OAI22_X1 port map( A1 => n6038, A2 => n5913, B1 => n5416, B2 => 
                           n5140, ZN => n3808);
   U1509 : OAI22_X1 port map( A1 => n6041, A2 => n5914, B1 => n5416, B2 => 
                           n2386, ZN => n3809);
   U1510 : OAI22_X1 port map( A1 => n6044, A2 => n5914, B1 => n5416, B2 => 
                           n5141, ZN => n3810);
   U1511 : OAI22_X1 port map( A1 => n6047, A2 => n5908, B1 => n5416, B2 => 
                           n5142, ZN => n3811);
   U1512 : OAI22_X1 port map( A1 => n6050, A2 => n5908, B1 => n5416, B2 => 
                           n5153, ZN => n3812);
   U1513 : OAI22_X1 port map( A1 => n6053, A2 => n5913, B1 => n5416, B2 => 
                           n5143, ZN => n3813);
   U1514 : OAI22_X1 port map( A1 => n6056, A2 => n5911, B1 => n5416, B2 => 
                           n5144, ZN => n3814);
   U1515 : OAI22_X1 port map( A1 => n6036, A2 => n5923, B1 => n5419, B2 => 
                           n2281, ZN => n3839);
   U1516 : OAI22_X1 port map( A1 => n6039, A2 => n5923, B1 => n5419, B2 => 
                           n2282, ZN => n3840);
   U1517 : OAI22_X1 port map( A1 => n6042, A2 => n5923, B1 => n5419, B2 => 
                           n2119, ZN => n3841);
   U1518 : OAI22_X1 port map( A1 => n6045, A2 => n5922, B1 => n5419, B2 => 
                           n2120, ZN => n3842);
   U1519 : OAI22_X1 port map( A1 => n6048, A2 => n5917, B1 => n5419, B2 => 
                           n2283, ZN => n3843);
   U1520 : OAI22_X1 port map( A1 => n6051, A2 => n5917, B1 => n5419, B2 => 
                           n2284, ZN => n3844);
   U1521 : OAI22_X1 port map( A1 => n6054, A2 => n5922, B1 => n5419, B2 => 
                           n2285, ZN => n3845);
   U1522 : OAI22_X1 port map( A1 => n6057, A2 => n5920, B1 => n5419, B2 => 
                           n2287, ZN => n3846);
   U1523 : OAI22_X1 port map( A1 => n6036, A2 => n5941, B1 => n5425, B2 => 
                           n2145, ZN => n3903);
   U1524 : OAI22_X1 port map( A1 => n6039, A2 => n5941, B1 => n5425, B2 => 
                           n2146, ZN => n3904);
   U1525 : OAI22_X1 port map( A1 => n6042, A2 => n5937, B1 => n5425, B2 => 
                           n2151, ZN => n3905);
   U1526 : OAI22_X1 port map( A1 => n6045, A2 => n5941, B1 => n5425, B2 => 
                           n2148, ZN => n3906);
   U1527 : OAI22_X1 port map( A1 => n6048, A2 => n5935, B1 => n5425, B2 => 
                           n2149, ZN => n3907);
   U1528 : OAI22_X1 port map( A1 => n6051, A2 => n5935, B1 => n5425, B2 => 
                           n2152, ZN => n3908);
   U1529 : OAI22_X1 port map( A1 => n6054, A2 => n5935, B1 => n5425, B2 => 
                           n2138, ZN => n3909);
   U1530 : OAI22_X1 port map( A1 => n6057, A2 => n5937, B1 => n5425, B2 => 
                           n2139, ZN => n3910);
   U1531 : OAI22_X1 port map( A1 => n6066, A2 => n5962, B1 => n6058, B2 => 
                           n2153, ZN => n3975);
   U1532 : OAI22_X1 port map( A1 => n6066, A2 => n5965, B1 => n6058, B2 => 
                           n2051, ZN => n3976);
   U1533 : OAI22_X1 port map( A1 => n6065, A2 => n5968, B1 => n6058, B2 => 
                           n2052, ZN => n3977);
   U1534 : OAI22_X1 port map( A1 => n6065, A2 => n5971, B1 => n6058, B2 => 
                           n2053, ZN => n3978);
   U1535 : OAI22_X1 port map( A1 => n6065, A2 => n5974, B1 => n6058, B2 => 
                           n2054, ZN => n3979);
   U1536 : OAI22_X1 port map( A1 => n6065, A2 => n5977, B1 => n6058, B2 => 
                           n2055, ZN => n3980);
   U1537 : OAI22_X1 port map( A1 => n6065, A2 => n5980, B1 => n6058, B2 => 
                           n2056, ZN => n3981);
   U1538 : OAI22_X1 port map( A1 => n6064, A2 => n5983, B1 => n6058, B2 => 
                           n2057, ZN => n3982);
   U1539 : OAI22_X1 port map( A1 => n6064, A2 => n5986, B1 => n6058, B2 => 
                           n2058, ZN => n3983);
   U1540 : OAI22_X1 port map( A1 => n6064, A2 => n5989, B1 => n6058, B2 => 
                           n2059, ZN => n3984);
   U1541 : OAI22_X1 port map( A1 => n6064, A2 => n5992, B1 => n6058, B2 => 
                           n2060, ZN => n3985);
   U1542 : OAI22_X1 port map( A1 => n6064, A2 => n5995, B1 => n6058, B2 => 
                           n2061, ZN => n3986);
   U1543 : OAI22_X1 port map( A1 => n6063, A2 => n5998, B1 => n6059, B2 => 
                           n2062, ZN => n3987);
   U1544 : OAI22_X1 port map( A1 => n6063, A2 => n6001, B1 => n6059, B2 => 
                           n2063, ZN => n3988);
   U1545 : OAI22_X1 port map( A1 => n6063, A2 => n6004, B1 => n6059, B2 => 
                           n2064, ZN => n3989);
   U1546 : OAI22_X1 port map( A1 => n6063, A2 => n6007, B1 => n6059, B2 => 
                           n2065, ZN => n3990);
   U1547 : OAI22_X1 port map( A1 => n6063, A2 => n6010, B1 => n6059, B2 => 
                           n2066, ZN => n3991);
   U1548 : OAI22_X1 port map( A1 => n6062, A2 => n6013, B1 => n6059, B2 => 
                           n2067, ZN => n3992);
   U1549 : OAI22_X1 port map( A1 => n6062, A2 => n6016, B1 => n6059, B2 => 
                           n2068, ZN => n3993);
   U1550 : OAI22_X1 port map( A1 => n6062, A2 => n6019, B1 => n6059, B2 => 
                           n2069, ZN => n3994);
   U1551 : OAI22_X1 port map( A1 => n6062, A2 => n6022, B1 => n6059, B2 => 
                           n2070, ZN => n3995);
   U1552 : OAI22_X1 port map( A1 => n6062, A2 => n6025, B1 => n6059, B2 => 
                           n2071, ZN => n3996);
   U1553 : OAI22_X1 port map( A1 => n6061, A2 => n6028, B1 => n6059, B2 => 
                           n2072, ZN => n3997);
   U1554 : OAI22_X1 port map( A1 => n6061, A2 => n6031, B1 => n6059, B2 => 
                           n2073, ZN => n3998);
   U1555 : BUF_X1 port map( A => n5456, Z => n5458);
   U1556 : BUF_X1 port map( A => n5457, Z => n5459);
   U1557 : OAI22_X1 port map( A1 => n6041, A2 => n5841, B1 => n5392, B2 => 
                           n2648, ZN => n3553);
   U1558 : OAI22_X1 port map( A1 => n6044, A2 => n5841, B1 => n5392, B2 => 
                           n2649, ZN => n3554);
   U1559 : OAI22_X1 port map( A1 => n6047, A2 => n5842, B1 => n5392, B2 => 
                           n2650, ZN => n3555);
   U1560 : OAI22_X1 port map( A1 => n6050, A2 => n5842, B1 => n5392, B2 => 
                           n2651, ZN => n3556);
   U1561 : OAI22_X1 port map( A1 => n6053, A2 => n5836, B1 => n5392, B2 => 
                           n2652, ZN => n3557);
   U1562 : OAI22_X1 port map( A1 => n6056, A2 => n5841, B1 => n5392, B2 => 
                           n2653, ZN => n3558);
   U1563 : OAI22_X1 port map( A1 => n6042, A2 => n5931, B1 => n5422, B2 => 
                           n2551, ZN => n3873);
   U1564 : OAI22_X1 port map( A1 => n6045, A2 => n5931, B1 => n5422, B2 => 
                           n2552, ZN => n3874);
   U1565 : OAI22_X1 port map( A1 => n6048, A2 => n5932, B1 => n5422, B2 => 
                           n2553, ZN => n3875);
   U1566 : OAI22_X1 port map( A1 => n6051, A2 => n5932, B1 => n5422, B2 => 
                           n2554, ZN => n3876);
   U1567 : OAI22_X1 port map( A1 => n6054, A2 => n5926, B1 => n5422, B2 => 
                           n2545, ZN => n3877);
   U1568 : OAI22_X1 port map( A1 => n6057, A2 => n5932, B1 => n5422, B2 => 
                           n2546, ZN => n3878);
   U1569 : BUF_X1 port map( A => n4501, Z => n5452);
   U1570 : OAI22_X1 port map( A1 => n5962, A2 => n5942, B1 => n5951, B2 => 
                           n5123, ZN => n3911);
   U1571 : OAI22_X1 port map( A1 => n5965, A2 => n5942, B1 => n5951, B2 => 
                           n5154, ZN => n3912);
   U1572 : OAI22_X1 port map( A1 => n5968, A2 => n5942, B1 => n5951, B2 => 
                           n5155, ZN => n3913);
   U1573 : OAI22_X1 port map( A1 => n5971, A2 => n5942, B1 => n5951, B2 => 
                           n5156, ZN => n3914);
   U1574 : OAI22_X1 port map( A1 => n5974, A2 => n5942, B1 => n5950, B2 => 
                           n5157, ZN => n3915);
   U1575 : OAI22_X1 port map( A1 => n5977, A2 => n5942, B1 => n5950, B2 => 
                           n5158, ZN => n3916);
   U1576 : OAI22_X1 port map( A1 => n5980, A2 => n5942, B1 => n5950, B2 => 
                           n5159, ZN => n3917);
   U1577 : OAI22_X1 port map( A1 => n5983, A2 => n5942, B1 => n5950, B2 => 
                           n5160, ZN => n3918);
   U1578 : OAI22_X1 port map( A1 => n5986, A2 => n5942, B1 => n5949, B2 => 
                           n5161, ZN => n3919);
   U1579 : OAI22_X1 port map( A1 => n5989, A2 => n5942, B1 => n5949, B2 => 
                           n5162, ZN => n3920);
   U1580 : OAI22_X1 port map( A1 => n5992, A2 => n5942, B1 => n5949, B2 => 
                           n5163, ZN => n3921);
   U1581 : OAI22_X1 port map( A1 => n5995, A2 => n5942, B1 => n5949, B2 => 
                           n5164, ZN => n3922);
   U1582 : OAI22_X1 port map( A1 => n5998, A2 => n5943, B1 => n5948, B2 => 
                           n5165, ZN => n3923);
   U1583 : OAI22_X1 port map( A1 => n6001, A2 => n5943, B1 => n5948, B2 => 
                           n5166, ZN => n3924);
   U1584 : OAI22_X1 port map( A1 => n6004, A2 => n5943, B1 => n5948, B2 => 
                           n5167, ZN => n3925);
   U1585 : OAI22_X1 port map( A1 => n6007, A2 => n5943, B1 => n5948, B2 => 
                           n5168, ZN => n3926);
   U1586 : OAI22_X1 port map( A1 => n6010, A2 => n5943, B1 => n5947, B2 => 
                           n5169, ZN => n3927);
   U1587 : OAI22_X1 port map( A1 => n6013, A2 => n5943, B1 => n5947, B2 => 
                           n5170, ZN => n3928);
   U1588 : OAI22_X1 port map( A1 => n6016, A2 => n5943, B1 => n5947, B2 => 
                           n5171, ZN => n3929);
   U1589 : OAI22_X1 port map( A1 => n6019, A2 => n5943, B1 => n5947, B2 => 
                           n5172, ZN => n3930);
   U1590 : OAI22_X1 port map( A1 => n6022, A2 => n5943, B1 => n5946, B2 => 
                           n5173, ZN => n3931);
   U1591 : OAI22_X1 port map( A1 => n6025, A2 => n5943, B1 => n5946, B2 => 
                           n5174, ZN => n3932);
   U1592 : OAI22_X1 port map( A1 => n6028, A2 => n5943, B1 => n5946, B2 => 
                           n5175, ZN => n3933);
   U1593 : OAI22_X1 port map( A1 => n6031, A2 => n5943, B1 => n5946, B2 => 
                           n5176, ZN => n3934);
   U1594 : OAI22_X1 port map( A1 => n6034, A2 => n5942, B1 => n5945, B2 => 
                           n5177, ZN => n3935);
   U1595 : OAI22_X1 port map( A1 => n6037, A2 => n5943, B1 => n5945, B2 => 
                           n5178, ZN => n3936);
   U1596 : OAI22_X1 port map( A1 => n6040, A2 => n5942, B1 => n5945, B2 => 
                           n5179, ZN => n3937);
   U1597 : OAI22_X1 port map( A1 => n6043, A2 => n5943, B1 => n5945, B2 => 
                           n2388, ZN => n3938);
   U1598 : OAI22_X1 port map( A1 => n6046, A2 => n5942, B1 => n5944, B2 => 
                           n5180, ZN => n3939);
   U1599 : OAI22_X1 port map( A1 => n6049, A2 => n5943, B1 => n5944, B2 => 
                           n5181, ZN => n3940);
   U1600 : OAI22_X1 port map( A1 => n6052, A2 => n5942, B1 => n5944, B2 => 
                           n5182, ZN => n3941);
   U1601 : OAI22_X1 port map( A1 => n6055, A2 => n5943, B1 => n5944, B2 => 
                           n5183, ZN => n3942);
   U1602 : BUF_X1 port map( A => n5484, Z => n5486);
   U1603 : BUF_X1 port map( A => n4502, Z => n5534);
   U1604 : BUF_X1 port map( A => n4512, Z => n5525);
   U1605 : BUF_X1 port map( A => n4504, Z => n5447);
   U1606 : BUF_X1 port map( A => n2704, Z => n5696);
   U1607 : BUF_X1 port map( A => n2704, Z => n5697);
   U1608 : BUF_X1 port map( A => n5485, Z => n5487);
   U1609 : BUF_X1 port map( A => n5438, Z => n5440);
   U1610 : BUF_X1 port map( A => n5439, Z => n5441);
   U1611 : NAND2_X1 port map( A1 => n2629, A2 => n1730, ZN => n2665);
   U1612 : NAND2_X1 port map( A1 => n2492, A2 => n1730, ZN => n2527);
   U1613 : NAND2_X1 port map( A1 => n2355, A2 => n1730, ZN => n2390);
   U1614 : NAND2_X1 port map( A1 => n2217, A2 => n1730, ZN => n2252);
   U1615 : NAND2_X1 port map( A1 => n2078, A2 => n1730, ZN => n2113);
   U1616 : NAND2_X1 port map( A1 => n1941, A2 => n1730, ZN => n1976);
   U1617 : NAND2_X1 port map( A1 => n1804, A2 => n1730, ZN => n1839);
   U1618 : NAND2_X1 port map( A1 => n5080, A2 => n5084, ZN => n4491);
   U1619 : NAND2_X1 port map( A1 => n2078, A2 => n1694, ZN => n2081);
   U1620 : NAND2_X1 port map( A1 => n2629, A2 => n1694, ZN => n2630);
   U1621 : NAND2_X1 port map( A1 => n2492, A2 => n1694, ZN => n2493);
   U1622 : NAND2_X1 port map( A1 => n2355, A2 => n1694, ZN => n2356);
   U1623 : NAND2_X1 port map( A1 => n2217, A2 => n1694, ZN => n2218);
   U1624 : NAND2_X1 port map( A1 => n1941, A2 => n1694, ZN => n1942);
   U1625 : NAND2_X1 port map( A1 => n1804, A2 => n1694, ZN => n1805);
   U1626 : BUF_X1 port map( A => n4481, Z => n5465);
   U1627 : NAND2_X1 port map( A1 => n2492, A2 => n1765, ZN => n2561);
   U1628 : NAND2_X1 port map( A1 => n2355, A2 => n1765, ZN => n2424);
   U1629 : NAND2_X1 port map( A1 => n2078, A2 => n1765, ZN => n2147);
   U1630 : NAND2_X1 port map( A1 => n1941, A2 => n1765, ZN => n2010);
   U1631 : NAND2_X1 port map( A1 => n1804, A2 => n1765, ZN => n1873);
   U1632 : NAND2_X1 port map( A1 => n1941, A2 => n1803, ZN => n1909);
   U1633 : NAND2_X1 port map( A1 => n2629, A2 => n1803, ZN => n2595);
   U1634 : NAND2_X1 port map( A1 => n2492, A2 => n1803, ZN => n2458);
   U1635 : NAND2_X1 port map( A1 => n2355, A2 => n1803, ZN => n2321);
   U1636 : NAND2_X1 port map( A1 => n2217, A2 => n1803, ZN => n2183);
   U1637 : NAND2_X1 port map( A1 => n2078, A2 => n1803, ZN => n2044);
   U1638 : BUF_X1 port map( A => n4480, Z => n5460);
   U1639 : BUF_X1 port map( A => n2704, Z => n5698);
   U1640 : BUF_X1 port map( A => n2749, Z => n5488);
   U1641 : BUF_X1 port map( A => n4506, Z => n5442);
   U1642 : AND3_X1 port map( A1 => n1766, A2 => n1767, A3 => n2320, ZN => n2217
                           );
   U1643 : AND3_X1 port map( A1 => n5078, A2 => n5503, A3 => n5079, ZN => n4484
                           );
   U1644 : AND3_X1 port map( A1 => n5078, A2 => n5503, A3 => n5085, ZN => n4508
                           );
   U1645 : AND3_X1 port map( A1 => n5067, A2 => n5506, A3 => n5070, ZN => n4478
                           );
   U1646 : AND3_X1 port map( A1 => n5067, A2 => n5504, A3 => n5085, ZN => n4513
                           );
   U1647 : AND2_X1 port map( A1 => n5080, A2 => n5070, ZN => n4494);
   U1648 : AND3_X1 port map( A1 => n1766, A2 => n1767, A3 => n1768, ZN => n1695
                           );
   U1649 : AND2_X1 port map( A1 => n5500, A2 => n5100, ZN => n5068);
   U1650 : NAND4_X1 port map( A1 => n5072, A2 => n5101, A3 => n5071, A4 => 
                           n5102, ZN => n5100);
   U1651 : NOR3_X1 port map( A1 => n5075, A2 => n2182, A3 => n5074, ZN => n5102
                           );
   U1652 : INV_X1 port map( A => n5076, ZN => n5101);
   U1653 : AND4_X1 port map( A1 => n5086, A2 => n5078, A3 => n5503, A4 => n5087
                           , ZN => n4509);
   U1654 : AND2_X1 port map( A1 => n5080, A2 => n5085, ZN => n5563);
   U1655 : AND2_X1 port map( A1 => n5080, A2 => n5085, ZN => n5564);
   U1656 : AND2_X1 port map( A1 => n5080, A2 => n5085, ZN => n4488);
   U1657 : BUF_X1 port map( A => n1690, Z => n5967);
   U1658 : BUF_X1 port map( A => n1688, Z => n5970);
   U1659 : BUF_X1 port map( A => n1686, Z => n5973);
   U1660 : BUF_X1 port map( A => n1684, Z => n5976);
   U1661 : BUF_X1 port map( A => n1682, Z => n5979);
   U1662 : BUF_X1 port map( A => n1680, Z => n5982);
   U1663 : BUF_X1 port map( A => n1678, Z => n5985);
   U1664 : BUF_X1 port map( A => n1676, Z => n5988);
   U1665 : BUF_X1 port map( A => n1674, Z => n5991);
   U1666 : BUF_X1 port map( A => n1672, Z => n5994);
   U1667 : BUF_X1 port map( A => n1670, Z => n5997);
   U1668 : BUF_X1 port map( A => n1668, Z => n6000);
   U1669 : BUF_X1 port map( A => n1666, Z => n6003);
   U1670 : BUF_X1 port map( A => n1664, Z => n6006);
   U1671 : BUF_X1 port map( A => n1662, Z => n6009);
   U1672 : BUF_X1 port map( A => n1660, Z => n6012);
   U1673 : BUF_X1 port map( A => n1658, Z => n6015);
   U1674 : BUF_X1 port map( A => n1656, Z => n6018);
   U1675 : BUF_X1 port map( A => n1654, Z => n6021);
   U1676 : BUF_X1 port map( A => n1652, Z => n6024);
   U1677 : BUF_X1 port map( A => n1650, Z => n6027);
   U1678 : BUF_X1 port map( A => n1648, Z => n6030);
   U1679 : BUF_X1 port map( A => n1646, Z => n6033);
   U1680 : BUF_X1 port map( A => n1644, Z => n6036);
   U1681 : BUF_X1 port map( A => n1642, Z => n6039);
   U1682 : BUF_X1 port map( A => n1640, Z => n6042);
   U1683 : BUF_X1 port map( A => n1638, Z => n6045);
   U1684 : BUF_X1 port map( A => n1636, Z => n6048);
   U1685 : BUF_X1 port map( A => n1634, Z => n6051);
   U1686 : BUF_X1 port map( A => n1632, Z => n6054);
   U1687 : BUF_X1 port map( A => n1629, Z => n6057);
   U1688 : OAI22_X1 port map( A1 => n2547, A2 => n5675, B1 => n2309, B2 => 
                           n5682, ZN => n4011);
   U1689 : OAI22_X1 port map( A1 => n2548, A2 => n5676, B1 => n2310, B2 => 
                           n2744, ZN => n2905);
   U1690 : OAI22_X1 port map( A1 => n2549, A2 => n5675, B1 => n2311, B2 => 
                           n5681, ZN => n2886);
   U1691 : OAI22_X1 port map( A1 => n2550, A2 => n5676, B1 => n2312, B2 => 
                           n5682, ZN => n2867);
   U1692 : OAI22_X1 port map( A1 => n2551, A2 => n5675, B1 => n2313, B2 => 
                           n2744, ZN => n2848);
   U1693 : OAI22_X1 port map( A1 => n2552, A2 => n5676, B1 => n2314, B2 => 
                           n5681, ZN => n2829);
   U1694 : OAI22_X1 port map( A1 => n2553, A2 => n5675, B1 => n2315, B2 => 
                           n5682, ZN => n2810);
   U1695 : OAI22_X1 port map( A1 => n2554, A2 => n5676, B1 => n2316, B2 => 
                           n2744, ZN => n2791);
   U1696 : BUF_X1 port map( A => n1692, Z => n5964);
   U1697 : NOR2_X1 port map( A1 => n4441, A2 => n4458, ZN => n4443);
   U1698 : AND2_X1 port map( A1 => n4429, A2 => n4439, ZN => n5655);
   U1699 : AND2_X1 port map( A1 => n4429, A2 => n4439, ZN => n5656);
   U1700 : AND2_X1 port map( A1 => n4429, A2 => n4439, ZN => n2723);
   U1701 : BUF_X1 port map( A => n2752, Z => n5466);
   U1702 : AND2_X1 port map( A1 => n4430, A2 => n4443, ZN => n2738);
   U1703 : AND3_X1 port map( A1 => n4433, A2 => n4434, A3 => n4439, ZN => n2733
                           );
   U1704 : AND2_X1 port map( A1 => n4426, A2 => n4439, ZN => n2739);
   U1705 : AND2_X1 port map( A1 => n4428, A2 => n4443, ZN => n2724);
   U1706 : BUF_X1 port map( A => n5489, Z => n5491);
   U1707 : BUF_X1 port map( A => n5489, Z => n5494);
   U1708 : BUF_X1 port map( A => n5490, Z => n5496);
   U1709 : BUF_X1 port map( A => n5490, Z => n5497);
   U1710 : BUF_X1 port map( A => n5490, Z => n5495);
   U1711 : BUF_X1 port map( A => n5490, Z => n5498);
   U1712 : BUF_X1 port map( A => n4476, Z => n5499);
   U1713 : BUF_X1 port map( A => n5489, Z => n5492);
   U1714 : BUF_X1 port map( A => n5489, Z => n5493);
   U1715 : BUF_X1 port map( A => n4476, Z => n5500);
   U1716 : BUF_X1 port map( A => rst, Z => n6073);
   U1717 : NOR3_X1 port map( A1 => n4461, A2 => n4434, A3 => n4459, ZN => n4438
                           );
   U1718 : NOR3_X1 port map( A1 => n5096, A2 => n5087, A3 => n5097, ZN => n5069
                           );
   U1719 : NAND2_X1 port map( A1 => n4429, A2 => n4443, ZN => n5642);
   U1720 : NAND2_X1 port map( A1 => n4429, A2 => n4443, ZN => n5643);
   U1721 : NAND2_X1 port map( A1 => n4429, A2 => n4443, ZN => n2725);
   U1722 : AND3_X1 port map( A1 => n4458, A2 => n4441, A3 => n4438, ZN => n5646
                           );
   U1723 : AND3_X1 port map( A1 => n4458, A2 => n4441, A3 => n4438, ZN => n5647
                           );
   U1724 : AND3_X1 port map( A1 => n4458, A2 => n4441, A3 => n4438, ZN => n2729
                           );
   U1725 : NAND2_X1 port map( A1 => n4428, A2 => n4439, ZN => n5648);
   U1726 : NAND2_X1 port map( A1 => n4428, A2 => n4439, ZN => n2720);
   U1727 : NAND2_X1 port map( A1 => n4439, A2 => n4435, ZN => n2730);
   U1728 : NAND2_X1 port map( A1 => n4443, A2 => n4435, ZN => n2735);
   U1729 : NAND2_X1 port map( A1 => n4439, A2 => n4430, ZN => n5606);
   U1730 : NAND2_X1 port map( A1 => n4439, A2 => n4430, ZN => n2736);
   U1731 : BUF_X1 port map( A => n2752, Z => n5467);
   U1732 : BUF_X1 port map( A => n2752, Z => n5468);
   U1733 : NAND3_X1 port map( A1 => n4458, A2 => n4441, A3 => n4435, ZN => 
                           n2721);
   U1734 : BUF_X1 port map( A => n4476, Z => n5501);
   U1735 : BUF_X1 port map( A => n4476, Z => n5502);
   U1736 : BUF_X1 port map( A => rst, Z => n6072);
   U1737 : NOR4_X1 port map( A1 => n5062, A2 => n5063, A3 => n5064, A4 => n5065
                           , ZN => n5061);
   U1738 : OAI221_X1 port map( B1 => n5962, B2 => n5585, C1 => net108129, C2 =>
                           n5494, A => n5066, ZN => n5065);
   U1739 : OAI221_X1 port map( B1 => n2116, B2 => n5459, C1 => n5312, C2 => 
                           n5464, A => n5077, ZN => n5064);
   U1740 : OAI221_X1 port map( B1 => n2224, B2 => n5561, C1 => n2511, C2 => 
                           n5454, A => n5082, ZN => n5063);
   U1741 : NOR4_X1 port map( A1 => n5044, A2 => n5045, A3 => n5046, A4 => n5047
                           , ZN => n5043);
   U1742 : OAI221_X1 port map( B1 => n5965, B2 => n5586, C1 => net108130, C2 =>
                           n5495, A => n5048, ZN => n5047);
   U1743 : OAI221_X1 port map( B1 => n2353, B2 => n5460, C1 => n5280, C2 => 
                           n5465, A => n5049, ZN => n5046);
   U1744 : OAI221_X1 port map( B1 => n2930, B2 => n5562, C1 => n2121, C2 => 
                           n5455, A => n5050, ZN => n5045);
   U1745 : NOR4_X1 port map( A1 => n5026, A2 => n5027, A3 => n5028, A4 => n5029
                           , ZN => n5025);
   U1746 : OAI221_X1 port map( B1 => n5968, B2 => n5584, C1 => net108131, C2 =>
                           n5496, A => n5030, ZN => n5029);
   U1747 : OAI221_X1 port map( B1 => n2354, B2 => n5458, C1 => n5281, C2 => 
                           n5463, A => n5031, ZN => n5028);
   U1748 : OAI221_X1 port map( B1 => n2931, B2 => n4485, C1 => n2122, C2 => 
                           n5453, A => n5032, ZN => n5027);
   U1749 : NOR4_X1 port map( A1 => n5008, A2 => n5009, A3 => n5010, A4 => n5011
                           , ZN => n5007);
   U1750 : OAI221_X1 port map( B1 => n5971, B2 => n5584, C1 => net108132, C2 =>
                           n5497, A => n5012, ZN => n5011);
   U1751 : OAI221_X1 port map( B1 => n2357, B2 => n5458, C1 => n5282, C2 => 
                           n5463, A => n5013, ZN => n5010);
   U1752 : OAI221_X1 port map( B1 => n2932, B2 => n5561, C1 => n2123, C2 => 
                           n5453, A => n5014, ZN => n5009);
   U1753 : NOR4_X1 port map( A1 => n4990, A2 => n4991, A3 => n4992, A4 => n4993
                           , ZN => n4989);
   U1754 : OAI221_X1 port map( B1 => n5974, B2 => n5585, C1 => net108133, C2 =>
                           n5498, A => n4994, ZN => n4993);
   U1755 : OAI221_X1 port map( B1 => n2358, B2 => n5459, C1 => n5283, C2 => 
                           n5464, A => n4995, ZN => n4992);
   U1756 : OAI221_X1 port map( B1 => n2933, B2 => n5562, C1 => n2124, C2 => 
                           n5454, A => n4996, ZN => n4991);
   U1757 : NOR4_X1 port map( A1 => n4972, A2 => n4973, A3 => n4974, A4 => n4975
                           , ZN => n4971);
   U1758 : OAI221_X1 port map( B1 => n5977, B2 => n5585, C1 => net108134, C2 =>
                           n5499, A => n4976, ZN => n4975);
   U1759 : OAI221_X1 port map( B1 => n2359, B2 => n5459, C1 => n5284, C2 => 
                           n5464, A => n4977, ZN => n4974);
   U1760 : OAI221_X1 port map( B1 => n2934, B2 => n4485, C1 => n2125, C2 => 
                           n5454, A => n4978, ZN => n4973);
   U1761 : NOR4_X1 port map( A1 => n4954, A2 => n4955, A3 => n4956, A4 => n4957
                           , ZN => n4953);
   U1762 : OAI221_X1 port map( B1 => n5980, B2 => n5586, C1 => net108135, C2 =>
                           n5500, A => n4958, ZN => n4957);
   U1763 : OAI221_X1 port map( B1 => n2360, B2 => n5460, C1 => n5285, C2 => 
                           n5465, A => n4959, ZN => n4956);
   U1764 : OAI221_X1 port map( B1 => n2935, B2 => n5561, C1 => n2126, C2 => 
                           n5455, A => n4960, ZN => n4955);
   U1765 : NOR4_X1 port map( A1 => n4936, A2 => n4937, A3 => n4938, A4 => n4939
                           , ZN => n4935);
   U1766 : OAI221_X1 port map( B1 => n5983, B2 => n5584, C1 => net108136, C2 =>
                           n5501, A => n4940, ZN => n4939);
   U1767 : OAI221_X1 port map( B1 => n2361, B2 => n5458, C1 => n5286, C2 => 
                           n5463, A => n4941, ZN => n4938);
   U1768 : OAI221_X1 port map( B1 => n2936, B2 => n5562, C1 => n2127, C2 => 
                           n5453, A => n4942, ZN => n4937);
   U1769 : NOR4_X1 port map( A1 => n4900, A2 => n4901, A3 => n4902, A4 => n4903
                           , ZN => n4899);
   U1770 : OAI221_X1 port map( B1 => n5989, B2 => n5585, C1 => net108138, C2 =>
                           n5496, A => n4904, ZN => n4903);
   U1771 : OAI221_X1 port map( B1 => n2362, B2 => n5459, C1 => n5287, C2 => 
                           n5464, A => n4905, ZN => n4902);
   U1772 : OAI221_X1 port map( B1 => n2937, B2 => n5561, C1 => n2128, C2 => 
                           n5454, A => n4906, ZN => n4901);
   U1773 : NOR4_X1 port map( A1 => n4882, A2 => n4883, A3 => n4884, A4 => n4885
                           , ZN => n4881);
   U1774 : OAI221_X1 port map( B1 => n5992, B2 => n5586, C1 => net108139, C2 =>
                           n5497, A => n4886, ZN => n4885);
   U1775 : OAI221_X1 port map( B1 => n2363, B2 => n5460, C1 => n5288, C2 => 
                           n5465, A => n4887, ZN => n4884);
   U1776 : OAI221_X1 port map( B1 => n2938, B2 => n5562, C1 => n2129, C2 => 
                           n5455, A => n4888, ZN => n4883);
   U1777 : NOR4_X1 port map( A1 => n4864, A2 => n4865, A3 => n4866, A4 => n4867
                           , ZN => n4863);
   U1778 : OAI221_X1 port map( B1 => n5995, B2 => n5584, C1 => net108140, C2 =>
                           n5494, A => n4868, ZN => n4867);
   U1779 : OAI221_X1 port map( B1 => n2364, B2 => n5458, C1 => n5289, C2 => 
                           n5463, A => n4869, ZN => n4866);
   U1780 : OAI221_X1 port map( B1 => n2939, B2 => n4485, C1 => n2130, C2 => 
                           n5453, A => n4870, ZN => n4865);
   U1781 : NOR4_X1 port map( A1 => n4846, A2 => n4847, A3 => n4848, A4 => n4849
                           , ZN => n4845);
   U1782 : OAI221_X1 port map( B1 => n5998, B2 => n5584, C1 => net108141, C2 =>
                           n5502, A => n4850, ZN => n4849);
   U1783 : OAI221_X1 port map( B1 => n2365, B2 => n5458, C1 => n5290, C2 => 
                           n5463, A => n4851, ZN => n4848);
   U1784 : OAI221_X1 port map( B1 => n2940, B2 => n5561, C1 => n2131, C2 => 
                           n5453, A => n4852, ZN => n4847);
   U1785 : NOR4_X1 port map( A1 => n4828, A2 => n4829, A3 => n4830, A4 => n4831
                           , ZN => n4827);
   U1786 : OAI221_X1 port map( B1 => n6001, B2 => n5585, C1 => net108142, C2 =>
                           n5491, A => n4832, ZN => n4831);
   U1787 : OAI221_X1 port map( B1 => n2366, B2 => n5459, C1 => n5291, C2 => 
                           n5464, A => n4833, ZN => n4830);
   U1788 : OAI221_X1 port map( B1 => n2941, B2 => n5562, C1 => n2132, C2 => 
                           n5454, A => n4834, ZN => n4829);
   U1789 : NOR4_X1 port map( A1 => n4810, A2 => n4811, A3 => n4812, A4 => n4813
                           , ZN => n4809);
   U1790 : OAI221_X1 port map( B1 => n6004, B2 => n5585, C1 => net108143, C2 =>
                           n5492, A => n4814, ZN => n4813);
   U1791 : OAI221_X1 port map( B1 => n2367, B2 => n5459, C1 => n5292, C2 => 
                           n5464, A => n4815, ZN => n4812);
   U1792 : OAI221_X1 port map( B1 => n2942, B2 => n4485, C1 => n2133, C2 => 
                           n5454, A => n4816, ZN => n4811);
   U1793 : NOR4_X1 port map( A1 => n4792, A2 => n4793, A3 => n4794, A4 => n4795
                           , ZN => n4791);
   U1794 : OAI221_X1 port map( B1 => n6007, B2 => n5586, C1 => net108144, C2 =>
                           n5493, A => n4796, ZN => n4795);
   U1795 : OAI221_X1 port map( B1 => n2368, B2 => n5460, C1 => n5293, C2 => 
                           n5465, A => n4797, ZN => n4794);
   U1796 : OAI221_X1 port map( B1 => n2943, B2 => n5561, C1 => n2134, C2 => 
                           n5455, A => n4798, ZN => n4793);
   U1797 : NOR4_X1 port map( A1 => n4774, A2 => n4775, A3 => n4776, A4 => n4777
                           , ZN => n4773);
   U1798 : OAI221_X1 port map( B1 => n6010, B2 => n5584, C1 => net108145, C2 =>
                           n5494, A => n4778, ZN => n4777);
   U1799 : OAI221_X1 port map( B1 => n2369, B2 => n5458, C1 => n5294, C2 => 
                           n5463, A => n4779, ZN => n4776);
   U1800 : OAI221_X1 port map( B1 => n2944, B2 => n5562, C1 => n2135, C2 => 
                           n5453, A => n4780, ZN => n4775);
   U1801 : NOR4_X1 port map( A1 => n4738, A2 => n4739, A3 => n4740, A4 => n4741
                           , ZN => n4737);
   U1802 : OAI221_X1 port map( B1 => n6016, B2 => n5585, C1 => net108147, C2 =>
                           n5496, A => n4742, ZN => n4741);
   U1803 : OAI221_X1 port map( B1 => n2370, B2 => n5459, C1 => n5295, C2 => 
                           n5464, A => n4743, ZN => n4740);
   U1804 : OAI221_X1 port map( B1 => n2945, B2 => n5561, C1 => n2136, C2 => 
                           n5454, A => n4744, ZN => n4739);
   U1805 : NOR4_X1 port map( A1 => n4720, A2 => n4721, A3 => n4722, A4 => n4723
                           , ZN => n4719);
   U1806 : OAI221_X1 port map( B1 => n6019, B2 => n5586, C1 => net108148, C2 =>
                           n5497, A => n4724, ZN => n4723);
   U1807 : OAI221_X1 port map( B1 => n2371, B2 => n5460, C1 => n5296, C2 => 
                           n5465, A => n4725, ZN => n4722);
   U1808 : OAI221_X1 port map( B1 => n2946, B2 => n5562, C1 => n2137, C2 => 
                           n5455, A => n4726, ZN => n4721);
   U1809 : NOR4_X1 port map( A1 => n4522, A2 => n4523, A3 => n4524, A4 => n4525
                           , ZN => n4521);
   U1810 : OAI221_X1 port map( B1 => n6052, B2 => n5584, C1 => net108159, C2 =>
                           n5492, A => n4526, ZN => n4525);
   U1811 : OAI221_X1 port map( B1 => n2372, B2 => n5458, C1 => n5297, C2 => 
                           n5463, A => n4527, ZN => n4524);
   U1812 : OAI221_X1 port map( B1 => n2947, B2 => n5561, C1 => n2138, C2 => 
                           n5453, A => n4528, ZN => n4523);
   U1813 : NOR4_X1 port map( A1 => n4471, A2 => n4472, A3 => n4473, A4 => n4474
                           , ZN => n4470);
   U1814 : OAI221_X1 port map( B1 => n6055, B2 => n5585, C1 => net108160, C2 =>
                           n5493, A => n4477, ZN => n4474);
   U1815 : OAI221_X1 port map( B1 => n2373, B2 => n5459, C1 => n5298, C2 => 
                           n5464, A => n4482, ZN => n4473);
   U1816 : OAI221_X1 port map( B1 => n2948, B2 => n5562, C1 => n2139, C2 => 
                           n5454, A => n4487, ZN => n4472);
   U1817 : NOR4_X1 port map( A1 => n4918, A2 => n4919, A3 => n4920, A4 => n4921
                           , ZN => n4917);
   U1818 : OAI221_X1 port map( B1 => n5986, B2 => n5586, C1 => net108137, C2 =>
                           n5492, A => n4922, ZN => n4921);
   U1819 : OAI221_X1 port map( B1 => n2374, B2 => n5460, C1 => n5299, C2 => 
                           n5465, A => n4923, ZN => n4920);
   U1820 : OAI221_X1 port map( B1 => n2949, B2 => n4485, C1 => n2140, C2 => 
                           n5455, A => n4924, ZN => n4919);
   U1821 : NOR4_X1 port map( A1 => n4702, A2 => n4703, A3 => n4704, A4 => n4705
                           , ZN => n4701);
   U1822 : OAI221_X1 port map( B1 => n6022, B2 => n5584, C1 => net108149, C2 =>
                           n5493, A => n4706, ZN => n4705);
   U1823 : OAI221_X1 port map( B1 => n2375, B2 => n5458, C1 => n5300, C2 => 
                           n5463, A => n4707, ZN => n4704);
   U1824 : OAI221_X1 port map( B1 => n4014, B2 => n4485, C1 => n2141, C2 => 
                           n5453, A => n4708, ZN => n4703);
   U1825 : NOR4_X1 port map( A1 => n4684, A2 => n4685, A3 => n4686, A4 => n4687
                           , ZN => n4683);
   U1826 : OAI221_X1 port map( B1 => n6025, B2 => n5584, C1 => net108150, C2 =>
                           n5498, A => n4688, ZN => n4687);
   U1827 : OAI221_X1 port map( B1 => n2376, B2 => n5458, C1 => n5301, C2 => 
                           n5463, A => n4689, ZN => n4686);
   U1828 : OAI221_X1 port map( B1 => n4033, B2 => n5561, C1 => n2142, C2 => 
                           n5453, A => n4690, ZN => n4685);
   U1829 : NOR4_X1 port map( A1 => n4666, A2 => n4667, A3 => n4668, A4 => n4669
                           , ZN => n4665);
   U1830 : OAI221_X1 port map( B1 => n6028, B2 => n5585, C1 => net108151, C2 =>
                           n5499, A => n4670, ZN => n4669);
   U1831 : OAI221_X1 port map( B1 => n2377, B2 => n5459, C1 => n5302, C2 => 
                           n5464, A => n4671, ZN => n4668);
   U1832 : OAI221_X1 port map( B1 => n4052, B2 => n5562, C1 => n2143, C2 => 
                           n5454, A => n4672, ZN => n4667);
   U1833 : NOR4_X1 port map( A1 => n4648, A2 => n4649, A3 => n4650, A4 => n4651
                           , ZN => n4647);
   U1834 : OAI221_X1 port map( B1 => n6031, B2 => n5585, C1 => net108152, C2 =>
                           n5495, A => n4652, ZN => n4651);
   U1835 : OAI221_X1 port map( B1 => n2378, B2 => n5459, C1 => n5303, C2 => 
                           n5464, A => n4653, ZN => n4650);
   U1836 : OAI221_X1 port map( B1 => n4071, B2 => n4485, C1 => n2144, C2 => 
                           n5454, A => n4654, ZN => n4649);
   U1837 : NOR4_X1 port map( A1 => n4630, A2 => n4631, A3 => n4632, A4 => n4633
                           , ZN => n4629);
   U1838 : OAI221_X1 port map( B1 => n6034, B2 => n5586, C1 => net108153, C2 =>
                           n5498, A => n4634, ZN => n4633);
   U1839 : OAI221_X1 port map( B1 => n2379, B2 => n5460, C1 => n5304, C2 => 
                           n5465, A => n4635, ZN => n4632);
   U1840 : OAI221_X1 port map( B1 => n4090, B2 => n5561, C1 => n2145, C2 => 
                           n5455, A => n4636, ZN => n4631);
   U1841 : NOR4_X1 port map( A1 => n4612, A2 => n4613, A3 => n4614, A4 => n4615
                           , ZN => n4611);
   U1842 : OAI221_X1 port map( B1 => n6037, B2 => n5584, C1 => net108154, C2 =>
                           n5499, A => n4616, ZN => n4615);
   U1843 : OAI221_X1 port map( B1 => n2380, B2 => n5458, C1 => n5305, C2 => 
                           n5463, A => n4617, ZN => n4614);
   U1844 : OAI221_X1 port map( B1 => n4109, B2 => n5562, C1 => n2146, C2 => 
                           n5453, A => n4618, ZN => n4613);
   U1845 : NOR4_X1 port map( A1 => n4576, A2 => n4577, A3 => n4578, A4 => n4579
                           , ZN => n4575);
   U1846 : OAI221_X1 port map( B1 => n6043, B2 => n5585, C1 => net108156, C2 =>
                           n5501, A => n4580, ZN => n4579);
   U1847 : OAI221_X1 port map( B1 => n2381, B2 => n5459, C1 => n5306, C2 => 
                           n5464, A => n4581, ZN => n4578);
   U1848 : OAI221_X1 port map( B1 => n4128, B2 => n5561, C1 => n2148, C2 => 
                           n5454, A => n4582, ZN => n4577);
   U1849 : NOR4_X1 port map( A1 => n4558, A2 => n4559, A3 => n4560, A4 => n4561
                           , ZN => n4557);
   U1850 : OAI221_X1 port map( B1 => n6046, B2 => n5586, C1 => net108157, C2 =>
                           n5502, A => n4562, ZN => n4561);
   U1851 : OAI221_X1 port map( B1 => n2382, B2 => n5460, C1 => n5307, C2 => 
                           n5465, A => n4563, ZN => n4560);
   U1852 : OAI221_X1 port map( B1 => n4147, B2 => n5562, C1 => n2149, C2 => 
                           n5455, A => n4564, ZN => n4559);
   U1853 : NOR4_X1 port map( A1 => n4756, A2 => n4757, A3 => n4758, A4 => n4759
                           , ZN => n4755);
   U1854 : OAI221_X1 port map( B1 => n6013, B2 => n5586, C1 => net108146, C2 =>
                           n5495, A => n4760, ZN => n4759);
   U1855 : OAI221_X1 port map( B1 => n2383, B2 => n5460, C1 => n5308, C2 => 
                           n5465, A => n4761, ZN => n4758);
   U1856 : OAI221_X1 port map( B1 => n4166, B2 => n4485, C1 => n2150, C2 => 
                           n5455, A => n4762, ZN => n4757);
   U1857 : NOR4_X1 port map( A1 => n4594, A2 => n4595, A3 => n4596, A4 => n4597
                           , ZN => n4593);
   U1858 : OAI221_X1 port map( B1 => n6040, B2 => n5586, C1 => net108155, C2 =>
                           n5500, A => n4598, ZN => n4597);
   U1859 : OAI221_X1 port map( B1 => n2384, B2 => n5460, C1 => n5309, C2 => 
                           n5465, A => n4599, ZN => n4596);
   U1860 : OAI221_X1 port map( B1 => n4185, B2 => n4485, C1 => n2151, C2 => 
                           n5455, A => n4600, ZN => n4595);
   U1861 : NOR4_X1 port map( A1 => n4540, A2 => n4541, A3 => n4542, A4 => n4543
                           , ZN => n4539);
   U1862 : OAI221_X1 port map( B1 => n6049, B2 => n5584, C1 => net108158, C2 =>
                           n5491, A => n4544, ZN => n4543);
   U1863 : OAI221_X1 port map( B1 => n2385, B2 => n5458, C1 => n5310, C2 => 
                           n5463, A => n4545, ZN => n4542);
   U1864 : OAI221_X1 port map( B1 => n4204, B2 => n4485, C1 => n2152, C2 => 
                           n5453, A => n4546, ZN => n4541);
   U1865 : NOR3_X1 port map( A1 => n2181, A2 => wr_addr(4), A3 => n2182, ZN => 
                           n1768);
   U1866 : INV_X1 port map( A => en, ZN => n2181);
   U1867 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_1_port, C1 => 
                           n5679, C2 => registers_9_1_port, A => n4400, ZN => 
                           n4399);
   U1868 : OAI222_X1 port map( A1 => n5184, A2 => n5687, B1 => n4401, B2 => 
                           n5593, C1 => n2423, C2 => n5684, ZN => n4400);
   U1869 : NOR4_X1 port map( A1 => n4402, A2 => n4403, A3 => n4404, A4 => n4405
                           , ZN => n4401);
   U1870 : OAI221_X1 port map( B1 => n5124, B2 => n5600, C1 => n2228, C2 => 
                           n5608, A => n4409, ZN => n4402);
   U1871 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_3_port, C1 => 
                           n2710, C2 => registers_9_3_port, A => n4362, ZN => 
                           n4361);
   U1872 : OAI222_X1 port map( A1 => n5185, A2 => n5686, B1 => n4363, B2 => 
                           n2714, C1 => n2425, C2 => n5683, ZN => n4362);
   U1873 : NOR4_X1 port map( A1 => n4364, A2 => n4365, A3 => n4366, A4 => n4367
                           , ZN => n4363);
   U1874 : OAI221_X1 port map( B1 => n5125, B2 => n5599, C1 => n2229, C2 => 
                           n5608, A => n4371, ZN => n4364);
   U1875 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_4_port, C1 => 
                           n5679, C2 => registers_9_4_port, A => n4343, ZN => 
                           n4342);
   U1876 : OAI222_X1 port map( A1 => n5186, A2 => n5687, B1 => n4344, B2 => 
                           n5593, C1 => n2426, C2 => n5685, ZN => n4343);
   U1877 : NOR4_X1 port map( A1 => n4345, A2 => n4346, A3 => n4347, A4 => n4348
                           , ZN => n4344);
   U1878 : OAI221_X1 port map( B1 => n5126, B2 => n5600, C1 => n2230, C2 => 
                           n5609, A => n4352, ZN => n4345);
   U1879 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_6_port, C1 => 
                           n2710, C2 => registers_9_6_port, A => n4305, ZN => 
                           n4304);
   U1880 : OAI222_X1 port map( A1 => n5187, A2 => n5686, B1 => n4306, B2 => 
                           n2714, C1 => n2427, C2 => n5684, ZN => n4305);
   U1881 : NOR4_X1 port map( A1 => n4307, A2 => n4308, A3 => n4309, A4 => n4310
                           , ZN => n4306);
   U1882 : OAI221_X1 port map( B1 => n5127, B2 => n5602, C1 => n2231, C2 => 
                           n5609, A => n4314, ZN => n4307);
   U1883 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_7_port, C1 => 
                           n5679, C2 => registers_9_7_port, A => n4286, ZN => 
                           n4285);
   U1884 : OAI222_X1 port map( A1 => n5188, A2 => n5687, B1 => n4287, B2 => 
                           n5593, C1 => n2428, C2 => n5683, ZN => n4286);
   U1885 : NOR4_X1 port map( A1 => n4288, A2 => n4289, A3 => n4290, A4 => n4291
                           , ZN => n4287);
   U1886 : OAI221_X1 port map( B1 => n5128, B2 => n5601, C1 => n2232, C2 => 
                           n5610, A => n4295, ZN => n4288);
   U1887 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_9_port, C1 => 
                           n2710, C2 => registers_9_9_port, A => n4248, ZN => 
                           n4247);
   U1888 : OAI222_X1 port map( A1 => n5189, A2 => n5686, B1 => n4249, B2 => 
                           n2714, C1 => n2429, C2 => n5685, ZN => n4248);
   U1889 : NOR4_X1 port map( A1 => n4250, A2 => n4251, A3 => n4252, A4 => n4253
                           , ZN => n4249);
   U1890 : OAI221_X1 port map( B1 => n5129, B2 => n5604, C1 => n2233, C2 => 
                           n5612, A => n4257, ZN => n4250);
   U1891 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_10_port, C1 => 
                           n5679, C2 => registers_9_10_port, A => n4229, ZN => 
                           n4228);
   U1892 : OAI222_X1 port map( A1 => n5190, A2 => n5687, B1 => n4230, B2 => 
                           n5593, C1 => n2430, C2 => n5684, ZN => n4229);
   U1893 : NOR4_X1 port map( A1 => n4231, A2 => n4232, A3 => n4233, A4 => n4234
                           , ZN => n4230);
   U1894 : OAI221_X1 port map( B1 => n5130, B2 => n5603, C1 => n2234, C2 => 
                           n5607, A => n4238, ZN => n4231);
   U1895 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_12_port, C1 => 
                           n2710, C2 => registers_9_12_port, A => n4191, ZN => 
                           n4190);
   U1896 : OAI222_X1 port map( A1 => n5191, A2 => n5686, B1 => n4192, B2 => 
                           n2714, C1 => n2431, C2 => n5683, ZN => n4191);
   U1897 : NOR4_X1 port map( A1 => n4193, A2 => n4194, A3 => n4195, A4 => n4196
                           , ZN => n4192);
   U1898 : OAI221_X1 port map( B1 => n5131, B2 => n5600, C1 => n2235, C2 => 
                           n5611, A => n4200, ZN => n4193);
   U1899 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_13_port, C1 => 
                           n5679, C2 => registers_9_13_port, A => n4172, ZN => 
                           n4171);
   U1900 : OAI222_X1 port map( A1 => n5192, A2 => n5687, B1 => n4173, B2 => 
                           n5593, C1 => n2432, C2 => n5685, ZN => n4172);
   U1901 : NOR4_X1 port map( A1 => n4174, A2 => n4175, A3 => n4176, A4 => n4177
                           , ZN => n4173);
   U1902 : OAI221_X1 port map( B1 => n5132, B2 => n5602, C1 => n2236, C2 => 
                           n5612, A => n4181, ZN => n4174);
   U1903 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_15_port, C1 => 
                           n2710, C2 => registers_9_15_port, A => n4134, ZN => 
                           n4133);
   U1904 : OAI222_X1 port map( A1 => n5193, A2 => n5686, B1 => n4135, B2 => 
                           n2714, C1 => n2433, C2 => n5684, ZN => n4134);
   U1905 : NOR4_X1 port map( A1 => n4136, A2 => n4137, A3 => n4138, A4 => n4139
                           , ZN => n4135);
   U1906 : OAI221_X1 port map( B1 => n5133, B2 => n5601, C1 => n2237, C2 => 
                           n5610, A => n4143, ZN => n4136);
   U1907 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_16_port, C1 => 
                           n5679, C2 => registers_9_16_port, A => n4115, ZN => 
                           n4114);
   U1908 : OAI222_X1 port map( A1 => n5194, A2 => n5687, B1 => n4116, B2 => 
                           n5593, C1 => n2434, C2 => n5683, ZN => n4115);
   U1909 : NOR4_X1 port map( A1 => n4117, A2 => n4118, A3 => n4119, A4 => n4120
                           , ZN => n4116);
   U1910 : OAI221_X1 port map( B1 => n5134, B2 => n5602, C1 => n2238, C2 => 
                           n5611, A => n4124, ZN => n4117);
   U1911 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_18_port, C1 => 
                           n2710, C2 => registers_9_18_port, A => n4077, ZN => 
                           n4076);
   U1912 : OAI222_X1 port map( A1 => n5195, A2 => n5686, B1 => n4078, B2 => 
                           n2714, C1 => n2435, C2 => n5685, ZN => n4077);
   U1913 : NOR4_X1 port map( A1 => n4079, A2 => n4080, A3 => n4081, A4 => n4082
                           , ZN => n4078);
   U1914 : OAI221_X1 port map( B1 => n5135, B2 => n5603, C1 => n2239, C2 => 
                           n5607, A => n4086, ZN => n4079);
   U1915 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_19_port, C1 => 
                           n5679, C2 => registers_9_19_port, A => n4058, ZN => 
                           n4057);
   U1916 : OAI222_X1 port map( A1 => n5196, A2 => n5687, B1 => n4059, B2 => 
                           n5593, C1 => n2436, C2 => n5684, ZN => n4058);
   U1917 : NOR4_X1 port map( A1 => n4060, A2 => n4061, A3 => n4062, A4 => n4063
                           , ZN => n4059);
   U1918 : OAI221_X1 port map( B1 => n5136, B2 => n5604, C1 => n2240, C2 => 
                           n5608, A => n4067, ZN => n4060);
   U1919 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_21_port, C1 => 
                           n2710, C2 => registers_9_21_port, A => n4020, ZN => 
                           n4019);
   U1920 : OAI222_X1 port map( A1 => n5197, A2 => n5686, B1 => n4021, B2 => 
                           n2714, C1 => n2437, C2 => n5683, ZN => n4020);
   U1921 : NOR4_X1 port map( A1 => n4022, A2 => n4023, A3 => n4024, A4 => n4025
                           , ZN => n4021);
   U1922 : OAI221_X1 port map( B1 => n5137, B2 => n5604, C1 => n2241, C2 => 
                           n5608, A => n4029, ZN => n4022);
   U1923 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_22_port, C1 => 
                           n5679, C2 => registers_9_22_port, A => n2914, ZN => 
                           n2913);
   U1924 : OAI222_X1 port map( A1 => n5198, A2 => n5687, B1 => n2915, B2 => 
                           n5593, C1 => n2438, C2 => n5685, ZN => n2914);
   U1925 : NOR4_X1 port map( A1 => n2916, A2 => n2917, A3 => n2918, A4 => n2950
                           , ZN => n2915);
   U1926 : OAI221_X1 port map( B1 => n5138, B2 => n5604, C1 => n2242, C2 => 
                           n5609, A => n4010, ZN => n2916);
   U1927 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_24_port, C1 => 
                           n2710, C2 => registers_9_24_port, A => n2876, ZN => 
                           n2875);
   U1928 : OAI222_X1 port map( A1 => n5199, A2 => n5686, B1 => n2877, B2 => 
                           n2714, C1 => n2439, C2 => n5684, ZN => n2876);
   U1929 : NOR4_X1 port map( A1 => n2878, A2 => n2879, A3 => n2880, A4 => n2881
                           , ZN => n2877);
   U1930 : OAI221_X1 port map( B1 => n5139, B2 => n5601, C1 => n2243, C2 => 
                           n5609, A => n2885, ZN => n2878);
   U1931 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_25_port, C1 => 
                           n5679, C2 => registers_9_25_port, A => n2857, ZN => 
                           n2856);
   U1932 : OAI222_X1 port map( A1 => n5200, A2 => n5687, B1 => n2858, B2 => 
                           n5593, C1 => n2440, C2 => n5683, ZN => n2857);
   U1933 : NOR4_X1 port map( A1 => n2859, A2 => n2860, A3 => n2861, A4 => n2862
                           , ZN => n2858);
   U1934 : OAI221_X1 port map( B1 => n5140, B2 => n5605, C1 => n2244, C2 => 
                           n5610, A => n2866, ZN => n2859);
   U1935 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_27_port, C1 => 
                           n2710, C2 => registers_9_27_port, A => n2819, ZN => 
                           n2818);
   U1936 : OAI222_X1 port map( A1 => n5201, A2 => n5686, B1 => n2820, B2 => 
                           n2714, C1 => n2441, C2 => n5685, ZN => n2819);
   U1937 : NOR4_X1 port map( A1 => n2821, A2 => n2822, A3 => n2823, A4 => n2824
                           , ZN => n2820);
   U1938 : OAI221_X1 port map( B1 => n5141, B2 => n5605, C1 => n2117, C2 => 
                           n5612, A => n2828, ZN => n2821);
   U1939 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_28_port, C1 => 
                           n5679, C2 => registers_9_28_port, A => n2800, ZN => 
                           n2799);
   U1940 : OAI222_X1 port map( A1 => n5202, A2 => n5687, B1 => n2801, B2 => 
                           n5593, C1 => n2442, C2 => n5684, ZN => n2800);
   U1941 : NOR4_X1 port map( A1 => n2802, A2 => n2803, A3 => n2804, A4 => n2805
                           , ZN => n2801);
   U1942 : OAI221_X1 port map( B1 => n5142, B2 => n5600, C1 => n2245, C2 => 
                           n5607, A => n2809, ZN => n2802);
   U1943 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_30_port, C1 => 
                           n2710, C2 => registers_9_30_port, A => n2762, ZN => 
                           n2761);
   U1944 : OAI222_X1 port map( A1 => n5203, A2 => n5686, B1 => n2763, B2 => 
                           n2714, C1 => n2443, C2 => n5683, ZN => n2762);
   U1945 : NOR4_X1 port map( A1 => n2764, A2 => n2765, A3 => n2766, A4 => n2767
                           , ZN => n2763);
   U1946 : OAI221_X1 port map( B1 => n5143, B2 => n5599, C1 => n2246, C2 => 
                           n5611, A => n2771, ZN => n2764);
   U1947 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_31_port, C1 => 
                           n5679, C2 => registers_9_31_port, A => n2711, ZN => 
                           n2708);
   U1948 : OAI222_X1 port map( A1 => n5204, A2 => n5687, B1 => n2713, B2 => 
                           n5593, C1 => n2444, C2 => n5685, ZN => n2711);
   U1949 : NOR4_X1 port map( A1 => n2716, A2 => n2717, A3 => n2718, A4 => n2719
                           , ZN => n2713);
   U1950 : OAI221_X1 port map( B1 => n5144, B2 => n5599, C1 => n2247, C2 => 
                           n5612, A => n2737, ZN => n2716);
   U1951 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_2_port, C1 => 
                           n5680, C2 => registers_9_2_port, A => n4381, ZN => 
                           n4380);
   U1952 : OAI222_X1 port map( A1 => n5205, A2 => n2712, B1 => n4382, B2 => 
                           n5594, C1 => n2445, C2 => n5683, ZN => n4381);
   U1953 : NOR4_X1 port map( A1 => n4383, A2 => n4384, A3 => n4385, A4 => n4386
                           , ZN => n4382);
   U1954 : OAI221_X1 port map( B1 => n5145, B2 => n5600, C1 => n2248, C2 => 
                           n5607, A => n4390, ZN => n4383);
   U1955 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_5_port, C1 => 
                           n5680, C2 => registers_9_5_port, A => n4324, ZN => 
                           n4323);
   U1956 : OAI222_X1 port map( A1 => n5206, A2 => n2712, B1 => n4325, B2 => 
                           n5594, C1 => n2446, C2 => n5684, ZN => n4324);
   U1957 : NOR4_X1 port map( A1 => n4326, A2 => n4327, A3 => n4328, A4 => n4329
                           , ZN => n4325);
   U1958 : OAI221_X1 port map( B1 => n5146, B2 => n5601, C1 => n2249, C2 => 
                           n5610, A => n4333, ZN => n4326);
   U1959 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_8_port, C1 => 
                           n5680, C2 => registers_9_8_port, A => n4267, ZN => 
                           n4266);
   U1960 : OAI222_X1 port map( A1 => n5207, A2 => n2712, B1 => n4268, B2 => 
                           n5594, C1 => n2447, C2 => n5685, ZN => n4267);
   U1961 : NOR4_X1 port map( A1 => n4269, A2 => n4270, A3 => n4271, A4 => n4272
                           , ZN => n4268);
   U1962 : OAI221_X1 port map( B1 => n5147, B2 => n5602, C1 => n2250, C2 => 
                           n5611, A => n4276, ZN => n4269);
   U1963 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_11_port, C1 => 
                           n5680, C2 => registers_9_11_port, A => n4210, ZN => 
                           n4209);
   U1964 : OAI222_X1 port map( A1 => n5208, A2 => n2712, B1 => n4211, B2 => 
                           n5594, C1 => n2448, C2 => n5683, ZN => n4210);
   U1965 : NOR4_X1 port map( A1 => n4212, A2 => n4213, A3 => n4214, A4 => n4215
                           , ZN => n4211);
   U1966 : OAI221_X1 port map( B1 => n5148, B2 => n5603, C1 => n2251, C2 => 
                           n5608, A => n4219, ZN => n4212);
   U1967 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_14_port, C1 => 
                           n5680, C2 => registers_9_14_port, A => n4153, ZN => 
                           n4152);
   U1968 : OAI222_X1 port map( A1 => n5209, A2 => n2712, B1 => n4154, B2 => 
                           n5594, C1 => n2449, C2 => n5684, ZN => n4153);
   U1969 : NOR4_X1 port map( A1 => n4155, A2 => n4156, A3 => n4157, A4 => n4158
                           , ZN => n4154);
   U1970 : OAI221_X1 port map( B1 => n5149, B2 => n5601, C1 => n2253, C2 => 
                           n5609, A => n4162, ZN => n4155);
   U1971 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_17_port, C1 => 
                           n5680, C2 => registers_9_17_port, A => n4096, ZN => 
                           n4095);
   U1972 : OAI222_X1 port map( A1 => n5210, A2 => n2712, B1 => n4097, B2 => 
                           n5594, C1 => n2450, C2 => n5685, ZN => n4096);
   U1973 : NOR4_X1 port map( A1 => n4098, A2 => n4099, A3 => n4100, A4 => n4101
                           , ZN => n4097);
   U1974 : OAI221_X1 port map( B1 => n5150, B2 => n5603, C1 => n2254, C2 => 
                           n5612, A => n4105, ZN => n4098);
   U1975 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_20_port, C1 => 
                           n5680, C2 => registers_9_20_port, A => n4039, ZN => 
                           n4038);
   U1976 : OAI222_X1 port map( A1 => n5211, A2 => n2712, B1 => n4040, B2 => 
                           n5594, C1 => n2451, C2 => n5683, ZN => n4039);
   U1977 : NOR4_X1 port map( A1 => n4041, A2 => n4042, A3 => n4043, A4 => n4044
                           , ZN => n4040);
   U1978 : OAI221_X1 port map( B1 => n5151, B2 => n5605, C1 => n2255, C2 => 
                           n5607, A => n4048, ZN => n4041);
   U1979 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_23_port, C1 => 
                           n5680, C2 => registers_9_23_port, A => n2895, ZN => 
                           n2894);
   U1980 : OAI222_X1 port map( A1 => n5212, A2 => n2712, B1 => n2896, B2 => 
                           n5594, C1 => n2452, C2 => n5684, ZN => n2895);
   U1981 : NOR4_X1 port map( A1 => n2897, A2 => n2898, A3 => n2899, A4 => n2900
                           , ZN => n2896);
   U1982 : OAI221_X1 port map( B1 => n5152, B2 => n5602, C1 => n2256, C2 => 
                           n5610, A => n2904, ZN => n2897);
   U1983 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_26_port, C1 => 
                           n5680, C2 => registers_9_26_port, A => n2838, ZN => 
                           n2837);
   U1984 : OAI222_X1 port map( A1 => n5213, A2 => n2712, B1 => n2839, B2 => 
                           n5594, C1 => n2453, C2 => n5685, ZN => n2838);
   U1985 : NOR4_X1 port map( A1 => n2840, A2 => n2841, A3 => n2842, A4 => n2843
                           , ZN => n2839);
   U1986 : OAI221_X1 port map( B1 => n2386, B2 => n5605, C1 => n2118, C2 => 
                           n5611, A => n2847, ZN => n2840);
   U1987 : AOI221_X1 port map( B1 => n2709, B2 => registers_13_29_port, C1 => 
                           n5680, C2 => registers_9_29_port, A => n2781, ZN => 
                           n2780);
   U1988 : OAI222_X1 port map( A1 => n5214, A2 => n2712, B1 => n2782, B2 => 
                           n5594, C1 => n2454, C2 => n5683, ZN => n2781);
   U1989 : NOR4_X1 port map( A1 => n2783, A2 => n2784, A3 => n2785, A4 => n2786
                           , ZN => n2782);
   U1990 : OAI221_X1 port map( B1 => n5153, B2 => n5605, C1 => n2257, C2 => 
                           n5608, A => n2790, ZN => n2783);
   U1991 : AOI221_X1 port map( B1 => n5664, B2 => registers_30_0_port, C1 => 
                           n4436, C2 => registers_15_0_port, A => n4437, ZN => 
                           n4420);
   U1992 : INV_X1 port map( A => n5479, ZN => n4436);
   U1993 : OAI222_X1 port map( A1 => n5279, A2 => n5482, B1 => n2422, B2 => 
                           n5666, C1 => n2116, C2 => n4414, ZN => n4437);
   U1994 : AOI22_X1 port map( A1 => en, A2 => link_en, B1 => n1765, B2 => n2629
                           , ZN => n4418);
   U1995 : AND3_X1 port map( A1 => rd1_addr(2), A2 => n5090, A3 => n5506, ZN =>
                           n5080);
   U1996 : NAND4_X1 port map( A1 => n5069, A2 => n5503, A3 => rd1_addr(2), A4 
                           => n5090, ZN => n4512);
   U1997 : NAND4_X1 port map( A1 => n5079, A2 => n5505, A3 => rd1_addr(2), A4 
                           => n5090, ZN => n4502);
   U1998 : NOR2_X1 port map( A1 => n4418, A2 => link_en, ZN => n2704);
   U1999 : XNOR2_X1 port map( A => wr_addr(4), B => n4459, ZN => n4450);
   U2000 : XNOR2_X1 port map( A => wr_addr(4), B => n5096, ZN => n5074);
   U2001 : XNOR2_X1 port map( A => n4441, B => wr_addr(2), ZN => n4451);
   U2002 : XNOR2_X1 port map( A => n5095, B => wr_addr(2), ZN => n5075);
   U2003 : XNOR2_X1 port map( A => wr_addr(0), B => rd1_addr(0), ZN => n5071);
   U2004 : XNOR2_X1 port map( A => wr_addr(0), B => rd2_addr(0), ZN => n4446);
   U2005 : XNOR2_X1 port map( A => wr_addr(1), B => rd1_addr(1), ZN => n5072);
   U2006 : XNOR2_X1 port map( A => wr_addr(1), B => rd2_addr(1), ZN => n4447);
   U2007 : XNOR2_X1 port map( A => rd2_addr(3), B => n1767, ZN => n4452);
   U2008 : XNOR2_X1 port map( A => rd1_addr(3), B => n1767, ZN => n5076);
   U2009 : INV_X1 port map( A => n2180, ZN => n3527);
   U2010 : AOI22_X1 port map( A1 => d_in(0), A2 => n5390, B1 => n5836, B2 => 
                           registers_15_0_port, ZN => n2180);
   U2011 : INV_X1 port map( A => n1838, ZN => n3847);
   U2012 : AOI22_X1 port map( A1 => d_in(0), A2 => n5420, B1 => n5926, B2 => 
                           registers_5_0_port, ZN => n1838);
   U2013 : INV_X1 port map( A => n2089, ZN => n3614);
   U2014 : AOI22_X1 port map( A1 => d_in(23), A2 => n5396, B1 => n5860, B2 => 
                           registers_13_23_port, ZN => n2089);
   U2015 : AOI22_X1 port map( A1 => n5565, A2 => registers_5_0_port, B1 => 
                           n5577, B2 => registers_8_0_port, ZN => n5082);
   U2016 : AOI22_X1 port map( A1 => n5579, A2 => registers_21_0_port, B1 => 
                           n5582, B2 => registers_26_0_port, ZN => n5077);
   U2017 : AOI22_X1 port map( A1 => n5588, A2 => registers_15_0_port, B1 => 
                           n5591, B2 => registers_31_0_port, ZN => n5066);
   U2018 : AOI22_X1 port map( A1 => n5566, A2 => registers_5_1_port, B1 => 
                           n5578, B2 => registers_8_1_port, ZN => n5050);
   U2019 : AOI22_X1 port map( A1 => n5580, A2 => registers_21_1_port, B1 => 
                           n5583, B2 => registers_26_1_port, ZN => n5049);
   U2020 : AOI22_X1 port map( A1 => n5589, A2 => registers_15_1_port, B1 => 
                           n5592, B2 => registers_31_1_port, ZN => n5048);
   U2021 : AOI22_X1 port map( A1 => n5567, A2 => registers_5_2_port, B1 => 
                           n4489, B2 => registers_8_2_port, ZN => n5032);
   U2022 : AOI22_X1 port map( A1 => n4483, A2 => registers_21_2_port, B1 => 
                           n5581, B2 => registers_26_2_port, ZN => n5031);
   U2023 : AOI22_X1 port map( A1 => n5587, A2 => registers_15_2_port, B1 => 
                           n5590, B2 => registers_31_2_port, ZN => n5030);
   U2024 : AOI22_X1 port map( A1 => n5568, A2 => registers_5_3_port, B1 => 
                           n5577, B2 => registers_8_3_port, ZN => n5014);
   U2025 : AOI22_X1 port map( A1 => n5579, A2 => registers_21_3_port, B1 => 
                           n5581, B2 => registers_26_3_port, ZN => n5013);
   U2026 : AOI22_X1 port map( A1 => n5587, A2 => registers_15_3_port, B1 => 
                           n5590, B2 => registers_31_3_port, ZN => n5012);
   U2027 : AOI22_X1 port map( A1 => n5569, A2 => registers_5_4_port, B1 => 
                           n5578, B2 => registers_8_4_port, ZN => n4996);
   U2028 : AOI22_X1 port map( A1 => n5580, A2 => registers_21_4_port, B1 => 
                           n5582, B2 => registers_26_4_port, ZN => n4995);
   U2029 : AOI22_X1 port map( A1 => n5588, A2 => registers_15_4_port, B1 => 
                           n5591, B2 => registers_31_4_port, ZN => n4994);
   U2030 : AOI22_X1 port map( A1 => n5570, A2 => registers_5_5_port, B1 => 
                           n4489, B2 => registers_8_5_port, ZN => n4978);
   U2031 : AOI22_X1 port map( A1 => n4483, A2 => registers_21_5_port, B1 => 
                           n5582, B2 => registers_26_5_port, ZN => n4977);
   U2032 : AOI22_X1 port map( A1 => n5588, A2 => registers_15_5_port, B1 => 
                           n5591, B2 => registers_31_5_port, ZN => n4976);
   U2033 : AOI22_X1 port map( A1 => n5571, A2 => registers_5_6_port, B1 => 
                           n5577, B2 => registers_8_6_port, ZN => n4960);
   U2034 : AOI22_X1 port map( A1 => n5579, A2 => registers_21_6_port, B1 => 
                           n5583, B2 => registers_26_6_port, ZN => n4959);
   U2035 : AOI22_X1 port map( A1 => n5589, A2 => registers_15_6_port, B1 => 
                           n5592, B2 => registers_31_6_port, ZN => n4958);
   U2036 : AOI22_X1 port map( A1 => n5572, A2 => registers_5_7_port, B1 => 
                           n5578, B2 => registers_8_7_port, ZN => n4942);
   U2037 : AOI22_X1 port map( A1 => n5580, A2 => registers_21_7_port, B1 => 
                           n5581, B2 => registers_26_7_port, ZN => n4941);
   U2038 : AOI22_X1 port map( A1 => n5587, A2 => registers_15_7_port, B1 => 
                           n5590, B2 => registers_31_7_port, ZN => n4940);
   U2039 : AOI22_X1 port map( A1 => n5565, A2 => registers_5_8_port, B1 => 
                           n4489, B2 => registers_8_8_port, ZN => n4924);
   U2040 : AOI22_X1 port map( A1 => n4483, A2 => registers_21_8_port, B1 => 
                           n5583, B2 => registers_26_8_port, ZN => n4923);
   U2041 : AOI22_X1 port map( A1 => n5589, A2 => registers_15_8_port, B1 => 
                           n5592, B2 => registers_31_8_port, ZN => n4922);
   U2042 : AOI22_X1 port map( A1 => n5566, A2 => registers_5_9_port, B1 => 
                           n5577, B2 => registers_8_9_port, ZN => n4906);
   U2043 : AOI22_X1 port map( A1 => n5579, A2 => registers_21_9_port, B1 => 
                           n5582, B2 => registers_26_9_port, ZN => n4905);
   U2044 : AOI22_X1 port map( A1 => n5588, A2 => registers_15_9_port, B1 => 
                           n5591, B2 => registers_31_9_port, ZN => n4904);
   U2045 : AOI22_X1 port map( A1 => n5567, A2 => registers_5_10_port, B1 => 
                           n5578, B2 => registers_8_10_port, ZN => n4888);
   U2046 : AOI22_X1 port map( A1 => n5580, A2 => registers_21_10_port, B1 => 
                           n5583, B2 => registers_26_10_port, ZN => n4887);
   U2047 : AOI22_X1 port map( A1 => n5589, A2 => registers_15_10_port, B1 => 
                           n5592, B2 => registers_31_10_port, ZN => n4886);
   U2048 : AOI22_X1 port map( A1 => n5568, A2 => registers_5_11_port, B1 => 
                           n4489, B2 => registers_8_11_port, ZN => n4870);
   U2049 : AOI22_X1 port map( A1 => n4483, A2 => registers_21_11_port, B1 => 
                           n5581, B2 => registers_26_11_port, ZN => n4869);
   U2050 : AOI22_X1 port map( A1 => n5587, A2 => registers_15_11_port, B1 => 
                           n5590, B2 => registers_31_11_port, ZN => n4868);
   U2051 : AOI22_X1 port map( A1 => n5573, A2 => registers_5_12_port, B1 => 
                           n5577, B2 => registers_8_12_port, ZN => n4852);
   U2052 : AOI22_X1 port map( A1 => n5579, A2 => registers_21_12_port, B1 => 
                           n5581, B2 => registers_26_12_port, ZN => n4851);
   U2053 : AOI22_X1 port map( A1 => n5587, A2 => registers_15_12_port, B1 => 
                           n5590, B2 => registers_31_12_port, ZN => n4850);
   U2054 : AOI22_X1 port map( A1 => n5574, A2 => registers_5_13_port, B1 => 
                           n5578, B2 => registers_8_13_port, ZN => n4834);
   U2055 : AOI22_X1 port map( A1 => n5580, A2 => registers_21_13_port, B1 => 
                           n5582, B2 => registers_26_13_port, ZN => n4833);
   U2056 : AOI22_X1 port map( A1 => n5588, A2 => registers_15_13_port, B1 => 
                           n5591, B2 => registers_31_13_port, ZN => n4832);
   U2057 : AOI22_X1 port map( A1 => n5575, A2 => registers_5_14_port, B1 => 
                           n4489, B2 => registers_8_14_port, ZN => n4816);
   U2058 : AOI22_X1 port map( A1 => n4483, A2 => registers_21_14_port, B1 => 
                           n5582, B2 => registers_26_14_port, ZN => n4815);
   U2059 : AOI22_X1 port map( A1 => n5588, A2 => registers_15_14_port, B1 => 
                           n5591, B2 => registers_31_14_port, ZN => n4814);
   U2060 : AOI22_X1 port map( A1 => n5576, A2 => registers_5_15_port, B1 => 
                           n5577, B2 => registers_8_15_port, ZN => n4798);
   U2061 : AOI22_X1 port map( A1 => n5579, A2 => registers_21_15_port, B1 => 
                           n5583, B2 => registers_26_15_port, ZN => n4797);
   U2062 : AOI22_X1 port map( A1 => n5589, A2 => registers_15_15_port, B1 => 
                           n5592, B2 => registers_31_15_port, ZN => n4796);
   U2063 : AOI22_X1 port map( A1 => n5565, A2 => registers_5_16_port, B1 => 
                           n5578, B2 => registers_8_16_port, ZN => n4780);
   U2065 : AOI22_X1 port map( A1 => n5580, A2 => registers_21_16_port, B1 => 
                           n5581, B2 => registers_26_16_port, ZN => n4779);
   U2066 : AOI22_X1 port map( A1 => n5587, A2 => registers_15_16_port, B1 => 
                           n5590, B2 => registers_31_16_port, ZN => n4778);
   U2067 : AOI22_X1 port map( A1 => n5566, A2 => registers_5_17_port, B1 => 
                           n4489, B2 => registers_8_17_port, ZN => n4762);
   U2068 : AOI22_X1 port map( A1 => n4483, A2 => registers_21_17_port, B1 => 
                           n5583, B2 => registers_26_17_port, ZN => n4761);
   U2069 : AOI22_X1 port map( A1 => n5589, A2 => registers_15_17_port, B1 => 
                           n5592, B2 => registers_31_17_port, ZN => n4760);
   U2071 : AOI22_X1 port map( A1 => n5567, A2 => registers_5_18_port, B1 => 
                           n5577, B2 => registers_8_18_port, ZN => n4744);
   U2072 : AOI22_X1 port map( A1 => n5579, A2 => registers_21_18_port, B1 => 
                           n5582, B2 => registers_26_18_port, ZN => n4743);
   U2073 : AOI22_X1 port map( A1 => n5588, A2 => registers_15_18_port, B1 => 
                           n5591, B2 => registers_31_18_port, ZN => n4742);
   U2074 : AOI22_X1 port map( A1 => n5568, A2 => registers_5_19_port, B1 => 
                           n5578, B2 => registers_8_19_port, ZN => n4726);
   U2075 : AOI22_X1 port map( A1 => n5580, A2 => registers_21_19_port, B1 => 
                           n5583, B2 => registers_26_19_port, ZN => n4725);
   U2076 : AOI22_X1 port map( A1 => n5589, A2 => registers_15_19_port, B1 => 
                           n5592, B2 => registers_31_19_port, ZN => n4724);
   U2077 : AOI22_X1 port map( A1 => n5569, A2 => registers_5_20_port, B1 => 
                           n4489, B2 => registers_8_20_port, ZN => n4708);
   U2078 : AOI22_X1 port map( A1 => n4483, A2 => registers_21_20_port, B1 => 
                           n5581, B2 => registers_26_20_port, ZN => n4707);
   U2079 : AOI22_X1 port map( A1 => n5587, A2 => registers_15_20_port, B1 => 
                           n5590, B2 => registers_31_20_port, ZN => n4706);
   U2080 : AOI22_X1 port map( A1 => n5570, A2 => registers_5_21_port, B1 => 
                           n5577, B2 => registers_8_21_port, ZN => n4690);
   U2081 : AOI22_X1 port map( A1 => n5579, A2 => registers_21_21_port, B1 => 
                           n5581, B2 => registers_26_21_port, ZN => n4689);
   U2082 : AOI22_X1 port map( A1 => n5587, A2 => registers_15_21_port, B1 => 
                           n5590, B2 => registers_31_21_port, ZN => n4688);
   U2083 : AOI22_X1 port map( A1 => n5571, A2 => registers_5_22_port, B1 => 
                           n5578, B2 => registers_8_22_port, ZN => n4672);
   U2084 : AOI22_X1 port map( A1 => n5580, A2 => registers_21_22_port, B1 => 
                           n5582, B2 => registers_26_22_port, ZN => n4671);
   U2085 : AOI22_X1 port map( A1 => n5588, A2 => registers_15_22_port, B1 => 
                           n5591, B2 => registers_31_22_port, ZN => n4670);
   U2086 : AOI22_X1 port map( A1 => n5572, A2 => registers_5_23_port, B1 => 
                           n4489, B2 => registers_8_23_port, ZN => n4654);
   U2087 : AOI22_X1 port map( A1 => n4483, A2 => registers_21_23_port, B1 => 
                           n5582, B2 => registers_26_23_port, ZN => n4653);
   U2088 : AOI22_X1 port map( A1 => n5588, A2 => registers_15_23_port, B1 => 
                           n5591, B2 => registers_31_23_port, ZN => n4652);
   U2089 : AOI22_X1 port map( A1 => n5569, A2 => registers_5_24_port, B1 => 
                           n5577, B2 => registers_8_24_port, ZN => n4636);
   U2090 : AOI22_X1 port map( A1 => n5579, A2 => registers_21_24_port, B1 => 
                           n5583, B2 => registers_26_24_port, ZN => n4635);
   U2091 : AOI22_X1 port map( A1 => n5589, A2 => registers_15_24_port, B1 => 
                           n5592, B2 => registers_31_24_port, ZN => n4634);
   U2092 : AOI22_X1 port map( A1 => n5570, A2 => registers_5_25_port, B1 => 
                           n5578, B2 => registers_8_25_port, ZN => n4618);
   U2093 : AOI22_X1 port map( A1 => n5580, A2 => registers_21_25_port, B1 => 
                           n5581, B2 => registers_26_25_port, ZN => n4617);
   U2094 : AOI22_X1 port map( A1 => n5587, A2 => registers_15_25_port, B1 => 
                           n5590, B2 => registers_31_25_port, ZN => n4616);
   U2095 : AOI22_X1 port map( A1 => n5571, A2 => registers_5_26_port, B1 => 
                           n4489, B2 => registers_8_26_port, ZN => n4600);
   U2096 : AOI22_X1 port map( A1 => n4483, A2 => registers_21_26_port, B1 => 
                           n5583, B2 => registers_26_26_port, ZN => n4599);
   U2097 : AOI22_X1 port map( A1 => n5589, A2 => registers_15_26_port, B1 => 
                           n5592, B2 => registers_31_26_port, ZN => n4598);
   U2098 : AOI22_X1 port map( A1 => n5572, A2 => registers_5_27_port, B1 => 
                           n5577, B2 => registers_8_27_port, ZN => n4582);
   U2099 : AOI22_X1 port map( A1 => n5579, A2 => registers_21_27_port, B1 => 
                           n5582, B2 => registers_26_27_port, ZN => n4581);
   U2100 : AOI22_X1 port map( A1 => n5588, A2 => registers_15_27_port, B1 => 
                           n5591, B2 => registers_31_27_port, ZN => n4580);
   U2101 : AOI22_X1 port map( A1 => n5573, A2 => registers_5_28_port, B1 => 
                           n5578, B2 => registers_8_28_port, ZN => n4564);
   U2102 : AOI22_X1 port map( A1 => n5580, A2 => registers_21_28_port, B1 => 
                           n5583, B2 => registers_26_28_port, ZN => n4563);
   U2103 : AOI22_X1 port map( A1 => n5589, A2 => registers_15_28_port, B1 => 
                           n5592, B2 => registers_31_28_port, ZN => n4562);
   U2104 : AOI22_X1 port map( A1 => n5574, A2 => registers_5_29_port, B1 => 
                           n4489, B2 => registers_8_29_port, ZN => n4546);
   U2106 : AOI22_X1 port map( A1 => n4483, A2 => registers_21_29_port, B1 => 
                           n5581, B2 => registers_26_29_port, ZN => n4545);
   U2107 : AOI22_X1 port map( A1 => n5587, A2 => registers_15_29_port, B1 => 
                           n5590, B2 => registers_31_29_port, ZN => n4544);
   U2108 : AOI22_X1 port map( A1 => n5575, A2 => registers_5_30_port, B1 => 
                           n5577, B2 => registers_8_30_port, ZN => n4528);
   U2109 : AOI22_X1 port map( A1 => n5579, A2 => registers_21_30_port, B1 => 
                           n5581, B2 => registers_26_30_port, ZN => n4527);
   U2110 : AOI22_X1 port map( A1 => n5587, A2 => registers_15_30_port, B1 => 
                           n5590, B2 => registers_31_30_port, ZN => n4526);
   U2111 : AOI22_X1 port map( A1 => n5576, A2 => registers_5_31_port, B1 => 
                           n5578, B2 => registers_8_31_port, ZN => n4487);
   U2112 : AOI22_X1 port map( A1 => n5580, A2 => registers_21_31_port, B1 => 
                           n5582, B2 => registers_26_31_port, ZN => n4482);
   U2113 : AOI22_X1 port map( A1 => n5588, A2 => registers_15_31_port, B1 => 
                           n5591, B2 => net108162, ZN => n4477);
   U2114 : OAI221_X1 port map( B1 => n2387, B2 => n5541, C1 => n5311, C2 => 
                           n5549, A => n5089, ZN => n5062);
   U2115 : AOI22_X1 port map( A1 => n5551, A2 => registers_17_0_port, B1 => 
                           n5559, B2 => registers_13_0_port, ZN => n5089);
   U2116 : OAI221_X1 port map( B1 => n4223, B2 => n5542, C1 => n2288, C2 => 
                           n5548, A => n5051, ZN => n5044);
   U2117 : AOI22_X1 port map( A1 => n5552, A2 => registers_17_1_port, B1 => 
                           n5555, B2 => registers_13_1_port, ZN => n5051);
   U2118 : OAI221_X1 port map( B1 => n4242, B2 => n4490, C1 => n2289, C2 => 
                           n5546, A => n5033, ZN => n5026);
   U2119 : AOI22_X1 port map( A1 => n4493, A2 => registers_17_2_port, B1 => 
                           n5559, B2 => registers_13_2_port, ZN => n5033);
   U2120 : OAI221_X1 port map( B1 => n4261, B2 => n5541, C1 => n2290, C2 => 
                           n5549, A => n5015, ZN => n5008);
   U2121 : AOI22_X1 port map( A1 => n5551, A2 => registers_17_3_port, B1 => 
                           n5556, B2 => registers_13_3_port, ZN => n5015);
   U2122 : OAI221_X1 port map( B1 => n4280, B2 => n5542, C1 => n2291, C2 => 
                           n5544, A => n4997, ZN => n4990);
   U2123 : AOI22_X1 port map( A1 => n5552, A2 => registers_17_4_port, B1 => 
                           n5557, B2 => registers_13_4_port, ZN => n4997);
   U2124 : OAI221_X1 port map( B1 => n4299, B2 => n4490, C1 => n2292, C2 => 
                           n5545, A => n4979, ZN => n4972);
   U2125 : AOI22_X1 port map( A1 => n4493, A2 => registers_17_5_port, B1 => 
                           n5556, B2 => registers_13_5_port, ZN => n4979);
   U2126 : OAI221_X1 port map( B1 => n4318, B2 => n5541, C1 => n2293, C2 => 
                           n5546, A => n4961, ZN => n4954);
   U2127 : AOI22_X1 port map( A1 => n5551, A2 => registers_17_6_port, B1 => 
                           n5558, B2 => registers_13_6_port, ZN => n4961);
   U2128 : OAI221_X1 port map( B1 => n4337, B2 => n5542, C1 => n2294, C2 => 
                           n5545, A => n4943, ZN => n4936);
   U2129 : AOI22_X1 port map( A1 => n5552, A2 => registers_17_7_port, B1 => 
                           n5560, B2 => registers_13_7_port, ZN => n4943);
   U2130 : OAI221_X1 port map( B1 => n4356, B2 => n4490, C1 => n2295, C2 => 
                           n5547, A => n4925, ZN => n4918);
   U2131 : AOI22_X1 port map( A1 => n4493, A2 => registers_17_8_port, B1 => 
                           n5555, B2 => registers_13_8_port, ZN => n4925);
   U2132 : OAI221_X1 port map( B1 => n4375, B2 => n5541, C1 => n2296, C2 => 
                           n5548, A => n4907, ZN => n4900);
   U2133 : AOI22_X1 port map( A1 => n5551, A2 => registers_17_9_port, B1 => 
                           n5557, B2 => registers_13_9_port, ZN => n4907);
   U2134 : OAI221_X1 port map( B1 => n4394, B2 => n5542, C1 => n2297, C2 => 
                           n5549, A => n4889, ZN => n4882);
   U2135 : AOI22_X1 port map( A1 => n5552, A2 => registers_17_10_port, B1 => 
                           n5557, B2 => registers_13_10_port, ZN => n4889);
   U2136 : OAI221_X1 port map( B1 => n4416, B2 => n4490, C1 => n2298, C2 => 
                           n5550, A => n4871, ZN => n4864);
   U2137 : AOI22_X1 port map( A1 => n4493, A2 => registers_17_11_port, B1 => 
                           n5558, B2 => registers_13_11_port, ZN => n4871);
   U2138 : OAI221_X1 port map( B1 => n4431, B2 => n5541, C1 => n2299, C2 => 
                           n5544, A => n4853, ZN => n4846);
   U2139 : AOI22_X1 port map( A1 => n5551, A2 => registers_17_12_port, B1 => 
                           n5559, B2 => registers_13_12_port, ZN => n4853);
   U2140 : OAI221_X1 port map( B1 => n5103, B2 => n5542, C1 => n2300, C2 => 
                           n5545, A => n4835, ZN => n4828);
   U2141 : AOI22_X1 port map( A1 => n5552, A2 => registers_17_13_port, B1 => 
                           n5559, B2 => registers_13_13_port, ZN => n4835);
   U2142 : OAI221_X1 port map( B1 => n5104, B2 => n4490, C1 => n2301, C2 => 
                           n5546, A => n4817, ZN => n4810);
   U2143 : AOI22_X1 port map( A1 => n4493, A2 => registers_17_14_port, B1 => 
                           n5557, B2 => registers_13_14_port, ZN => n4817);
   U2144 : OAI221_X1 port map( B1 => n5105, B2 => n5541, C1 => n2302, C2 => 
                           n5545, A => n4799, ZN => n4792);
   U2145 : AOI22_X1 port map( A1 => n5551, A2 => registers_17_15_port, B1 => 
                           n5558, B2 => registers_13_15_port, ZN => n4799);
   U2146 : OAI221_X1 port map( B1 => n5106, B2 => n5542, C1 => n2303, C2 => 
                           n5547, A => n4781, ZN => n4774);
   U2147 : AOI22_X1 port map( A1 => n5552, A2 => registers_17_16_port, B1 => 
                           n5559, B2 => registers_13_16_port, ZN => n4781);
   U2148 : OAI221_X1 port map( B1 => n5107, B2 => n4490, C1 => n2304, C2 => 
                           n5548, A => n4763, ZN => n4756);
   U2149 : AOI22_X1 port map( A1 => n4493, A2 => registers_17_17_port, B1 => 
                           n5559, B2 => registers_13_17_port, ZN => n4763);
   U2150 : OAI221_X1 port map( B1 => n5108, B2 => n5541, C1 => n2305, C2 => 
                           n5549, A => n4745, ZN => n4738);
   U2151 : AOI22_X1 port map( A1 => n5551, A2 => registers_17_18_port, B1 => 
                           n5560, B2 => registers_13_18_port, ZN => n4745);
   U2152 : OAI221_X1 port map( B1 => n5109, B2 => n5542, C1 => n2306, C2 => 
                           n5550, A => n4727, ZN => n4720);
   U2153 : AOI22_X1 port map( A1 => n5552, A2 => registers_17_19_port, B1 => 
                           n5560, B2 => registers_13_19_port, ZN => n4727);
   U2154 : OAI221_X1 port map( B1 => n5110, B2 => n4490, C1 => n2307, C2 => 
                           n5544, A => n4709, ZN => n4702);
   U2155 : AOI22_X1 port map( A1 => n4493, A2 => registers_17_20_port, B1 => 
                           n5560, B2 => registers_13_20_port, ZN => n4709);
   U2156 : OAI221_X1 port map( B1 => n5111, B2 => n5541, C1 => n2308, C2 => 
                           n5544, A => n4691, ZN => n4684);
   U2157 : AOI22_X1 port map( A1 => n5551, A2 => registers_17_21_port, B1 => 
                           n5560, B2 => registers_13_21_port, ZN => n4691);
   U2158 : OAI221_X1 port map( B1 => n5112, B2 => n5542, C1 => n2309, C2 => 
                           n5549, A => n4673, ZN => n4666);
   U2159 : AOI22_X1 port map( A1 => n5552, A2 => registers_17_22_port, B1 => 
                           n5560, B2 => registers_13_22_port, ZN => n4673);
   U2160 : OAI221_X1 port map( B1 => n5113, B2 => n4490, C1 => n2310, C2 => 
                           n5546, A => n4655, ZN => n4648);
   U2161 : AOI22_X1 port map( A1 => n4493, A2 => registers_17_23_port, B1 => 
                           n5555, B2 => registers_13_23_port, ZN => n4655);
   U2162 : OAI221_X1 port map( B1 => n5114, B2 => n5541, C1 => n2311, C2 => 
                           n5550, A => n4637, ZN => n4630);
   U2163 : AOI22_X1 port map( A1 => n5551, A2 => registers_17_24_port, B1 => 
                           n5555, B2 => registers_13_24_port, ZN => n4637);
   U2164 : OAI221_X1 port map( B1 => n5115, B2 => n5542, C1 => n2312, C2 => 
                           n5544, A => n4619, ZN => n4612);
   U2165 : AOI22_X1 port map( A1 => n5552, A2 => registers_17_25_port, B1 => 
                           n5556, B2 => registers_13_25_port, ZN => n4619);
   U2166 : OAI221_X1 port map( B1 => n5116, B2 => n4490, C1 => n2313, C2 => 
                           n5546, A => n4601, ZN => n4594);
   U2167 : AOI22_X1 port map( A1 => n4493, A2 => registers_17_26_port, B1 => 
                           n5557, B2 => registers_13_26_port, ZN => n4601);
   U2168 : OAI221_X1 port map( B1 => n5117, B2 => n5541, C1 => n2314, C2 => 
                           n5548, A => n4583, ZN => n4576);
   U2169 : AOI22_X1 port map( A1 => n5551, A2 => registers_17_27_port, B1 => 
                           n5556, B2 => registers_13_27_port, ZN => n4583);
   U2170 : OAI221_X1 port map( B1 => n5118, B2 => n5542, C1 => n2315, C2 => 
                           n5550, A => n4565, ZN => n4558);
   U2171 : AOI22_X1 port map( A1 => n5552, A2 => registers_17_28_port, B1 => 
                           n5555, B2 => registers_13_28_port, ZN => n4565);
   U2172 : OAI221_X1 port map( B1 => n5119, B2 => n4490, C1 => n2316, C2 => 
                           n5547, A => n4547, ZN => n4540);
   U2173 : AOI22_X1 port map( A1 => n4493, A2 => registers_17_29_port, B1 => 
                           n5557, B2 => registers_13_29_port, ZN => n4547);
   U2174 : OAI221_X1 port map( B1 => n5120, B2 => n5541, C1 => n2317, C2 => 
                           n5547, A => n4529, ZN => n4522);
   U2175 : AOI22_X1 port map( A1 => n5551, A2 => registers_17_30_port, B1 => 
                           n5558, B2 => registers_13_30_port, ZN => n4529);
   U2176 : OAI221_X1 port map( B1 => n5121, B2 => n5542, C1 => n2318, C2 => 
                           n5550, A => n4492, ZN => n4471);
   U2177 : AOI22_X1 port map( A1 => n5552, A2 => registers_17_31_port, B1 => 
                           n5558, B2 => registers_13_31_port, ZN => n4492);
   U2178 : INV_X1 port map( A => wr_addr(3), ZN => n1767);
   U2179 : INV_X1 port map( A => n1706, ZN => n3966);
   U2180 : AOI22_X1 port map( A1 => d_in(23), A2 => n5953, B1 => n5956, B2 => 
                           registers_2_23_port, ZN => n1706);
   U2181 : OAI21_X1 port map( B1 => n2700, B2 => n5314, A => n4186, ZN => n3008
                           );
   U2182 : AOI22_X1 port map( A1 => d_link(12), A2 => n5694, B1 => n5696, B2 =>
                           d_in(12), ZN => n4186);
   U2183 : AND3_X1 port map( A1 => wr_addr(3), A2 => wr_addr(2), A3 => n2320, 
                           ZN => n2629);
   U2184 : AND3_X1 port map( A1 => n1768, A2 => n1767, A3 => wr_addr(2), ZN => 
                           n1804);
   U2185 : AND3_X1 port map( A1 => wr_addr(2), A2 => n1767, A3 => n2320, ZN => 
                           n2355);
   U2186 : AND3_X1 port map( A1 => wr_addr(2), A2 => n1768, A3 => wr_addr(3), 
                           ZN => n2078);
   U2187 : AND3_X1 port map( A1 => wr_addr(3), A2 => n1766, A3 => n2320, ZN => 
                           n2492);
   U2188 : AND3_X1 port map( A1 => n1768, A2 => n1766, A3 => wr_addr(3), ZN => 
                           n1941);
   U2189 : OAI21_X1 port map( B1 => n2700, B2 => n5315, A => n4319, ZN => n2994
                           );
   U2190 : AOI22_X1 port map( A1 => d_link(5), A2 => n5691, B1 => n5697, B2 => 
                           d_in(5), ZN => n4319);
   U2191 : INV_X1 port map( A => wr_addr(2), ZN => n1766);
   U2192 : INV_X1 port map( A => wr_addr(0), ZN => n2664);
   U2193 : INV_X1 port map( A => wr_addr(1), ZN => n2699);
   U2194 : AND2_X1 port map( A1 => link_en, A2 => n2700, ZN => n2703);
   U2195 : NAND4_X1 port map( A1 => n4419, A2 => n4420, A3 => n4421, A4 => 
                           n4422, ZN => n2983);
   U2196 : AOI221_X1 port map( B1 => registers_31_0_port, B2 => n5595, C1 => 
                           n5468, C2 => d_out2_0_port, A => n4444, ZN => n4419)
                           ;
   U2197 : AOI221_X1 port map( B1 => n5680, B2 => registers_9_0_port, C1 => 
                           n4423, C2 => registers_12_0_port, A => n4424, ZN => 
                           n4422);
   U2198 : AOI221_X1 port map( B1 => n5669, B2 => registers_5_0_port, C1 => 
                           n5677, C2 => registers_8_0_port, A => n4432, ZN => 
                           n4421);
   U2199 : NAND4_X1 port map( A1 => n4396, A2 => n4397, A3 => n4398, A4 => 
                           n4399, ZN => n2985);
   U2200 : AOI221_X1 port map( B1 => registers_31_1_port, B2 => n5597, C1 => 
                           n5466, C2 => d_out2_1_port, A => n4415, ZN => n4396)
                           ;
   U2201 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_1_port, C1 => 
                           n5663, C2 => registers_30_1_port, A => n4413, ZN => 
                           n4397);
   U2202 : AOI221_X1 port map( B1 => n5678, B2 => registers_8_1_port, C1 => 
                           n2741, C2 => registers_20_1_port, A => n4411, ZN => 
                           n4398);
   U2203 : NAND4_X1 port map( A1 => n4377, A2 => n4378, A3 => n4379, A4 => 
                           n4380, ZN => n2987);
   U2204 : AOI221_X1 port map( B1 => registers_31_2_port, B2 => n5596, C1 => 
                           n5467, C2 => d_out2_2_port, A => n4393, ZN => n4377)
                           ;
   U2205 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_2_port, C1 => 
                           n2746, C2 => registers_30_2_port, A => n4392, ZN => 
                           n4378);
   U2206 : AOI221_X1 port map( B1 => n2740, B2 => registers_8_2_port, C1 => 
                           n2741, C2 => registers_20_2_port, A => n4391, ZN => 
                           n4379);
   U2207 : NAND4_X1 port map( A1 => n4358, A2 => n4359, A3 => n4360, A4 => 
                           n4361, ZN => n2989);
   U2208 : AOI221_X1 port map( B1 => registers_31_3_port, B2 => n5596, C1 => 
                           n5467, C2 => d_out2_3_port, A => n4374, ZN => n4358)
                           ;
   U2209 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_3_port, C1 => 
                           n2746, C2 => registers_30_3_port, A => n4373, ZN => 
                           n4359);
   U2210 : AOI221_X1 port map( B1 => n5677, B2 => registers_8_3_port, C1 => 
                           n2741, C2 => registers_20_3_port, A => n4372, ZN => 
                           n4360);
   U2211 : NAND4_X1 port map( A1 => n4339, A2 => n4340, A3 => n4341, A4 => 
                           n4342, ZN => n2991);
   U2212 : AOI221_X1 port map( B1 => registers_31_4_port, B2 => n5595, C1 => 
                           n5468, C2 => d_out2_4_port, A => n4355, ZN => n4339)
                           ;
   U2213 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_4_port, C1 => 
                           n5663, C2 => registers_30_4_port, A => n4354, ZN => 
                           n4340);
   U2214 : AOI221_X1 port map( B1 => n5678, B2 => registers_8_4_port, C1 => 
                           n2741, C2 => registers_20_4_port, A => n4353, ZN => 
                           n4341);
   U2215 : NAND4_X1 port map( A1 => n4320, A2 => n4321, A3 => n4322, A4 => 
                           n4323, ZN => n2993);
   U2216 : AOI221_X1 port map( B1 => registers_31_5_port, B2 => n5597, C1 => 
                           n5468, C2 => d_out2_5_port, A => n4336, ZN => n4320)
                           ;
   U2217 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_5_port, C1 => 
                           n5664, C2 => registers_30_5_port, A => n4335, ZN => 
                           n4321);
   U2218 : AOI221_X1 port map( B1 => n2740, B2 => registers_8_5_port, C1 => 
                           n2741, C2 => registers_20_5_port, A => n4334, ZN => 
                           n4322);
   U2219 : NAND4_X1 port map( A1 => n4301, A2 => n4302, A3 => n4303, A4 => 
                           n4304, ZN => n2995);
   U2220 : AOI221_X1 port map( B1 => registers_31_6_port, B2 => n5597, C1 => 
                           n5466, C2 => d_out2_6_port, A => n4317, ZN => n4301)
                           ;
   U2221 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_6_port, C1 => 
                           n2746, C2 => registers_30_6_port, A => n4316, ZN => 
                           n4302);
   U2222 : AOI221_X1 port map( B1 => n5677, B2 => registers_8_6_port, C1 => 
                           n2741, C2 => registers_20_6_port, A => n4315, ZN => 
                           n4303);
   U2223 : NAND4_X1 port map( A1 => n4282, A2 => n4283, A3 => n4284, A4 => 
                           n4285, ZN => n2997);
   U2224 : AOI221_X1 port map( B1 => registers_31_7_port, B2 => n5596, C1 => 
                           n5467, C2 => d_out2_7_port, A => n4298, ZN => n4282)
                           ;
   U2225 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_7_port, C1 => 
                           n5663, C2 => registers_30_7_port, A => n4297, ZN => 
                           n4283);
   U2226 : AOI221_X1 port map( B1 => n5678, B2 => registers_8_7_port, C1 => 
                           n2741, C2 => registers_20_7_port, A => n4296, ZN => 
                           n4284);
   U2227 : NAND4_X1 port map( A1 => n4263, A2 => n4264, A3 => n4265, A4 => 
                           n4266, ZN => n2999);
   U2228 : AOI221_X1 port map( B1 => registers_31_8_port, B2 => n5595, C1 => 
                           n5466, C2 => d_out2_8_port, A => n4279, ZN => n4263)
                           ;
   U2229 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_8_port, C1 => 
                           n5664, C2 => registers_30_8_port, A => n4278, ZN => 
                           n4264);
   U2230 : AOI221_X1 port map( B1 => n2740, B2 => registers_8_8_port, C1 => 
                           n2741, C2 => registers_20_8_port, A => n4277, ZN => 
                           n4265);
   U2231 : NAND4_X1 port map( A1 => n4244, A2 => n4245, A3 => n4246, A4 => 
                           n4247, ZN => n3001);
   U2232 : AOI221_X1 port map( B1 => registers_31_9_port, B2 => n5595, C1 => 
                           n5468, C2 => d_out2_9_port, A => n4260, ZN => n4244)
                           ;
   U2233 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_9_port, C1 => 
                           n2746, C2 => registers_30_9_port, A => n4259, ZN => 
                           n4245);
   U2234 : AOI221_X1 port map( B1 => n5677, B2 => registers_8_9_port, C1 => 
                           n2741, C2 => registers_20_9_port, A => n4258, ZN => 
                           n4246);
   U2235 : NAND4_X1 port map( A1 => n4225, A2 => n4226, A3 => n4227, A4 => 
                           n4228, ZN => n3003);
   U2236 : AOI221_X1 port map( B1 => registers_31_10_port, B2 => n5597, C1 => 
                           n5466, C2 => d_out2_10_port, A => n4241, ZN => n4225
                           );
   U2237 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_10_port, C1 => 
                           n5663, C2 => registers_30_10_port, A => n4240, ZN =>
                           n4226);
   U2238 : AOI221_X1 port map( B1 => n5678, B2 => registers_8_10_port, C1 => 
                           n2741, C2 => registers_20_10_port, A => n4239, ZN =>
                           n4227);
   U2239 : NAND4_X1 port map( A1 => n4206, A2 => n4207, A3 => n4208, A4 => 
                           n4209, ZN => n3005);
   U2240 : AOI221_X1 port map( B1 => registers_31_11_port, B2 => n5596, C1 => 
                           n5467, C2 => d_out2_11_port, A => n4222, ZN => n4206
                           );
   U2241 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_11_port, C1 => 
                           n5664, C2 => registers_30_11_port, A => n4221, ZN =>
                           n4207);
   U2242 : AOI221_X1 port map( B1 => n2740, B2 => registers_8_11_port, C1 => 
                           n2741, C2 => registers_20_11_port, A => n4220, ZN =>
                           n4208);
   U2243 : NAND4_X1 port map( A1 => n4187, A2 => n4188, A3 => n4189, A4 => 
                           n4190, ZN => n3007);
   U2244 : AOI221_X1 port map( B1 => registers_31_12_port, B2 => n5596, C1 => 
                           n5467, C2 => d_out2_12_port, A => n4203, ZN => n4187
                           );
   U2245 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_12_port, C1 => 
                           n2746, C2 => registers_30_12_port, A => n4202, ZN =>
                           n4188);
   U2246 : AOI221_X1 port map( B1 => n5677, B2 => registers_8_12_port, C1 => 
                           n2741, C2 => registers_20_12_port, A => n4201, ZN =>
                           n4189);
   U2247 : NAND4_X1 port map( A1 => n4168, A2 => n4169, A3 => n4170, A4 => 
                           n4171, ZN => n3009);
   U2248 : AOI221_X1 port map( B1 => registers_31_13_port, B2 => n5595, C1 => 
                           n5468, C2 => d_out2_13_port, A => n4184, ZN => n4168
                           );
   U2249 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_13_port, C1 => 
                           n5663, C2 => registers_30_13_port, A => n4183, ZN =>
                           n4169);
   U2250 : AOI221_X1 port map( B1 => n5678, B2 => registers_8_13_port, C1 => 
                           n2741, C2 => registers_20_13_port, A => n4182, ZN =>
                           n4170);
   U2251 : NAND4_X1 port map( A1 => n4149, A2 => n4150, A3 => n4151, A4 => 
                           n4152, ZN => n3011);
   U2252 : AOI221_X1 port map( B1 => registers_31_14_port, B2 => n5597, C1 => 
                           n5468, C2 => d_out2_14_port, A => n4165, ZN => n4149
                           );
   U2253 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_14_port, C1 => 
                           n5664, C2 => registers_30_14_port, A => n4164, ZN =>
                           n4150);
   U2254 : AOI221_X1 port map( B1 => n2740, B2 => registers_8_14_port, C1 => 
                           n2741, C2 => registers_20_14_port, A => n4163, ZN =>
                           n4151);
   U2255 : NAND4_X1 port map( A1 => n4130, A2 => n4131, A3 => n4132, A4 => 
                           n4133, ZN => n3013);
   U2256 : AOI221_X1 port map( B1 => registers_31_15_port, B2 => n5597, C1 => 
                           n5466, C2 => d_out2_15_port, A => n4146, ZN => n4130
                           );
   U2257 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_15_port, C1 => 
                           n2746, C2 => registers_30_15_port, A => n4145, ZN =>
                           n4131);
   U2258 : AOI221_X1 port map( B1 => n5677, B2 => registers_8_15_port, C1 => 
                           n2741, C2 => registers_20_15_port, A => n4144, ZN =>
                           n4132);
   U2259 : NAND4_X1 port map( A1 => n4111, A2 => n4112, A3 => n4113, A4 => 
                           n4114, ZN => n3015);
   U2260 : AOI221_X1 port map( B1 => registers_31_16_port, B2 => n5596, C1 => 
                           n5467, C2 => d_out2_16_port, A => n4127, ZN => n4111
                           );
   U2261 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_16_port, C1 => 
                           n5663, C2 => registers_30_16_port, A => n4126, ZN =>
                           n4112);
   U2262 : AOI221_X1 port map( B1 => n5678, B2 => registers_8_16_port, C1 => 
                           n2741, C2 => registers_20_16_port, A => n4125, ZN =>
                           n4113);
   U2263 : NAND4_X1 port map( A1 => n4092, A2 => n4093, A3 => n4094, A4 => 
                           n4095, ZN => n3017);
   U2264 : AOI221_X1 port map( B1 => registers_31_17_port, B2 => n5595, C1 => 
                           n5466, C2 => d_out2_17_port, A => n4108, ZN => n4092
                           );
   U2265 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_17_port, C1 => 
                           n5664, C2 => registers_30_17_port, A => n4107, ZN =>
                           n4093);
   U2266 : AOI221_X1 port map( B1 => n2740, B2 => registers_8_17_port, C1 => 
                           n2741, C2 => registers_20_17_port, A => n4106, ZN =>
                           n4094);
   U2267 : NAND4_X1 port map( A1 => n4073, A2 => n4074, A3 => n4075, A4 => 
                           n4076, ZN => n3019);
   U2268 : AOI221_X1 port map( B1 => registers_31_18_port, B2 => n5595, C1 => 
                           n5468, C2 => d_out2_18_port, A => n4089, ZN => n4073
                           );
   U2269 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_18_port, C1 => 
                           n2746, C2 => registers_30_18_port, A => n4088, ZN =>
                           n4074);
   U2270 : AOI221_X1 port map( B1 => n5677, B2 => registers_8_18_port, C1 => 
                           n2741, C2 => registers_20_18_port, A => n4087, ZN =>
                           n4075);
   U2271 : NAND4_X1 port map( A1 => n4054, A2 => n4055, A3 => n4056, A4 => 
                           n4057, ZN => n3021);
   U2272 : AOI221_X1 port map( B1 => registers_31_19_port, B2 => n5597, C1 => 
                           n5466, C2 => d_out2_19_port, A => n4070, ZN => n4054
                           );
   U2273 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_19_port, C1 => 
                           n5663, C2 => registers_30_19_port, A => n4069, ZN =>
                           n4055);
   U2274 : AOI221_X1 port map( B1 => n5678, B2 => registers_8_19_port, C1 => 
                           n2741, C2 => registers_20_19_port, A => n4068, ZN =>
                           n4056);
   U2275 : NAND4_X1 port map( A1 => n4035, A2 => n4036, A3 => n4037, A4 => 
                           n4038, ZN => n3023);
   U2276 : AOI221_X1 port map( B1 => registers_31_20_port, B2 => n5596, C1 => 
                           n5467, C2 => d_out2_20_port, A => n4051, ZN => n4035
                           );
   U2277 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_20_port, C1 => 
                           n5664, C2 => registers_30_20_port, A => n4050, ZN =>
                           n4036);
   U2278 : AOI221_X1 port map( B1 => n2740, B2 => registers_8_20_port, C1 => 
                           n2741, C2 => registers_20_20_port, A => n4049, ZN =>
                           n4037);
   U2279 : NAND4_X1 port map( A1 => n4016, A2 => n4017, A3 => n4018, A4 => 
                           n4019, ZN => n3025);
   U2280 : AOI221_X1 port map( B1 => registers_31_21_port, B2 => n5596, C1 => 
                           n5467, C2 => d_out2_21_port, A => n4032, ZN => n4016
                           );
   U2281 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_21_port, C1 => 
                           n2746, C2 => registers_30_21_port, A => n4031, ZN =>
                           n4017);
   U2282 : AOI221_X1 port map( B1 => n5677, B2 => registers_8_21_port, C1 => 
                           n2741, C2 => registers_20_21_port, A => n4030, ZN =>
                           n4018);
   U2283 : NAND4_X1 port map( A1 => n2910, A2 => n2911, A3 => n2912, A4 => 
                           n2913, ZN => n3027);
   U2284 : AOI221_X1 port map( B1 => registers_31_22_port, B2 => n5595, C1 => 
                           n5468, C2 => d_out2_22_port, A => n4013, ZN => n2910
                           );
   U2285 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_22_port, C1 => 
                           n5663, C2 => registers_30_22_port, A => n4012, ZN =>
                           n2911);
   U2286 : AOI221_X1 port map( B1 => n5678, B2 => registers_8_22_port, C1 => 
                           n2741, C2 => registers_20_22_port, A => n4011, ZN =>
                           n2912);
   U2287 : NAND4_X1 port map( A1 => n2891, A2 => n2892, A3 => n2893, A4 => 
                           n2894, ZN => n3029);
   U2288 : AOI221_X1 port map( B1 => registers_31_23_port, B2 => n5597, C1 => 
                           n5468, C2 => d_out2_23_port, A => n2907, ZN => n2891
                           );
   U2289 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_23_port, C1 => 
                           n5664, C2 => registers_30_23_port, A => n2906, ZN =>
                           n2892);
   U2290 : AOI221_X1 port map( B1 => n2740, B2 => registers_8_23_port, C1 => 
                           n2741, C2 => registers_20_23_port, A => n2905, ZN =>
                           n2893);
   U2291 : NAND4_X1 port map( A1 => n2872, A2 => n2873, A3 => n2874, A4 => 
                           n2875, ZN => n3031);
   U2292 : AOI221_X1 port map( B1 => registers_31_24_port, B2 => n5597, C1 => 
                           n5466, C2 => d_out2_24_port, A => n2888, ZN => n2872
                           );
   U2293 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_24_port, C1 => 
                           n2746, C2 => registers_30_24_port, A => n2887, ZN =>
                           n2873);
   U2294 : AOI221_X1 port map( B1 => n5677, B2 => registers_8_24_port, C1 => 
                           n2741, C2 => registers_20_24_port, A => n2886, ZN =>
                           n2874);
   U2295 : NAND4_X1 port map( A1 => n2853, A2 => n2854, A3 => n2855, A4 => 
                           n2856, ZN => n3033);
   U2296 : AOI221_X1 port map( B1 => registers_31_25_port, B2 => n5596, C1 => 
                           n5467, C2 => d_out2_25_port, A => n2869, ZN => n2853
                           );
   U2297 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_25_port, C1 => 
                           n5663, C2 => registers_30_25_port, A => n2868, ZN =>
                           n2854);
   U2298 : AOI221_X1 port map( B1 => n5678, B2 => registers_8_25_port, C1 => 
                           n2741, C2 => registers_20_25_port, A => n2867, ZN =>
                           n2855);
   U2299 : NAND4_X1 port map( A1 => n2834, A2 => n2835, A3 => n2836, A4 => 
                           n2837, ZN => n3035);
   U2300 : AOI221_X1 port map( B1 => registers_31_26_port, B2 => n5595, C1 => 
                           n5466, C2 => d_out2_26_port, A => n2850, ZN => n2834
                           );
   U2301 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_26_port, C1 => 
                           n5664, C2 => registers_30_26_port, A => n2849, ZN =>
                           n2835);
   U2302 : AOI221_X1 port map( B1 => n2740, B2 => registers_8_26_port, C1 => 
                           n2741, C2 => registers_20_26_port, A => n2848, ZN =>
                           n2836);
   U2303 : NAND4_X1 port map( A1 => n2815, A2 => n2816, A3 => n2817, A4 => 
                           n2818, ZN => n3037);
   U2304 : AOI221_X1 port map( B1 => registers_31_27_port, B2 => n5595, C1 => 
                           n5468, C2 => d_out2_27_port, A => n2831, ZN => n2815
                           );
   U2305 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_27_port, C1 => 
                           n2746, C2 => registers_30_27_port, A => n2830, ZN =>
                           n2816);
   U2306 : AOI221_X1 port map( B1 => n5677, B2 => registers_8_27_port, C1 => 
                           n2741, C2 => registers_20_27_port, A => n2829, ZN =>
                           n2817);
   U2307 : NAND4_X1 port map( A1 => n2796, A2 => n2797, A3 => n2798, A4 => 
                           n2799, ZN => n3039);
   U2308 : AOI221_X1 port map( B1 => registers_31_28_port, B2 => n5597, C1 => 
                           n5466, C2 => d_out2_28_port, A => n2812, ZN => n2796
                           );
   U2309 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_28_port, C1 => 
                           n5663, C2 => registers_30_28_port, A => n2811, ZN =>
                           n2797);
   U2310 : AOI221_X1 port map( B1 => n5678, B2 => registers_8_28_port, C1 => 
                           n2741, C2 => registers_20_28_port, A => n2810, ZN =>
                           n2798);
   U2311 : NAND4_X1 port map( A1 => n2777, A2 => n2778, A3 => n2779, A4 => 
                           n2780, ZN => n3041);
   U2312 : AOI221_X1 port map( B1 => registers_31_29_port, B2 => n5596, C1 => 
                           n5467, C2 => d_out2_29_port, A => n2793, ZN => n2777
                           );
   U2313 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_29_port, C1 => 
                           n5664, C2 => registers_30_29_port, A => n2792, ZN =>
                           n2778);
   U2314 : AOI221_X1 port map( B1 => n2740, B2 => registers_8_29_port, C1 => 
                           n2741, C2 => registers_20_29_port, A => n2791, ZN =>
                           n2779);
   U2315 : NAND4_X1 port map( A1 => n2758, A2 => n2759, A3 => n2760, A4 => 
                           n2761, ZN => n3043);
   U2316 : AOI221_X1 port map( B1 => registers_31_30_port, B2 => n5596, C1 => 
                           n5467, C2 => d_out2_30_port, A => n2774, ZN => n2758
                           );
   U2317 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_30_port, C1 => 
                           n2746, C2 => registers_30_30_port, A => n2773, ZN =>
                           n2759);
   U2318 : AOI221_X1 port map( B1 => n5677, B2 => registers_8_30_port, C1 => 
                           n2741, C2 => registers_20_30_port, A => n2772, ZN =>
                           n2760);
   U2319 : NAND4_X1 port map( A1 => n2705, A2 => n2706, A3 => n2707, A4 => 
                           n2708, ZN => n3045);
   U2320 : AOI221_X1 port map( B1 => n5595, B2 => net108162, C1 => n5468, C2 =>
                           d_out2_31_port, A => n2753, ZN => n2705);
   U2321 : AOI221_X1 port map( B1 => n2745, B2 => registers_27_31_port, C1 => 
                           n5663, C2 => registers_30_31_port, A => n2747, ZN =>
                           n2706);
   U2322 : AOI221_X1 port map( B1 => n5678, B2 => registers_8_31_port, C1 => 
                           n2741, C2 => registers_20_31_port, A => n2742, ZN =>
                           n2707);
   U2323 : NAND4_X1 port map( A1 => n5058, A2 => n5059, A3 => n5060, A4 => 
                           n5061, ZN => n2951);
   U2324 : AOI221_X1 port map( B1 => n5508, B2 => registers_7_0_port, C1 => 
                           n5510, C2 => registers_16_0_port, A => n5099, ZN => 
                           n5058);
   U2325 : AOI221_X1 port map( B1 => n5513, B2 => registers_3_0_port, C1 => 
                           n5517, C2 => registers_2_0_port, A => n5098, ZN => 
                           n5059);
   U2326 : NOR4_X1 port map( A1 => n5091, A2 => n5092, A3 => n5093, A4 => n5094
                           , ZN => n5060);
   U2327 : NAND4_X1 port map( A1 => n5040, A2 => n5041, A3 => n5042, A4 => 
                           n5043, ZN => n2952);
   U2328 : AOI221_X1 port map( B1 => n5509, B2 => registers_7_1_port, C1 => 
                           n5511, C2 => registers_16_1_port, A => n5057, ZN => 
                           n5040);
   U2329 : AOI221_X1 port map( B1 => n5514, B2 => registers_3_1_port, C1 => 
                           n5521, C2 => registers_2_1_port, A => n5056, ZN => 
                           n5041);
   U2330 : NOR4_X1 port map( A1 => n5052, A2 => n5053, A3 => n5054, A4 => n5055
                           , ZN => n5042);
   U2331 : NAND4_X1 port map( A1 => n5022, A2 => n5023, A3 => n5024, A4 => 
                           n5025, ZN => n2953);
   U2332 : AOI221_X1 port map( B1 => n5507, B2 => registers_7_2_port, C1 => 
                           n4514, C2 => registers_16_2_port, A => n5039, ZN => 
                           n5022);
   U2333 : AOI221_X1 port map( B1 => n5512, B2 => registers_3_2_port, C1 => 
                           n5522, C2 => registers_2_2_port, A => n5038, ZN => 
                           n5023);
   U2334 : NOR4_X1 port map( A1 => n5034, A2 => n5035, A3 => n5036, A4 => n5037
                           , ZN => n5024);
   U2335 : NAND4_X1 port map( A1 => n5004, A2 => n5005, A3 => n5006, A4 => 
                           n5007, ZN => n2954);
   U2336 : AOI221_X1 port map( B1 => n5507, B2 => registers_7_3_port, C1 => 
                           n5510, C2 => registers_16_3_port, A => n5021, ZN => 
                           n5004);
   U2337 : AOI221_X1 port map( B1 => n5512, B2 => registers_3_3_port, C1 => 
                           n5518, C2 => registers_2_3_port, A => n5020, ZN => 
                           n5005);
   U2338 : NOR4_X1 port map( A1 => n5016, A2 => n5017, A3 => n5018, A4 => n5019
                           , ZN => n5006);
   U2339 : NAND4_X1 port map( A1 => n4986, A2 => n4987, A3 => n4988, A4 => 
                           n4989, ZN => n2955);
   U2340 : AOI221_X1 port map( B1 => n5508, B2 => registers_7_4_port, C1 => 
                           n5511, C2 => registers_16_4_port, A => n5003, ZN => 
                           n4986);
   U2341 : AOI221_X1 port map( B1 => n5513, B2 => registers_3_4_port, C1 => 
                           n5519, C2 => registers_2_4_port, A => n5002, ZN => 
                           n4987);
   U2342 : NOR4_X1 port map( A1 => n4998, A2 => n4999, A3 => n5000, A4 => n5001
                           , ZN => n4988);
   U2343 : NAND4_X1 port map( A1 => n4968, A2 => n4969, A3 => n4970, A4 => 
                           n4971, ZN => n2956);
   U2344 : AOI221_X1 port map( B1 => n5508, B2 => registers_7_5_port, C1 => 
                           n4514, C2 => registers_16_5_port, A => n4985, ZN => 
                           n4968);
   U2345 : AOI221_X1 port map( B1 => n5513, B2 => registers_3_5_port, C1 => 
                           n5518, C2 => registers_2_5_port, A => n4984, ZN => 
                           n4969);
   U2346 : NOR4_X1 port map( A1 => n4980, A2 => n4981, A3 => n4982, A4 => n4983
                           , ZN => n4970);
   U2347 : NAND4_X1 port map( A1 => n4950, A2 => n4951, A3 => n4952, A4 => 
                           n4953, ZN => n2957);
   U2348 : AOI221_X1 port map( B1 => n5509, B2 => registers_7_6_port, C1 => 
                           n5510, C2 => registers_16_6_port, A => n4967, ZN => 
                           n4950);
   U2349 : AOI221_X1 port map( B1 => n5514, B2 => registers_3_6_port, C1 => 
                           n5520, C2 => registers_2_6_port, A => n4966, ZN => 
                           n4951);
   U2350 : NOR4_X1 port map( A1 => n4962, A2 => n4963, A3 => n4964, A4 => n4965
                           , ZN => n4952);
   U2351 : NAND4_X1 port map( A1 => n4932, A2 => n4933, A3 => n4934, A4 => 
                           n4935, ZN => n2958);
   U2352 : AOI221_X1 port map( B1 => n5507, B2 => registers_7_7_port, C1 => 
                           n5511, C2 => registers_16_7_port, A => n4949, ZN => 
                           n4932);
   U2353 : AOI221_X1 port map( B1 => n5512, B2 => registers_3_7_port, C1 => 
                           n5522, C2 => registers_2_7_port, A => n4948, ZN => 
                           n4933);
   U2354 : NOR4_X1 port map( A1 => n4944, A2 => n4945, A3 => n4946, A4 => n4947
                           , ZN => n4934);
   U2355 : NAND4_X1 port map( A1 => n4914, A2 => n4915, A3 => n4916, A4 => 
                           n4917, ZN => n2959);
   U2356 : AOI221_X1 port map( B1 => n5509, B2 => registers_7_8_port, C1 => 
                           n4514, C2 => registers_16_8_port, A => n4931, ZN => 
                           n4914);
   U2357 : AOI221_X1 port map( B1 => n5514, B2 => registers_3_8_port, C1 => 
                           n5520, C2 => registers_2_8_port, A => n4930, ZN => 
                           n4915);
   U2358 : NOR4_X1 port map( A1 => n4926, A2 => n4927, A3 => n4928, A4 => n4929
                           , ZN => n4916);
   U2359 : NAND4_X1 port map( A1 => n4896, A2 => n4897, A3 => n4898, A4 => 
                           n4899, ZN => n2960);
   U2360 : AOI221_X1 port map( B1 => n5508, B2 => registers_7_9_port, C1 => 
                           n5510, C2 => registers_16_9_port, A => n4913, ZN => 
                           n4896);
   U2361 : AOI221_X1 port map( B1 => n5513, B2 => registers_3_9_port, C1 => 
                           n5519, C2 => registers_2_9_port, A => n4912, ZN => 
                           n4897);
   U2362 : NOR4_X1 port map( A1 => n4908, A2 => n4909, A3 => n4910, A4 => n4911
                           , ZN => n4898);
   U2363 : NAND4_X1 port map( A1 => n4878, A2 => n4879, A3 => n4880, A4 => 
                           n4881, ZN => n2961);
   U2364 : AOI221_X1 port map( B1 => n5509, B2 => registers_7_10_port, C1 => 
                           n5511, C2 => registers_16_10_port, A => n4895, ZN =>
                           n4878);
   U2365 : AOI221_X1 port map( B1 => n5514, B2 => registers_3_10_port, C1 => 
                           n5519, C2 => registers_2_10_port, A => n4894, ZN => 
                           n4879);
   U2366 : NOR4_X1 port map( A1 => n4890, A2 => n4891, A3 => n4892, A4 => n4893
                           , ZN => n4880);
   U2367 : NAND4_X1 port map( A1 => n4860, A2 => n4861, A3 => n4862, A4 => 
                           n4863, ZN => n2962);
   U2368 : AOI221_X1 port map( B1 => n5507, B2 => registers_7_11_port, C1 => 
                           n4514, C2 => registers_16_11_port, A => n4877, ZN =>
                           n4860);
   U2369 : AOI221_X1 port map( B1 => n5512, B2 => registers_3_11_port, C1 => 
                           n5520, C2 => registers_2_11_port, A => n4876, ZN => 
                           n4861);
   U2370 : NOR4_X1 port map( A1 => n4872, A2 => n4873, A3 => n4874, A4 => n4875
                           , ZN => n4862);
   U2371 : NAND4_X1 port map( A1 => n4842, A2 => n4843, A3 => n4844, A4 => 
                           n4845, ZN => n2963);
   U2372 : AOI221_X1 port map( B1 => n5507, B2 => registers_7_12_port, C1 => 
                           n5510, C2 => registers_16_12_port, A => n4859, ZN =>
                           n4842);
   U2373 : AOI221_X1 port map( B1 => n5512, B2 => registers_3_12_port, C1 => 
                           n5521, C2 => registers_2_12_port, A => n4858, ZN => 
                           n4843);
   U2374 : NOR4_X1 port map( A1 => n4854, A2 => n4855, A3 => n4856, A4 => n4857
                           , ZN => n4844);
   U2375 : NAND4_X1 port map( A1 => n4824, A2 => n4825, A3 => n4826, A4 => 
                           n4827, ZN => n2964);
   U2376 : AOI221_X1 port map( B1 => n5508, B2 => registers_7_13_port, C1 => 
                           n5511, C2 => registers_16_13_port, A => n4841, ZN =>
                           n4824);
   U2377 : AOI221_X1 port map( B1 => n5513, B2 => registers_3_13_port, C1 => 
                           n5521, C2 => registers_2_13_port, A => n4840, ZN => 
                           n4825);
   U2378 : NOR4_X1 port map( A1 => n4836, A2 => n4837, A3 => n4838, A4 => n4839
                           , ZN => n4826);
   U2379 : NAND4_X1 port map( A1 => n4806, A2 => n4807, A3 => n4808, A4 => 
                           n4809, ZN => n2965);
   U2380 : AOI221_X1 port map( B1 => n5508, B2 => registers_7_14_port, C1 => 
                           n4514, C2 => registers_16_14_port, A => n4823, ZN =>
                           n4806);
   U2381 : AOI221_X1 port map( B1 => n5513, B2 => registers_3_14_port, C1 => 
                           n5519, C2 => registers_2_14_port, A => n4822, ZN => 
                           n4807);
   U2382 : NOR4_X1 port map( A1 => n4818, A2 => n4819, A3 => n4820, A4 => n4821
                           , ZN => n4808);
   U2383 : NAND4_X1 port map( A1 => n4788, A2 => n4789, A3 => n4790, A4 => 
                           n4791, ZN => n2966);
   U2384 : AOI221_X1 port map( B1 => n5509, B2 => registers_7_15_port, C1 => 
                           n5510, C2 => registers_16_15_port, A => n4805, ZN =>
                           n4788);
   U2385 : AOI221_X1 port map( B1 => n5514, B2 => registers_3_15_port, C1 => 
                           n5520, C2 => registers_2_15_port, A => n4804, ZN => 
                           n4789);
   U2386 : NOR4_X1 port map( A1 => n4800, A2 => n4801, A3 => n4802, A4 => n4803
                           , ZN => n4790);
   U2387 : NAND4_X1 port map( A1 => n4770, A2 => n4771, A3 => n4772, A4 => 
                           n4773, ZN => n2967);
   U2388 : AOI221_X1 port map( B1 => n5507, B2 => registers_7_16_port, C1 => 
                           n5511, C2 => registers_16_16_port, A => n4787, ZN =>
                           n4770);
   U2389 : AOI221_X1 port map( B1 => n5512, B2 => registers_3_16_port, C1 => 
                           n5521, C2 => registers_2_16_port, A => n4786, ZN => 
                           n4771);
   U2390 : NOR4_X1 port map( A1 => n4782, A2 => n4783, A3 => n4784, A4 => n4785
                           , ZN => n4772);
   U2391 : NAND4_X1 port map( A1 => n4752, A2 => n4753, A3 => n4754, A4 => 
                           n4755, ZN => n2968);
   U2392 : AOI221_X1 port map( B1 => n5509, B2 => registers_7_17_port, C1 => 
                           n4514, C2 => registers_16_17_port, A => n4769, ZN =>
                           n4752);
   U2393 : AOI221_X1 port map( B1 => n5514, B2 => registers_3_17_port, C1 => 
                           n5521, C2 => registers_2_17_port, A => n4768, ZN => 
                           n4753);
   U2394 : NOR4_X1 port map( A1 => n4764, A2 => n4765, A3 => n4766, A4 => n4767
                           , ZN => n4754);
   U2395 : NAND4_X1 port map( A1 => n4734, A2 => n4735, A3 => n4736, A4 => 
                           n4737, ZN => n2969);
   U2396 : AOI221_X1 port map( B1 => n5508, B2 => registers_7_18_port, C1 => 
                           n5510, C2 => registers_16_18_port, A => n4751, ZN =>
                           n4734);
   U2397 : AOI221_X1 port map( B1 => n5513, B2 => registers_3_18_port, C1 => 
                           n5522, C2 => registers_2_18_port, A => n4750, ZN => 
                           n4735);
   U2398 : NOR4_X1 port map( A1 => n4746, A2 => n4747, A3 => n4748, A4 => n4749
                           , ZN => n4736);
   U2399 : NAND4_X1 port map( A1 => n4716, A2 => n4717, A3 => n4718, A4 => 
                           n4719, ZN => n2970);
   U2400 : AOI221_X1 port map( B1 => n5509, B2 => registers_7_19_port, C1 => 
                           n5511, C2 => registers_16_19_port, A => n4733, ZN =>
                           n4716);
   U2401 : AOI221_X1 port map( B1 => n5514, B2 => registers_3_19_port, C1 => 
                           n5522, C2 => registers_2_19_port, A => n4732, ZN => 
                           n4717);
   U2402 : NOR4_X1 port map( A1 => n4728, A2 => n4729, A3 => n4730, A4 => n4731
                           , ZN => n4718);
   U2403 : NAND4_X1 port map( A1 => n4698, A2 => n4699, A3 => n4700, A4 => 
                           n4701, ZN => n2971);
   U2404 : AOI221_X1 port map( B1 => n5507, B2 => registers_7_20_port, C1 => 
                           n4514, C2 => registers_16_20_port, A => n4715, ZN =>
                           n4698);
   U2405 : AOI221_X1 port map( B1 => n5512, B2 => registers_3_20_port, C1 => 
                           n5522, C2 => registers_2_20_port, A => n4714, ZN => 
                           n4699);
   U2406 : NOR4_X1 port map( A1 => n4710, A2 => n4711, A3 => n4712, A4 => n4713
                           , ZN => n4700);
   U2407 : NAND4_X1 port map( A1 => n4680, A2 => n4681, A3 => n4682, A4 => 
                           n4683, ZN => n2972);
   U2408 : AOI221_X1 port map( B1 => n5507, B2 => registers_7_21_port, C1 => 
                           n5510, C2 => registers_16_21_port, A => n4697, ZN =>
                           n4680);
   U2409 : AOI221_X1 port map( B1 => n5512, B2 => registers_3_21_port, C1 => 
                           n5522, C2 => registers_2_21_port, A => n4696, ZN => 
                           n4681);
   U2410 : NOR4_X1 port map( A1 => n4692, A2 => n4693, A3 => n4694, A4 => n4695
                           , ZN => n4682);
   U2411 : NAND4_X1 port map( A1 => n4662, A2 => n4663, A3 => n4664, A4 => 
                           n4665, ZN => n2973);
   U2412 : AOI221_X1 port map( B1 => n5508, B2 => registers_7_22_port, C1 => 
                           n5511, C2 => registers_16_22_port, A => n4679, ZN =>
                           n4662);
   U2413 : AOI221_X1 port map( B1 => n5513, B2 => registers_3_22_port, C1 => 
                           n5517, C2 => registers_2_22_port, A => n4678, ZN => 
                           n4663);
   U2414 : NOR4_X1 port map( A1 => n4674, A2 => n4675, A3 => n4676, A4 => n4677
                           , ZN => n4664);
   U2415 : NAND4_X1 port map( A1 => n4644, A2 => n4645, A3 => n4646, A4 => 
                           n4647, ZN => n2974);
   U2416 : AOI221_X1 port map( B1 => n5508, B2 => registers_7_23_port, C1 => 
                           n4514, C2 => registers_16_23_port, A => n4661, ZN =>
                           n4644);
   U2417 : AOI221_X1 port map( B1 => n5513, B2 => registers_3_23_port, C1 => 
                           n5521, C2 => registers_2_23_port, A => n4660, ZN => 
                           n4645);
   U2418 : NOR4_X1 port map( A1 => n4656, A2 => n4657, A3 => n4658, A4 => n4659
                           , ZN => n4646);
   U2419 : NAND4_X1 port map( A1 => n4626, A2 => n4627, A3 => n4628, A4 => 
                           n4629, ZN => n2975);
   U2420 : AOI221_X1 port map( B1 => n5509, B2 => registers_7_24_port, C1 => 
                           n5510, C2 => registers_16_24_port, A => n4643, ZN =>
                           n4626);
   U2421 : AOI221_X1 port map( B1 => n5514, B2 => registers_3_24_port, C1 => 
                           n5517, C2 => registers_2_24_port, A => n4642, ZN => 
                           n4627);
   U2422 : NOR4_X1 port map( A1 => n4638, A2 => n4639, A3 => n4640, A4 => n4641
                           , ZN => n4628);
   U2423 : NAND4_X1 port map( A1 => n4608, A2 => n4609, A3 => n4610, A4 => 
                           n4611, ZN => n2976);
   U2424 : AOI221_X1 port map( B1 => n5507, B2 => registers_7_25_port, C1 => 
                           n5511, C2 => registers_16_25_port, A => n4625, ZN =>
                           n4608);
   U2425 : AOI221_X1 port map( B1 => n5512, B2 => registers_3_25_port, C1 => 
                           n5518, C2 => registers_2_25_port, A => n4624, ZN => 
                           n4609);
   U2426 : NOR4_X1 port map( A1 => n4620, A2 => n4621, A3 => n4622, A4 => n4623
                           , ZN => n4610);
   U2427 : NAND4_X1 port map( A1 => n4590, A2 => n4591, A3 => n4592, A4 => 
                           n4593, ZN => n2977);
   U2428 : AOI221_X1 port map( B1 => n5509, B2 => registers_7_26_port, C1 => 
                           n4514, C2 => registers_16_26_port, A => n4607, ZN =>
                           n4590);
   U2429 : AOI221_X1 port map( B1 => n5514, B2 => registers_3_26_port, C1 => 
                           n5519, C2 => registers_2_26_port, A => n4606, ZN => 
                           n4591);
   U2430 : NOR4_X1 port map( A1 => n4602, A2 => n4603, A3 => n4604, A4 => n4605
                           , ZN => n4592);
   U2431 : NAND4_X1 port map( A1 => n4572, A2 => n4573, A3 => n4574, A4 => 
                           n4575, ZN => n2978);
   U2432 : AOI221_X1 port map( B1 => n5508, B2 => registers_7_27_port, C1 => 
                           n5510, C2 => registers_16_27_port, A => n4589, ZN =>
                           n4572);
   U2433 : AOI221_X1 port map( B1 => n5513, B2 => registers_3_27_port, C1 => 
                           n5518, C2 => registers_2_27_port, A => n4588, ZN => 
                           n4573);
   U2434 : NOR4_X1 port map( A1 => n4584, A2 => n4585, A3 => n4586, A4 => n4587
                           , ZN => n4574);
   U2435 : NAND4_X1 port map( A1 => n4554, A2 => n4555, A3 => n4556, A4 => 
                           n4557, ZN => n2979);
   U2436 : AOI221_X1 port map( B1 => n5509, B2 => registers_7_28_port, C1 => 
                           n5511, C2 => registers_16_28_port, A => n4571, ZN =>
                           n4554);
   U2437 : AOI221_X1 port map( B1 => n5514, B2 => registers_3_28_port, C1 => 
                           n5517, C2 => registers_2_28_port, A => n4570, ZN => 
                           n4555);
   U2438 : NOR4_X1 port map( A1 => n4566, A2 => n4567, A3 => n4568, A4 => n4569
                           , ZN => n4556);
   U2439 : NAND4_X1 port map( A1 => n4536, A2 => n4537, A3 => n4538, A4 => 
                           n4539, ZN => n2980);
   U2440 : AOI221_X1 port map( B1 => n5507, B2 => registers_7_29_port, C1 => 
                           n4514, C2 => registers_16_29_port, A => n4553, ZN =>
                           n4536);
   U2441 : AOI221_X1 port map( B1 => n5512, B2 => registers_3_29_port, C1 => 
                           n5517, C2 => registers_2_29_port, A => n4552, ZN => 
                           n4537);
   U2442 : NOR4_X1 port map( A1 => n4548, A2 => n4549, A3 => n4550, A4 => n4551
                           , ZN => n4538);
   U2443 : NAND4_X1 port map( A1 => n4518, A2 => n4519, A3 => n4520, A4 => 
                           n4521, ZN => n2981);
   U2444 : AOI221_X1 port map( B1 => n5507, B2 => registers_7_30_port, C1 => 
                           n5510, C2 => registers_16_30_port, A => n4535, ZN =>
                           n4518);
   U2445 : AOI221_X1 port map( B1 => n5512, B2 => registers_3_30_port, C1 => 
                           n5519, C2 => registers_2_30_port, A => n4534, ZN => 
                           n4519);
   U2446 : NOR4_X1 port map( A1 => n4530, A2 => n4531, A3 => n4532, A4 => n4533
                           , ZN => n4520);
   U2447 : NAND4_X1 port map( A1 => n4467, A2 => n4468, A3 => n4469, A4 => 
                           n4470, ZN => n2982);
   U2448 : AOI221_X1 port map( B1 => n5508, B2 => registers_7_31_port, C1 => 
                           n5511, C2 => registers_16_31_port, A => n4515, ZN =>
                           n4467);
   U2449 : AOI221_X1 port map( B1 => n5513, B2 => registers_3_31_port, C1 => 
                           n5520, C2 => registers_2_31_port, A => n4510, ZN => 
                           n4468);
   U2450 : NOR4_X1 port map( A1 => n4495, A2 => n4496, A3 => n4497, A4 => n4498
                           , ZN => n4469);
   U2451 : OAI21_X1 port map( B1 => n2700, B2 => n5316, A => n4417, ZN => n2984
                           );
   U2452 : AOI22_X1 port map( A1 => d_link(0), A2 => n5689, B1 => n5697, B2 => 
                           d_in(0), ZN => n4417);
   U2453 : OAI21_X1 port map( B1 => n2700, B2 => n5317, A => n4395, ZN => n2986
                           );
   U2454 : AOI22_X1 port map( A1 => d_link(1), A2 => n5690, B1 => n5698, B2 => 
                           d_in(1), ZN => n4395);
   U2455 : OAI21_X1 port map( B1 => n2700, B2 => n5318, A => n4376, ZN => n2988
                           );
   U2456 : AOI22_X1 port map( A1 => d_link(2), A2 => n5690, B1 => n5696, B2 => 
                           d_in(2), ZN => n4376);
   U2457 : OAI21_X1 port map( B1 => n2700, B2 => n5319, A => n4357, ZN => n2990
                           );
   U2458 : AOI22_X1 port map( A1 => d_link(3), A2 => n5691, B1 => n5696, B2 => 
                           d_in(3), ZN => n4357);
   U2459 : OAI21_X1 port map( B1 => n2700, B2 => n5320, A => n4338, ZN => n2992
                           );
   U2460 : AOI22_X1 port map( A1 => d_link(4), A2 => n5692, B1 => n5697, B2 => 
                           d_in(4), ZN => n4338);
   U2461 : OAI21_X1 port map( B1 => n2700, B2 => n5321, A => n4300, ZN => n2996
                           );
   U2462 : AOI22_X1 port map( A1 => d_link(6), A2 => n5693, B1 => n5698, B2 => 
                           d_in(6), ZN => n4300);
   U2463 : OAI21_X1 port map( B1 => n2700, B2 => n5322, A => n4281, ZN => n2998
                           );
   U2464 : AOI22_X1 port map( A1 => d_link(7), A2 => n5689, B1 => n5696, B2 => 
                           d_in(7), ZN => n4281);
   U2465 : OAI21_X1 port map( B1 => n2700, B2 => n5323, A => n4262, ZN => n3000
                           );
   U2466 : AOI22_X1 port map( A1 => d_link(8), A2 => n5689, B1 => n5698, B2 => 
                           d_in(8), ZN => n4262);
   U2467 : OAI21_X1 port map( B1 => n2700, B2 => n5324, A => n4243, ZN => n3002
                           );
   U2468 : AOI22_X1 port map( A1 => d_link(9), A2 => n5692, B1 => n5697, B2 => 
                           d_in(9), ZN => n4243);
   U2469 : OAI21_X1 port map( B1 => n2700, B2 => n5325, A => n4224, ZN => n3004
                           );
   U2470 : AOI22_X1 port map( A1 => d_link(10), A2 => n5692, B1 => n5698, B2 =>
                           d_in(10), ZN => n4224);
   U2471 : OAI21_X1 port map( B1 => n2700, B2 => n5326, A => n4205, ZN => n3006
                           );
   U2472 : AOI22_X1 port map( A1 => d_link(11), A2 => n5693, B1 => n5696, B2 =>
                           d_in(11), ZN => n4205);
   U2473 : OAI21_X1 port map( B1 => n2700, B2 => n5327, A => n4167, ZN => n3010
                           );
   U2474 : AOI22_X1 port map( A1 => d_link(13), A2 => n5694, B1 => n5697, B2 =>
                           d_in(13), ZN => n4167);
   U2475 : OAI21_X1 port map( B1 => n2700, B2 => n5328, A => n4148, ZN => n3012
                           );
   U2476 : AOI22_X1 port map( A1 => d_link(14), A2 => n5692, B1 => n5697, B2 =>
                           d_in(14), ZN => n4148);
   U2477 : OAI21_X1 port map( B1 => n2700, B2 => n5329, A => n4129, ZN => n3014
                           );
   U2478 : AOI22_X1 port map( A1 => d_link(15), A2 => n5693, B1 => n5698, B2 =>
                           d_in(15), ZN => n4129);
   U2479 : OAI21_X1 port map( B1 => n2700, B2 => n5330, A => n4110, ZN => n3016
                           );
   U2480 : AOI22_X1 port map( A1 => d_link(16), A2 => n5694, B1 => n5696, B2 =>
                           d_in(16), ZN => n4110);
   U2481 : OAI21_X1 port map( B1 => n2700, B2 => n5331, A => n4091, ZN => n3018
                           );
   U2482 : AOI22_X1 port map( A1 => d_link(17), A2 => n5694, B1 => n5698, B2 =>
                           d_in(17), ZN => n4091);
   U2483 : OAI21_X1 port map( B1 => n2700, B2 => n5332, A => n4072, ZN => n3020
                           );
   U2484 : AOI22_X1 port map( A1 => d_link(18), A2 => n5695, B1 => n5697, B2 =>
                           d_in(18), ZN => n4072);
   U2485 : OAI21_X1 port map( B1 => n2700, B2 => n5333, A => n4053, ZN => n3022
                           );
   U2486 : AOI22_X1 port map( A1 => d_link(19), A2 => n5695, B1 => n5698, B2 =>
                           d_in(19), ZN => n4053);
   U2487 : OAI21_X1 port map( B1 => n2700, B2 => n5334, A => n4034, ZN => n3024
                           );
   U2488 : AOI22_X1 port map( A1 => d_link(20), A2 => n5695, B1 => n5696, B2 =>
                           d_in(20), ZN => n4034);
   U2489 : OAI21_X1 port map( B1 => n2700, B2 => n5335, A => n4015, ZN => n3026
                           );
   U2490 : AOI22_X1 port map( A1 => d_link(21), A2 => n5695, B1 => n5696, B2 =>
                           d_in(21), ZN => n4015);
   U2491 : OAI21_X1 port map( B1 => n2700, B2 => n5336, A => n2909, ZN => n3028
                           );
   U2492 : AOI22_X1 port map( A1 => d_link(22), A2 => n5689, B1 => n5697, B2 =>
                           d_in(22), ZN => n2909);
   U2493 : OAI21_X1 port map( B1 => n2700, B2 => n5337, A => n2890, ZN => n3030
                           );
   U2494 : AOI22_X1 port map( A1 => d_link(23), A2 => n5690, B1 => n5697, B2 =>
                           d_in(23), ZN => n2890);
   U2495 : OAI21_X1 port map( B1 => n2700, B2 => n5338, A => n2871, ZN => n3032
                           );
   U2496 : AOI22_X1 port map( A1 => d_link(24), A2 => n5689, B1 => n5698, B2 =>
                           d_in(24), ZN => n2871);
   U2497 : OAI21_X1 port map( B1 => n2700, B2 => n5339, A => n2852, ZN => n3034
                           );
   U2498 : AOI22_X1 port map( A1 => d_link(25), A2 => n5691, B1 => n5696, B2 =>
                           d_in(25), ZN => n2852);
   U2499 : OAI21_X1 port map( B1 => n2700, B2 => n5340, A => n2833, ZN => n3036
                           );
   U2500 : AOI22_X1 port map( A1 => d_link(26), A2 => n5691, B1 => n5698, B2 =>
                           d_in(26), ZN => n2833);
   U2501 : OAI21_X1 port map( B1 => n2700, B2 => n5341, A => n2814, ZN => n3038
                           );
   U2502 : AOI22_X1 port map( A1 => d_link(27), A2 => n5690, B1 => n5697, B2 =>
                           d_in(27), ZN => n2814);
   U2503 : OAI21_X1 port map( B1 => n2700, B2 => n5342, A => n2795, ZN => n3040
                           );
   U2504 : AOI22_X1 port map( A1 => d_link(28), A2 => n5692, B1 => n5698, B2 =>
                           d_in(28), ZN => n2795);
   U2505 : OAI21_X1 port map( B1 => n2700, B2 => n5343, A => n2776, ZN => n3042
                           );
   U2506 : AOI22_X1 port map( A1 => d_link(29), A2 => n5695, B1 => n5696, B2 =>
                           d_in(29), ZN => n2776);
   U2507 : OAI21_X1 port map( B1 => n2700, B2 => n5344, A => n2757, ZN => n3044
                           );
   U2508 : AOI22_X1 port map( A1 => d_link(30), A2 => n5693, B1 => n5696, B2 =>
                           d_in(30), ZN => n2757);
   U2509 : OAI21_X1 port map( B1 => n2700, B2 => n5313, A => n2702, ZN => n3046
                           );
   U2510 : AOI22_X1 port map( A1 => d_link(31), A2 => n5693, B1 => n5697, B2 =>
                           d_in(31), ZN => n2702);
   U2511 : AND3_X1 port map( A1 => wr_en, A2 => en, A3 => wr_addr(4), ZN => 
                           n2320);
   U2512 : INV_X1 port map( A => d_in(0), ZN => n1692);
   U2513 : INV_X1 port map( A => d_in(23), ZN => n1646);
   U2514 : INV_X1 port map( A => d_in(1), ZN => n1690);
   U2515 : INV_X1 port map( A => d_in(2), ZN => n1688);
   U2516 : INV_X1 port map( A => d_in(3), ZN => n1686);
   U2517 : INV_X1 port map( A => d_in(4), ZN => n1684);
   U2518 : INV_X1 port map( A => d_in(5), ZN => n1682);
   U2519 : INV_X1 port map( A => d_in(6), ZN => n1680);
   U2520 : INV_X1 port map( A => d_in(7), ZN => n1678);
   U2521 : INV_X1 port map( A => d_in(8), ZN => n1676);
   U2522 : INV_X1 port map( A => d_in(9), ZN => n1674);
   U2523 : INV_X1 port map( A => d_in(10), ZN => n1672);
   U2524 : INV_X1 port map( A => d_in(11), ZN => n1670);
   U2525 : INV_X1 port map( A => d_in(12), ZN => n1668);
   U2526 : INV_X1 port map( A => d_in(13), ZN => n1666);
   U2527 : INV_X1 port map( A => d_in(14), ZN => n1664);
   U2528 : INV_X1 port map( A => d_in(15), ZN => n1662);
   U2529 : INV_X1 port map( A => d_in(16), ZN => n1660);
   U2530 : INV_X1 port map( A => d_in(17), ZN => n1658);
   U2531 : INV_X1 port map( A => d_in(18), ZN => n1656);
   U2532 : INV_X1 port map( A => d_in(19), ZN => n1654);
   U2533 : INV_X1 port map( A => d_in(20), ZN => n1652);
   U2534 : INV_X1 port map( A => d_in(21), ZN => n1650);
   U2535 : INV_X1 port map( A => d_in(22), ZN => n1648);
   U2536 : INV_X1 port map( A => d_in(24), ZN => n1644);
   U2537 : INV_X1 port map( A => d_in(25), ZN => n1642);
   U2538 : INV_X1 port map( A => d_in(26), ZN => n1640);
   U2539 : INV_X1 port map( A => d_in(27), ZN => n1638);
   U2540 : INV_X1 port map( A => d_in(28), ZN => n1636);
   U2541 : INV_X1 port map( A => d_in(29), ZN => n1634);
   U2542 : INV_X1 port map( A => d_in(30), ZN => n1632);
   U2543 : INV_X1 port map( A => d_in(31), ZN => n1629);
   U2544 : INV_X1 port map( A => n1729, ZN => n3943);
   U2545 : AOI22_X1 port map( A1 => d_in(0), A2 => n5954, B1 => n5961, B2 => 
                           registers_2_0_port, ZN => n1729);
   U2546 : INV_X1 port map( A => n1728, ZN => n3944);
   U2547 : AOI22_X1 port map( A1 => d_in(1), A2 => n5953, B1 => n5961, B2 => 
                           registers_2_1_port, ZN => n1728);
   U2548 : INV_X1 port map( A => n1727, ZN => n3945);
   U2549 : AOI22_X1 port map( A1 => d_in(2), A2 => n5954, B1 => n5960, B2 => 
                           registers_2_2_port, ZN => n1727);
   U2550 : INV_X1 port map( A => n1726, ZN => n3946);
   U2551 : AOI22_X1 port map( A1 => d_in(3), A2 => n5953, B1 => n5960, B2 => 
                           registers_2_3_port, ZN => n1726);
   U2552 : INV_X1 port map( A => n1725, ZN => n3947);
   U2553 : AOI22_X1 port map( A1 => d_in(4), A2 => n5954, B1 => n5960, B2 => 
                           registers_2_4_port, ZN => n1725);
   U2554 : INV_X1 port map( A => n1724, ZN => n3948);
   U2555 : AOI22_X1 port map( A1 => d_in(5), A2 => n5953, B1 => n5960, B2 => 
                           registers_2_5_port, ZN => n1724);
   U2556 : INV_X1 port map( A => n1723, ZN => n3949);
   U2557 : AOI22_X1 port map( A1 => d_in(6), A2 => n5954, B1 => n5960, B2 => 
                           registers_2_6_port, ZN => n1723);
   U2558 : INV_X1 port map( A => n1722, ZN => n3950);
   U2559 : AOI22_X1 port map( A1 => d_in(7), A2 => n5953, B1 => n5959, B2 => 
                           registers_2_7_port, ZN => n1722);
   U2560 : INV_X1 port map( A => n1940, ZN => n3751);
   U2561 : AOI22_X1 port map( A1 => d_in(0), A2 => n5411, B1 => n5899, B2 => 
                           registers_8_0_port, ZN => n1940);
   U2562 : INV_X1 port map( A => n1917, ZN => n3774);
   U2563 : AOI22_X1 port map( A1 => d_in(23), A2 => n5412, B1 => n5904, B2 => 
                           registers_8_23_port, ZN => n1917);
   U2564 : INV_X1 port map( A => n2111, ZN => n3592);
   U2565 : AOI22_X1 port map( A1 => d_in(1), A2 => n5398, B1 => n5855, B2 => 
                           registers_13_1_port, ZN => n2111);
   U2566 : INV_X1 port map( A => n2110, ZN => n3593);
   U2567 : AOI22_X1 port map( A1 => d_in(2), A2 => n5398, B1 => n5858, B2 => 
                           registers_13_2_port, ZN => n2110);
   U2568 : INV_X1 port map( A => n2109, ZN => n3594);
   U2569 : AOI22_X1 port map( A1 => d_in(3), A2 => n5398, B1 => n5855, B2 => 
                           registers_13_3_port, ZN => n2109);
   U2570 : INV_X1 port map( A => n2108, ZN => n3595);
   U2571 : AOI22_X1 port map( A1 => d_in(4), A2 => n5398, B1 => n5856, B2 => 
                           registers_13_4_port, ZN => n2108);
   U2572 : INV_X1 port map( A => n2107, ZN => n3596);
   U2573 : AOI22_X1 port map( A1 => d_in(5), A2 => n5398, B1 => n5855, B2 => 
                           registers_13_5_port, ZN => n2107);
   U2574 : INV_X1 port map( A => n2106, ZN => n3597);
   U2575 : AOI22_X1 port map( A1 => d_in(6), A2 => n5398, B1 => n5857, B2 => 
                           registers_13_6_port, ZN => n2106);
   U2576 : INV_X1 port map( A => n2105, ZN => n3598);
   U2577 : AOI22_X1 port map( A1 => d_in(7), A2 => n5398, B1 => n5857, B2 => 
                           registers_13_7_port, ZN => n2105);
   U2578 : INV_X1 port map( A => n2104, ZN => n3599);
   U2579 : AOI22_X1 port map( A1 => d_in(8), A2 => n5397, B1 => n5858, B2 => 
                           registers_13_8_port, ZN => n2104);
   U2580 : INV_X1 port map( A => n2103, ZN => n3600);
   U2581 : AOI22_X1 port map( A1 => d_in(9), A2 => n5397, B1 => n5858, B2 => 
                           registers_13_9_port, ZN => n2103);
   U2582 : INV_X1 port map( A => n2102, ZN => n3601);
   U2583 : AOI22_X1 port map( A1 => d_in(10), A2 => n5397, B1 => n5860, B2 => 
                           registers_13_10_port, ZN => n2102);
   U2584 : INV_X1 port map( A => n2101, ZN => n3602);
   U2585 : AOI22_X1 port map( A1 => d_in(11), A2 => n5397, B1 => n5859, B2 => 
                           registers_13_11_port, ZN => n2101);
   U2586 : INV_X1 port map( A => n2100, ZN => n3603);
   U2587 : AOI22_X1 port map( A1 => d_in(12), A2 => n5397, B1 => n5860, B2 => 
                           registers_13_12_port, ZN => n2100);
   U2588 : INV_X1 port map( A => n2099, ZN => n3604);
   U2589 : AOI22_X1 port map( A1 => d_in(13), A2 => n5397, B1 => n5854, B2 => 
                           registers_13_13_port, ZN => n2099);
   U2590 : INV_X1 port map( A => n2098, ZN => n3605);
   U2591 : AOI22_X1 port map( A1 => d_in(14), A2 => n5397, B1 => n5855, B2 => 
                           registers_13_14_port, ZN => n2098);
   U2592 : INV_X1 port map( A => n2097, ZN => n3606);
   U2593 : AOI22_X1 port map( A1 => d_in(15), A2 => n5397, B1 => n5856, B2 => 
                           registers_13_15_port, ZN => n2097);
   U2594 : INV_X1 port map( A => n2096, ZN => n3607);
   U2595 : AOI22_X1 port map( A1 => d_in(16), A2 => n5397, B1 => n5856, B2 => 
                           registers_13_16_port, ZN => n2096);
   U2596 : INV_X1 port map( A => n2095, ZN => n3608);
   U2597 : AOI22_X1 port map( A1 => d_in(17), A2 => n5397, B1 => n5857, B2 => 
                           registers_13_17_port, ZN => n2095);
   U2598 : INV_X1 port map( A => n2094, ZN => n3609);
   U2599 : AOI22_X1 port map( A1 => d_in(18), A2 => n5397, B1 => n5857, B2 => 
                           registers_13_18_port, ZN => n2094);
   U2600 : INV_X1 port map( A => n2093, ZN => n3610);
   U2601 : AOI22_X1 port map( A1 => d_in(19), A2 => n5397, B1 => n5858, B2 => 
                           registers_13_19_port, ZN => n2093);
   U2602 : INV_X1 port map( A => n2092, ZN => n3611);
   U2603 : AOI22_X1 port map( A1 => d_in(20), A2 => n5396, B1 => n5857, B2 => 
                           registers_13_20_port, ZN => n2092);
   U2604 : INV_X1 port map( A => n2091, ZN => n3612);
   U2605 : AOI22_X1 port map( A1 => d_in(21), A2 => n5396, B1 => n5860, B2 => 
                           registers_13_21_port, ZN => n2091);
   U2606 : INV_X1 port map( A => n2090, ZN => n3613);
   U2607 : AOI22_X1 port map( A1 => d_in(22), A2 => n5396, B1 => n5859, B2 => 
                           registers_13_22_port, ZN => n2090);
   U2608 : INV_X1 port map( A => n2088, ZN => n3615);
   U2609 : AOI22_X1 port map( A1 => d_in(24), A2 => n5396, B1 => n5859, B2 => 
                           registers_13_24_port, ZN => n2088);
   U2610 : INV_X1 port map( A => n2087, ZN => n3616);
   U2611 : AOI22_X1 port map( A1 => d_in(25), A2 => n5396, B1 => n5860, B2 => 
                           registers_13_25_port, ZN => n2087);
   U2612 : INV_X1 port map( A => n2086, ZN => n3617);
   U2613 : AOI22_X1 port map( A1 => d_in(26), A2 => n5396, B1 => n5854, B2 => 
                           registers_13_26_port, ZN => n2086);
   U2614 : INV_X1 port map( A => n2085, ZN => n3618);
   U2615 : AOI22_X1 port map( A1 => d_in(27), A2 => n5396, B1 => n5854, B2 => 
                           registers_13_27_port, ZN => n2085);
   U2616 : INV_X1 port map( A => n2084, ZN => n3619);
   U2617 : AOI22_X1 port map( A1 => d_in(28), A2 => n5396, B1 => n5854, B2 => 
                           registers_13_28_port, ZN => n2084);
   U2618 : INV_X1 port map( A => n2083, ZN => n3620);
   U2619 : AOI22_X1 port map( A1 => d_in(29), A2 => n5396, B1 => n5856, B2 => 
                           registers_13_29_port, ZN => n2083);
   U2620 : INV_X1 port map( A => n2082, ZN => n3621);
   U2621 : AOI22_X1 port map( A1 => d_in(30), A2 => n5396, B1 => n5856, B2 => 
                           registers_13_30_port, ZN => n2082);
   U2622 : INV_X1 port map( A => n2079, ZN => n3622);
   U2623 : AOI22_X1 port map( A1 => d_in(31), A2 => n5396, B1 => n5859, B2 => 
                           registers_13_31_port, ZN => n2079);
   U2624 : INV_X1 port map( A => n1939, ZN => n3752);
   U2625 : AOI22_X1 port map( A1 => d_in(1), A2 => n5411, B1 => n5904, B2 => 
                           registers_8_1_port, ZN => n1939);
   U2626 : INV_X1 port map( A => n1938, ZN => n3753);
   U2627 : AOI22_X1 port map( A1 => d_in(2), A2 => n5411, B1 => n5901, B2 => 
                           registers_8_2_port, ZN => n1938);
   U2628 : INV_X1 port map( A => n1937, ZN => n3754);
   U2629 : AOI22_X1 port map( A1 => d_in(3), A2 => n5411, B1 => n5902, B2 => 
                           registers_8_3_port, ZN => n1937);
   U2630 : INV_X1 port map( A => n1936, ZN => n3755);
   U2631 : AOI22_X1 port map( A1 => d_in(4), A2 => n5411, B1 => n5900, B2 => 
                           registers_8_4_port, ZN => n1936);
   U2632 : INV_X1 port map( A => n1935, ZN => n3756);
   U2633 : AOI22_X1 port map( A1 => d_in(5), A2 => n5411, B1 => n5901, B2 => 
                           registers_8_5_port, ZN => n1935);
   U2634 : INV_X1 port map( A => n1934, ZN => n3757);
   U2635 : AOI22_X1 port map( A1 => d_in(6), A2 => n5411, B1 => n5901, B2 => 
                           registers_8_6_port, ZN => n1934);
   U2636 : INV_X1 port map( A => n1933, ZN => n3758);
   U2637 : AOI22_X1 port map( A1 => d_in(7), A2 => n5411, B1 => n5905, B2 => 
                           registers_8_7_port, ZN => n1933);
   U2638 : INV_X1 port map( A => n1932, ZN => n3759);
   U2639 : AOI22_X1 port map( A1 => d_in(8), A2 => n5411, B1 => n5902, B2 => 
                           registers_8_8_port, ZN => n1932);
   U2640 : INV_X1 port map( A => n1931, ZN => n3760);
   U2641 : AOI22_X1 port map( A1 => d_in(9), A2 => n5411, B1 => n5903, B2 => 
                           registers_8_9_port, ZN => n1931);
   U2642 : INV_X1 port map( A => n1930, ZN => n3761);
   U2643 : AOI22_X1 port map( A1 => d_in(10), A2 => n5411, B1 => n5903, B2 => 
                           registers_8_10_port, ZN => n1930);
   U2644 : INV_X1 port map( A => n1929, ZN => n3762);
   U2645 : AOI22_X1 port map( A1 => d_in(11), A2 => n5411, B1 => n5904, B2 => 
                           registers_8_11_port, ZN => n1929);
   U2646 : INV_X1 port map( A => n1928, ZN => n3763);
   U2647 : AOI22_X1 port map( A1 => d_in(12), A2 => n5412, B1 => n5899, B2 => 
                           registers_8_12_port, ZN => n1928);
   U2648 : INV_X1 port map( A => n1927, ZN => n3764);
   U2649 : AOI22_X1 port map( A1 => d_in(13), A2 => n5412, B1 => n5900, B2 => 
                           registers_8_13_port, ZN => n1927);
   U2650 : INV_X1 port map( A => n1926, ZN => n3765);
   U2651 : AOI22_X1 port map( A1 => d_in(14), A2 => n5412, B1 => n5901, B2 => 
                           registers_8_14_port, ZN => n1926);
   U2652 : INV_X1 port map( A => n1925, ZN => n3766);
   U2653 : AOI22_X1 port map( A1 => d_in(15), A2 => n5412, B1 => n5900, B2 => 
                           registers_8_15_port, ZN => n1925);
   U2654 : INV_X1 port map( A => n1924, ZN => n3767);
   U2655 : AOI22_X1 port map( A1 => d_in(16), A2 => n5412, B1 => n5905, B2 => 
                           registers_8_16_port, ZN => n1924);
   U2656 : INV_X1 port map( A => n1923, ZN => n3768);
   U2657 : AOI22_X1 port map( A1 => d_in(17), A2 => n5412, B1 => n5902, B2 => 
                           registers_8_17_port, ZN => n1923);
   U2658 : INV_X1 port map( A => n1922, ZN => n3769);
   U2659 : AOI22_X1 port map( A1 => d_in(18), A2 => n5412, B1 => n5903, B2 => 
                           registers_8_18_port, ZN => n1922);
   U2660 : INV_X1 port map( A => n1921, ZN => n3770);
   U2661 : AOI22_X1 port map( A1 => d_in(19), A2 => n5412, B1 => n5902, B2 => 
                           registers_8_19_port, ZN => n1921);
   U2662 : INV_X1 port map( A => n1920, ZN => n3771);
   U2663 : AOI22_X1 port map( A1 => d_in(20), A2 => n5412, B1 => n5904, B2 => 
                           registers_8_20_port, ZN => n1920);
   U2664 : INV_X1 port map( A => n1919, ZN => n3772);
   U2665 : AOI22_X1 port map( A1 => d_in(21), A2 => n5412, B1 => n5905, B2 => 
                           registers_8_21_port, ZN => n1919);
   U2666 : INV_X1 port map( A => n1918, ZN => n3773);
   U2667 : AOI22_X1 port map( A1 => d_in(22), A2 => n5412, B1 => n5904, B2 => 
                           registers_8_22_port, ZN => n1918);
   U2668 : INV_X1 port map( A => n1916, ZN => n3775);
   U2669 : AOI22_X1 port map( A1 => d_in(24), A2 => n5413, B1 => n5905, B2 => 
                           registers_8_24_port, ZN => n1916);
   U2670 : INV_X1 port map( A => n1915, ZN => n3776);
   U2671 : AOI22_X1 port map( A1 => d_in(25), A2 => n5413, B1 => n5905, B2 => 
                           registers_8_25_port, ZN => n1915);
   U2672 : INV_X1 port map( A => n1914, ZN => n3777);
   U2673 : AOI22_X1 port map( A1 => d_in(26), A2 => n5413, B1 => n5899, B2 => 
                           registers_8_26_port, ZN => n1914);
   U2674 : INV_X1 port map( A => n1913, ZN => n3778);
   U2675 : AOI22_X1 port map( A1 => d_in(27), A2 => n5413, B1 => n5899, B2 => 
                           registers_8_27_port, ZN => n1913);
   U2676 : INV_X1 port map( A => n1912, ZN => n3779);
   U2677 : AOI22_X1 port map( A1 => d_in(28), A2 => n5413, B1 => n5899, B2 => 
                           registers_8_28_port, ZN => n1912);
   U2678 : INV_X1 port map( A => n1911, ZN => n3780);
   U2679 : AOI22_X1 port map( A1 => d_in(29), A2 => n5413, B1 => n5902, B2 => 
                           registers_8_29_port, ZN => n1911);
   U2680 : INV_X1 port map( A => n1910, ZN => n3781);
   U2681 : AOI22_X1 port map( A1 => d_in(30), A2 => n5413, B1 => n5900, B2 => 
                           registers_8_30_port, ZN => n1910);
   U2682 : INV_X1 port map( A => n1907, ZN => n3782);
   U2683 : AOI22_X1 port map( A1 => d_in(31), A2 => n5413, B1 => n5903, B2 => 
                           registers_8_31_port, ZN => n1907);
   U2684 : INV_X1 port map( A => n1721, ZN => n3951);
   U2685 : AOI22_X1 port map( A1 => d_in(8), A2 => n5954, B1 => n5959, B2 => 
                           registers_2_8_port, ZN => n1721);
   U2686 : INV_X1 port map( A => n1720, ZN => n3952);
   U2687 : AOI22_X1 port map( A1 => d_in(9), A2 => n5954, B1 => n5959, B2 => 
                           registers_2_9_port, ZN => n1720);
   U2688 : INV_X1 port map( A => n1719, ZN => n3953);
   U2689 : AOI22_X1 port map( A1 => d_in(10), A2 => n5954, B1 => n5959, B2 => 
                           registers_2_10_port, ZN => n1719);
   U2690 : INV_X1 port map( A => n1718, ZN => n3954);
   U2691 : AOI22_X1 port map( A1 => d_in(11), A2 => n5954, B1 => n5959, B2 => 
                           registers_2_11_port, ZN => n1718);
   U2692 : INV_X1 port map( A => n1717, ZN => n3955);
   U2693 : AOI22_X1 port map( A1 => d_in(12), A2 => n5954, B1 => n5958, B2 => 
                           registers_2_12_port, ZN => n1717);
   U2694 : INV_X1 port map( A => n1716, ZN => n3956);
   U2695 : AOI22_X1 port map( A1 => d_in(13), A2 => n5954, B1 => n5958, B2 => 
                           registers_2_13_port, ZN => n1716);
   U2696 : INV_X1 port map( A => n1715, ZN => n3957);
   U2697 : AOI22_X1 port map( A1 => d_in(14), A2 => n5954, B1 => n5958, B2 => 
                           registers_2_14_port, ZN => n1715);
   U2698 : INV_X1 port map( A => n1714, ZN => n3958);
   U2699 : AOI22_X1 port map( A1 => d_in(15), A2 => n5954, B1 => n5958, B2 => 
                           registers_2_15_port, ZN => n1714);
   U2700 : INV_X1 port map( A => n1713, ZN => n3959);
   U2701 : AOI22_X1 port map( A1 => d_in(16), A2 => n5954, B1 => n5958, B2 => 
                           registers_2_16_port, ZN => n1713);
   U2702 : INV_X1 port map( A => n1712, ZN => n3960);
   U2703 : AOI22_X1 port map( A1 => d_in(17), A2 => n5954, B1 => n5957, B2 => 
                           registers_2_17_port, ZN => n1712);
   U2704 : INV_X1 port map( A => n1711, ZN => n3961);
   U2705 : AOI22_X1 port map( A1 => d_in(18), A2 => n5954, B1 => n5957, B2 => 
                           registers_2_18_port, ZN => n1711);
   U2706 : INV_X1 port map( A => n1710, ZN => n3962);
   U2707 : AOI22_X1 port map( A1 => d_in(19), A2 => n5954, B1 => n5957, B2 => 
                           registers_2_19_port, ZN => n1710);
   U2708 : INV_X1 port map( A => n1709, ZN => n3963);
   U2709 : AOI22_X1 port map( A1 => d_in(20), A2 => n5953, B1 => n5957, B2 => 
                           registers_2_20_port, ZN => n1709);
   U2710 : INV_X1 port map( A => n1708, ZN => n3964);
   U2711 : AOI22_X1 port map( A1 => d_in(21), A2 => n5953, B1 => n5957, B2 => 
                           registers_2_21_port, ZN => n1708);
   U2712 : INV_X1 port map( A => n1707, ZN => n3965);
   U2713 : AOI22_X1 port map( A1 => d_in(22), A2 => n5953, B1 => n5956, B2 => 
                           registers_2_22_port, ZN => n1707);
   U2714 : INV_X1 port map( A => n1705, ZN => n3967);
   U2715 : AOI22_X1 port map( A1 => d_in(24), A2 => n5953, B1 => n5956, B2 => 
                           registers_2_24_port, ZN => n1705);
   U2716 : INV_X1 port map( A => n1704, ZN => n3968);
   U2717 : AOI22_X1 port map( A1 => d_in(25), A2 => n5953, B1 => n5956, B2 => 
                           registers_2_25_port, ZN => n1704);
   U2718 : INV_X1 port map( A => n1703, ZN => n3969);
   U2719 : AOI22_X1 port map( A1 => d_in(26), A2 => n5953, B1 => n5956, B2 => 
                           registers_2_26_port, ZN => n1703);
   U2720 : INV_X1 port map( A => n1702, ZN => n3970);
   U2721 : AOI22_X1 port map( A1 => d_in(27), A2 => n5953, B1 => n5955, B2 => 
                           registers_2_27_port, ZN => n1702);
   U2722 : INV_X1 port map( A => n1701, ZN => n3971);
   U2723 : AOI22_X1 port map( A1 => d_in(28), A2 => n5953, B1 => n5955, B2 => 
                           registers_2_28_port, ZN => n1701);
   U2724 : INV_X1 port map( A => n1700, ZN => n3972);
   U2725 : AOI22_X1 port map( A1 => d_in(29), A2 => n5953, B1 => n5955, B2 => 
                           registers_2_29_port, ZN => n1700);
   U2726 : INV_X1 port map( A => n1699, ZN => n3973);
   U2727 : AOI22_X1 port map( A1 => d_in(30), A2 => n5953, B1 => n5955, B2 => 
                           registers_2_30_port, ZN => n1699);
   U2728 : INV_X1 port map( A => n1696, ZN => n3974);
   U2729 : AOI22_X1 port map( A1 => d_in(31), A2 => n5953, B1 => n5955, B2 => 
                           registers_2_31_port, ZN => n1696);
   U2730 : OAI221_X1 port map( B1 => n2223, B2 => n5642, C1 => n2512, C2 => 
                           n5473, A => n4460, ZN => n4455);
   U2731 : AOI22_X1 port map( A1 => n5644, A2 => registers_28_0_port, B1 => 
                           n5646, B2 => registers_25_0_port, ZN => n4460);
   U2732 : OAI221_X1 port map( B1 => n2155, B2 => n5643, C1 => n2488, C2 => 
                           n5474, A => n4407, ZN => n4404);
   U2733 : AOI22_X1 port map( A1 => n5645, A2 => registers_28_1_port, B1 => 
                           n5647, B2 => registers_25_1_port, ZN => n4407);
   U2734 : OAI221_X1 port map( B1 => n2156, B2 => n5642, C1 => n2489, C2 => 
                           n5472, A => n4369, ZN => n4366);
   U2735 : AOI22_X1 port map( A1 => n5644, A2 => registers_28_3_port, B1 => 
                           n5646, B2 => registers_25_3_port, ZN => n4369);
   U2736 : OAI221_X1 port map( B1 => n2157, B2 => n5643, C1 => n2490, C2 => 
                           n5473, A => n4350, ZN => n4347);
   U2737 : AOI22_X1 port map( A1 => n5645, A2 => registers_28_4_port, B1 => 
                           n5647, B2 => registers_25_4_port, ZN => n4350);
   U2738 : OAI221_X1 port map( B1 => n2158, B2 => n5642, C1 => n2491, C2 => 
                           n5474, A => n4312, ZN => n4309);
   U2739 : AOI22_X1 port map( A1 => n5644, A2 => registers_28_6_port, B1 => 
                           n5646, B2 => registers_25_6_port, ZN => n4312);
   U2740 : OAI221_X1 port map( B1 => n2159, B2 => n5643, C1 => n2494, C2 => 
                           n5472, A => n4293, ZN => n4290);
   U2741 : AOI22_X1 port map( A1 => n5645, A2 => registers_28_7_port, B1 => 
                           n5647, B2 => registers_25_7_port, ZN => n4293);
   U2742 : OAI221_X1 port map( B1 => n2160, B2 => n5642, C1 => n2495, C2 => 
                           n5473, A => n4255, ZN => n4252);
   U2743 : AOI22_X1 port map( A1 => n5644, A2 => registers_28_9_port, B1 => 
                           n5646, B2 => registers_25_9_port, ZN => n4255);
   U2744 : OAI221_X1 port map( B1 => n2161, B2 => n5643, C1 => n2496, C2 => 
                           n5474, A => n4236, ZN => n4233);
   U2745 : AOI22_X1 port map( A1 => n5645, A2 => registers_28_10_port, B1 => 
                           n5647, B2 => registers_25_10_port, ZN => n4236);
   U2746 : OAI221_X1 port map( B1 => n2162, B2 => n5642, C1 => n2497, C2 => 
                           n5472, A => n4198, ZN => n4195);
   U2747 : AOI22_X1 port map( A1 => n5644, A2 => registers_28_12_port, B1 => 
                           n5646, B2 => registers_25_12_port, ZN => n4198);
   U2748 : OAI221_X1 port map( B1 => n2163, B2 => n5643, C1 => n2498, C2 => 
                           n5473, A => n4179, ZN => n4176);
   U2749 : AOI22_X1 port map( A1 => n5645, A2 => registers_28_13_port, B1 => 
                           n5647, B2 => registers_25_13_port, ZN => n4179);
   U2750 : OAI221_X1 port map( B1 => n2164, B2 => n5642, C1 => n2499, C2 => 
                           n5474, A => n4141, ZN => n4138);
   U2751 : AOI22_X1 port map( A1 => n5644, A2 => registers_28_15_port, B1 => 
                           n5646, B2 => registers_25_15_port, ZN => n4141);
   U2752 : OAI221_X1 port map( B1 => n2165, B2 => n5643, C1 => n2500, C2 => 
                           n5472, A => n4122, ZN => n4119);
   U2753 : AOI22_X1 port map( A1 => n5645, A2 => registers_28_16_port, B1 => 
                           n5647, B2 => registers_25_16_port, ZN => n4122);
   U2754 : OAI221_X1 port map( B1 => n2166, B2 => n5642, C1 => n2501, C2 => 
                           n5473, A => n4084, ZN => n4081);
   U2755 : AOI22_X1 port map( A1 => n5644, A2 => registers_28_18_port, B1 => 
                           n5646, B2 => registers_25_18_port, ZN => n4084);
   U2756 : OAI221_X1 port map( B1 => n2167, B2 => n5643, C1 => n2502, C2 => 
                           n5474, A => n4065, ZN => n4062);
   U2757 : AOI22_X1 port map( A1 => n5645, A2 => registers_28_19_port, B1 => 
                           n5647, B2 => registers_25_19_port, ZN => n4065);
   U2758 : OAI221_X1 port map( B1 => n2168, B2 => n5642, C1 => n2503, C2 => 
                           n5472, A => n4027, ZN => n4024);
   U2759 : AOI22_X1 port map( A1 => n5644, A2 => registers_28_21_port, B1 => 
                           n5646, B2 => registers_25_21_port, ZN => n4027);
   U2760 : OAI221_X1 port map( B1 => n2169, B2 => n5643, C1 => n2504, C2 => 
                           n5473, A => n4008, ZN => n2918);
   U2761 : AOI22_X1 port map( A1 => n5645, A2 => registers_28_22_port, B1 => 
                           n5647, B2 => registers_25_22_port, ZN => n4008);
   U2762 : OAI221_X1 port map( B1 => n2170, B2 => n5642, C1 => n2505, C2 => 
                           n5474, A => n2883, ZN => n2880);
   U2763 : AOI22_X1 port map( A1 => n5644, A2 => registers_28_24_port, B1 => 
                           n5646, B2 => registers_25_24_port, ZN => n2883);
   U2764 : OAI221_X1 port map( B1 => n2171, B2 => n5643, C1 => n2506, C2 => 
                           n5472, A => n2864, ZN => n2861);
   U2765 : AOI22_X1 port map( A1 => n5645, A2 => registers_28_25_port, B1 => 
                           n5647, B2 => registers_25_25_port, ZN => n2864);
   U2766 : OAI221_X1 port map( B1 => n2172, B2 => n5642, C1 => n2507, C2 => 
                           n5473, A => n2826, ZN => n2823);
   U2767 : AOI22_X1 port map( A1 => n5644, A2 => registers_28_27_port, B1 => 
                           n5646, B2 => registers_25_27_port, ZN => n2826);
   U2768 : OAI221_X1 port map( B1 => n2173, B2 => n5643, C1 => n2508, C2 => 
                           n5474, A => n2807, ZN => n2804);
   U2769 : AOI22_X1 port map( A1 => n5645, A2 => registers_28_28_port, B1 => 
                           n5647, B2 => registers_25_28_port, ZN => n2807);
   U2770 : OAI221_X1 port map( B1 => n2174, B2 => n5642, C1 => n2509, C2 => 
                           n5472, A => n2769, ZN => n2766);
   U2771 : AOI22_X1 port map( A1 => n5644, A2 => registers_28_30_port, B1 => 
                           n5646, B2 => registers_25_30_port, ZN => n2769);
   U2772 : OAI221_X1 port map( B1 => n2175, B2 => n5643, C1 => n2510, C2 => 
                           n5473, A => n2727, ZN => n2718);
   U2773 : AOI22_X1 port map( A1 => n5645, A2 => registers_28_31_port, B1 => 
                           n5647, B2 => registers_25_31_port, ZN => n2727);
   U2774 : OAI221_X1 port map( B1 => n2176, B2 => n2725, C1 => n2513, C2 => 
                           n5472, A => n4388, ZN => n4385);
   U2775 : AOI22_X1 port map( A1 => n2728, A2 => registers_28_2_port, B1 => 
                           n2729, B2 => registers_25_2_port, ZN => n4388);
   U2776 : OAI221_X1 port map( B1 => n2177, B2 => n2725, C1 => n2514, C2 => 
                           n5473, A => n4331, ZN => n4328);
   U2777 : AOI22_X1 port map( A1 => n2728, A2 => registers_28_5_port, B1 => 
                           n2729, B2 => registers_25_5_port, ZN => n4331);
   U2778 : OAI221_X1 port map( B1 => n2178, B2 => n2725, C1 => n2515, C2 => 
                           n5474, A => n4274, ZN => n4271);
   U2779 : AOI22_X1 port map( A1 => n2728, A2 => registers_28_8_port, B1 => 
                           n2729, B2 => registers_25_8_port, ZN => n4274);
   U2780 : OAI221_X1 port map( B1 => n2179, B2 => n2725, C1 => n2516, C2 => 
                           n5472, A => n4217, ZN => n4214);
   U2781 : AOI22_X1 port map( A1 => n2728, A2 => registers_28_11_port, B1 => 
                           n2729, B2 => registers_25_11_port, ZN => n4217);
   U2782 : OAI221_X1 port map( B1 => n2184, B2 => n2725, C1 => n2517, C2 => 
                           n5473, A => n4160, ZN => n4157);
   U2783 : AOI22_X1 port map( A1 => n2728, A2 => registers_28_14_port, B1 => 
                           n2729, B2 => registers_25_14_port, ZN => n4160);
   U2784 : OAI221_X1 port map( B1 => n2185, B2 => n2725, C1 => n2518, C2 => 
                           n5474, A => n4103, ZN => n4100);
   U2785 : AOI22_X1 port map( A1 => n2728, A2 => registers_28_17_port, B1 => 
                           n2729, B2 => registers_25_17_port, ZN => n4103);
   U2786 : OAI221_X1 port map( B1 => n2186, B2 => n2725, C1 => n2519, C2 => 
                           n5472, A => n4046, ZN => n4043);
   U2787 : AOI22_X1 port map( A1 => n2728, A2 => registers_28_20_port, B1 => 
                           n2729, B2 => registers_25_20_port, ZN => n4046);
   U2788 : OAI221_X1 port map( B1 => n2187, B2 => n2725, C1 => n2520, C2 => 
                           n5473, A => n2902, ZN => n2899);
   U2789 : AOI22_X1 port map( A1 => n2728, A2 => registers_28_23_port, B1 => 
                           n2729, B2 => registers_25_23_port, ZN => n2902);
   U2790 : OAI221_X1 port map( B1 => n2188, B2 => n2725, C1 => n2521, C2 => 
                           n5474, A => n2845, ZN => n2842);
   U2791 : AOI22_X1 port map( A1 => n2728, A2 => registers_28_26_port, B1 => 
                           n2729, B2 => registers_25_26_port, ZN => n2845);
   U2792 : OAI221_X1 port map( B1 => n2189, B2 => n2725, C1 => n2522, C2 => 
                           n5472, A => n2788, ZN => n2785);
   U2793 : AOI22_X1 port map( A1 => n2728, A2 => registers_28_29_port, B1 => 
                           n2729, B2 => registers_25_29_port, ZN => n2788);
   U2794 : OAI221_X1 port map( B1 => n2225, B2 => n5649, C1 => n2153, C2 => 
                           n5476, A => n4457, ZN => n4456);
   U2795 : AOI22_X1 port map( A1 => n5655, A2 => registers_19_0_port, B1 => 
                           n5658, B2 => registers_22_0_port, ZN => n4457);
   U2796 : OAI221_X1 port map( B1 => n2190, B2 => n5650, C1 => n2051, C2 => 
                           n5477, A => n4406, ZN => n4405);
   U2797 : AOI22_X1 port map( A1 => n5656, A2 => registers_19_1_port, B1 => 
                           n5659, B2 => registers_22_1_port, ZN => n4406);
   U2798 : OAI221_X1 port map( B1 => n2191, B2 => n5649, C1 => n2052, C2 => 
                           n5475, A => n4387, ZN => n4386);
   U2799 : AOI22_X1 port map( A1 => n2723, A2 => registers_19_2_port, B1 => 
                           n5657, B2 => registers_22_2_port, ZN => n4387);
   U2800 : OAI221_X1 port map( B1 => n2192, B2 => n5650, C1 => n2053, C2 => 
                           n5475, A => n4368, ZN => n4367);
   U2801 : AOI22_X1 port map( A1 => n5655, A2 => registers_19_3_port, B1 => 
                           n5657, B2 => registers_22_3_port, ZN => n4368);
   U2802 : OAI221_X1 port map( B1 => n2193, B2 => n5651, C1 => n2054, C2 => 
                           n5476, A => n4349, ZN => n4348);
   U2803 : AOI22_X1 port map( A1 => n5656, A2 => registers_19_4_port, B1 => 
                           n5658, B2 => registers_22_4_port, ZN => n4349);
   U2804 : OAI221_X1 port map( B1 => n2194, B2 => n5652, C1 => n2055, C2 => 
                           n5476, A => n4330, ZN => n4329);
   U2805 : AOI22_X1 port map( A1 => n2723, A2 => registers_19_5_port, B1 => 
                           n5658, B2 => registers_22_5_port, ZN => n4330);
   U2806 : OAI221_X1 port map( B1 => n2195, B2 => n5651, C1 => n2056, C2 => 
                           n5477, A => n4311, ZN => n4310);
   U2807 : AOI22_X1 port map( A1 => n5655, A2 => registers_19_6_port, B1 => 
                           n5659, B2 => registers_22_6_port, ZN => n4311);
   U2808 : OAI221_X1 port map( B1 => n2196, B2 => n5652, C1 => n2057, C2 => 
                           n5475, A => n4292, ZN => n4291);
   U2809 : AOI22_X1 port map( A1 => n5656, A2 => registers_19_7_port, B1 => 
                           n5657, B2 => registers_22_7_port, ZN => n4292);
   U2810 : OAI221_X1 port map( B1 => n2197, B2 => n5653, C1 => n2058, C2 => 
                           n5477, A => n4273, ZN => n4272);
   U2811 : AOI22_X1 port map( A1 => n2723, A2 => registers_19_8_port, B1 => 
                           n5659, B2 => registers_22_8_port, ZN => n4273);
   U2812 : OAI221_X1 port map( B1 => n2198, B2 => n5654, C1 => n2059, C2 => 
                           n5476, A => n4254, ZN => n4253);
   U2813 : AOI22_X1 port map( A1 => n5655, A2 => registers_19_9_port, B1 => 
                           n5658, B2 => registers_22_9_port, ZN => n4254);
   U2814 : OAI221_X1 port map( B1 => n2199, B2 => n5649, C1 => n2060, C2 => 
                           n5477, A => n4235, ZN => n4234);
   U2815 : AOI22_X1 port map( A1 => n5656, A2 => registers_19_10_port, B1 => 
                           n5659, B2 => registers_22_10_port, ZN => n4235);
   U2816 : OAI221_X1 port map( B1 => n2200, B2 => n5650, C1 => n2061, C2 => 
                           n5475, A => n4216, ZN => n4215);
   U2817 : AOI22_X1 port map( A1 => n2723, A2 => registers_19_11_port, B1 => 
                           n5657, B2 => registers_22_11_port, ZN => n4216);
   U2818 : OAI221_X1 port map( B1 => n2201, B2 => n5653, C1 => n2062, C2 => 
                           n5475, A => n4197, ZN => n4196);
   U2819 : AOI22_X1 port map( A1 => n5655, A2 => registers_19_12_port, B1 => 
                           n5657, B2 => registers_22_12_port, ZN => n4197);
   U2820 : OAI221_X1 port map( B1 => n2202, B2 => n5654, C1 => n2063, C2 => 
                           n5476, A => n4178, ZN => n4177);
   U2821 : AOI22_X1 port map( A1 => n5656, A2 => registers_19_13_port, B1 => 
                           n5658, B2 => registers_22_13_port, ZN => n4178);
   U2822 : OAI221_X1 port map( B1 => n2203, B2 => n5651, C1 => n2064, C2 => 
                           n5476, A => n4159, ZN => n4158);
   U2823 : AOI22_X1 port map( A1 => n2723, A2 => registers_19_14_port, B1 => 
                           n5658, B2 => registers_22_14_port, ZN => n4159);
   U2824 : OAI221_X1 port map( B1 => n2204, B2 => n5652, C1 => n2065, C2 => 
                           n5477, A => n4140, ZN => n4139);
   U2825 : AOI22_X1 port map( A1 => n5655, A2 => registers_19_15_port, B1 => 
                           n5659, B2 => registers_22_15_port, ZN => n4140);
   U2826 : OAI221_X1 port map( B1 => n2205, B2 => n5653, C1 => n2066, C2 => 
                           n5475, A => n4121, ZN => n4120);
   U2827 : AOI22_X1 port map( A1 => n5656, A2 => registers_19_16_port, B1 => 
                           n5657, B2 => registers_22_16_port, ZN => n4121);
   U2828 : OAI221_X1 port map( B1 => n2206, B2 => n5654, C1 => n2067, C2 => 
                           n5477, A => n4102, ZN => n4101);
   U2829 : AOI22_X1 port map( A1 => n2723, A2 => registers_19_17_port, B1 => 
                           n5659, B2 => registers_22_17_port, ZN => n4102);
   U2830 : OAI221_X1 port map( B1 => n2207, B2 => n5649, C1 => n2068, C2 => 
                           n5476, A => n4083, ZN => n4082);
   U2831 : AOI22_X1 port map( A1 => n5655, A2 => registers_19_18_port, B1 => 
                           n5658, B2 => registers_22_18_port, ZN => n4083);
   U2832 : OAI221_X1 port map( B1 => n2208, B2 => n5650, C1 => n2069, C2 => 
                           n5477, A => n4064, ZN => n4063);
   U2833 : AOI22_X1 port map( A1 => n5656, A2 => registers_19_19_port, B1 => 
                           n5659, B2 => registers_22_19_port, ZN => n4064);
   U2834 : OAI221_X1 port map( B1 => n2209, B2 => n5649, C1 => n2070, C2 => 
                           n5475, A => n4045, ZN => n4044);
   U2835 : AOI22_X1 port map( A1 => n2723, A2 => registers_19_20_port, B1 => 
                           n5657, B2 => registers_22_20_port, ZN => n4045);
   U2836 : OAI221_X1 port map( B1 => n2210, B2 => n5650, C1 => n2071, C2 => 
                           n5475, A => n4026, ZN => n4025);
   U2837 : AOI22_X1 port map( A1 => n5655, A2 => registers_19_21_port, B1 => 
                           n5657, B2 => registers_22_21_port, ZN => n4026);
   U2838 : OAI221_X1 port map( B1 => n2211, B2 => n5651, C1 => n2072, C2 => 
                           n5476, A => n4007, ZN => n2950);
   U2839 : AOI22_X1 port map( A1 => n5656, A2 => registers_19_22_port, B1 => 
                           n5658, B2 => registers_22_22_port, ZN => n4007);
   U2840 : OAI221_X1 port map( B1 => n2212, B2 => n5652, C1 => n2073, C2 => 
                           n5476, A => n2901, ZN => n2900);
   U2841 : AOI22_X1 port map( A1 => n2723, A2 => registers_19_23_port, B1 => 
                           n5658, B2 => registers_22_23_port, ZN => n2901);
   U2842 : OAI221_X1 port map( B1 => n2213, B2 => n5651, C1 => n2074, C2 => 
                           n5477, A => n2882, ZN => n2881);
   U2843 : AOI22_X1 port map( A1 => n5655, A2 => registers_19_24_port, B1 => 
                           n5659, B2 => registers_22_24_port, ZN => n2882);
   U2844 : OAI221_X1 port map( B1 => n2214, B2 => n5652, C1 => n2075, C2 => 
                           n5475, A => n2863, ZN => n2862);
   U2845 : AOI22_X1 port map( A1 => n5656, A2 => registers_19_25_port, B1 => 
                           n5657, B2 => registers_22_25_port, ZN => n2863);
   U2846 : OAI221_X1 port map( B1 => n2215, B2 => n5653, C1 => n2076, C2 => 
                           n5477, A => n2844, ZN => n2843);
   U2847 : AOI22_X1 port map( A1 => n2723, A2 => registers_19_26_port, B1 => 
                           n5659, B2 => registers_22_26_port, ZN => n2844);
   U2848 : OAI221_X1 port map( B1 => n2216, B2 => n5654, C1 => n2077, C2 => 
                           n5476, A => n2825, ZN => n2824);
   U2849 : AOI22_X1 port map( A1 => n5655, A2 => registers_19_27_port, B1 => 
                           n5658, B2 => registers_22_27_port, ZN => n2825);
   U2850 : OAI221_X1 port map( B1 => n2219, B2 => n5649, C1 => n2080, C2 => 
                           n5477, A => n2806, ZN => n2805);
   U2851 : AOI22_X1 port map( A1 => n5656, A2 => registers_19_28_port, B1 => 
                           n5659, B2 => registers_22_28_port, ZN => n2806);
   U2852 : OAI221_X1 port map( B1 => n2220, B2 => n5650, C1 => n2112, C2 => 
                           n5475, A => n2787, ZN => n2786);
   U2853 : AOI22_X1 port map( A1 => n2723, A2 => registers_19_29_port, B1 => 
                           n5657, B2 => registers_22_29_port, ZN => n2787);
   U2854 : OAI221_X1 port map( B1 => n2221, B2 => n5653, C1 => n2114, C2 => 
                           n5475, A => n2768, ZN => n2767);
   U2855 : AOI22_X1 port map( A1 => n5655, A2 => registers_19_30_port, B1 => 
                           n5657, B2 => registers_22_30_port, ZN => n2768);
   U2856 : OAI221_X1 port map( B1 => n2222, B2 => n5654, C1 => n2115, C2 => 
                           n5476, A => n2722, ZN => n2719);
   U2857 : AOI22_X1 port map( A1 => n5656, A2 => registers_19_31_port, B1 => 
                           n5658, B2 => registers_22_31_port, ZN => n2722);
   U2858 : OAI221_X1 port map( B1 => n5154, B2 => n5636, C1 => n2258, C2 => 
                           n5471, A => n4408, ZN => n4403);
   U2859 : AOI22_X1 port map( A1 => n5639, A2 => registers_2_1_port, B1 => 
                           n5641, B2 => registers_29_1_port, ZN => n4408);
   U2860 : OAI221_X1 port map( B1 => n5155, B2 => n5632, C1 => n2259, C2 => 
                           n5469, A => n4389, ZN => n4384);
   U2861 : AOI22_X1 port map( A1 => n5637, A2 => registers_2_2_port, B1 => 
                           n2734, B2 => registers_29_2_port, ZN => n4389);
   U2862 : OAI221_X1 port map( B1 => n5156, B2 => n5635, C1 => n2260, C2 => 
                           n5469, A => n4370, ZN => n4365);
   U2863 : AOI22_X1 port map( A1 => n5637, A2 => registers_2_3_port, B1 => 
                           n5640, B2 => registers_29_3_port, ZN => n4370);
   U2864 : OAI221_X1 port map( B1 => n5157, B2 => n5630, C1 => n2261, C2 => 
                           n5470, A => n4351, ZN => n4346);
   U2865 : AOI22_X1 port map( A1 => n5638, A2 => registers_2_4_port, B1 => 
                           n5641, B2 => registers_29_4_port, ZN => n4351);
   U2866 : OAI221_X1 port map( B1 => n5158, B2 => n5632, C1 => n2262, C2 => 
                           n5470, A => n4332, ZN => n4327);
   U2867 : AOI22_X1 port map( A1 => n5638, A2 => registers_2_5_port, B1 => 
                           n2734, B2 => registers_29_5_port, ZN => n4332);
   U2868 : OAI221_X1 port map( B1 => n5159, B2 => n5631, C1 => n2263, C2 => 
                           n5471, A => n4313, ZN => n4308);
   U2869 : AOI22_X1 port map( A1 => n5639, A2 => registers_2_6_port, B1 => 
                           n5640, B2 => registers_29_6_port, ZN => n4313);
   U2870 : OAI221_X1 port map( B1 => n5160, B2 => n5632, C1 => n2264, C2 => 
                           n5469, A => n4294, ZN => n4289);
   U2871 : AOI22_X1 port map( A1 => n5637, A2 => registers_2_7_port, B1 => 
                           n5641, B2 => registers_29_7_port, ZN => n4294);
   U2872 : OAI221_X1 port map( B1 => n5161, B2 => n5631, C1 => n2265, C2 => 
                           n5471, A => n4275, ZN => n4270);
   U2873 : AOI22_X1 port map( A1 => n5639, A2 => registers_2_8_port, B1 => 
                           n2734, B2 => registers_29_8_port, ZN => n4275);
   U2874 : OAI221_X1 port map( B1 => n5162, B2 => n5634, C1 => n2266, C2 => 
                           n5470, A => n4256, ZN => n4251);
   U2875 : AOI22_X1 port map( A1 => n5638, A2 => registers_2_9_port, B1 => 
                           n5640, B2 => registers_29_9_port, ZN => n4256);
   U2876 : OAI221_X1 port map( B1 => n5163, B2 => n5633, C1 => n2267, C2 => 
                           n5471, A => n4237, ZN => n4232);
   U2877 : AOI22_X1 port map( A1 => n5639, A2 => registers_2_10_port, B1 => 
                           n5641, B2 => registers_29_10_port, ZN => n4237);
   U2878 : OAI221_X1 port map( B1 => n5164, B2 => n5634, C1 => n2268, C2 => 
                           n5469, A => n4218, ZN => n4213);
   U2879 : AOI22_X1 port map( A1 => n5637, A2 => registers_2_11_port, B1 => 
                           n2734, B2 => registers_29_11_port, ZN => n4218);
   U2880 : OAI221_X1 port map( B1 => n5165, B2 => n5630, C1 => n2269, C2 => 
                           n5469, A => n4199, ZN => n4194);
   U2881 : AOI22_X1 port map( A1 => n5637, A2 => registers_2_12_port, B1 => 
                           n5640, B2 => registers_29_12_port, ZN => n4199);
   U2882 : OAI221_X1 port map( B1 => n5166, B2 => n5631, C1 => n2270, C2 => 
                           n5470, A => n4180, ZN => n4175);
   U2883 : AOI22_X1 port map( A1 => n5638, A2 => registers_2_13_port, B1 => 
                           n5641, B2 => registers_29_13_port, ZN => n4180);
   U2884 : OAI221_X1 port map( B1 => n5167, B2 => n5631, C1 => n2271, C2 => 
                           n5470, A => n4161, ZN => n4156);
   U2885 : AOI22_X1 port map( A1 => n5638, A2 => registers_2_14_port, B1 => 
                           n2734, B2 => registers_29_14_port, ZN => n4161);
   U2886 : OAI221_X1 port map( B1 => n5168, B2 => n5632, C1 => n2272, C2 => 
                           n5471, A => n4142, ZN => n4137);
   U2887 : AOI22_X1 port map( A1 => n5639, A2 => registers_2_15_port, B1 => 
                           n5640, B2 => registers_29_15_port, ZN => n4142);
   U2888 : OAI221_X1 port map( B1 => n5169, B2 => n5632, C1 => n2273, C2 => 
                           n5469, A => n4123, ZN => n4118);
   U2889 : AOI22_X1 port map( A1 => n5637, A2 => registers_2_16_port, B1 => 
                           n5641, B2 => registers_29_16_port, ZN => n4123);
   U2890 : OAI221_X1 port map( B1 => n5170, B2 => n5636, C1 => n2274, C2 => 
                           n5471, A => n4104, ZN => n4099);
   U2891 : AOI22_X1 port map( A1 => n5639, A2 => registers_2_17_port, B1 => 
                           n2734, B2 => registers_29_17_port, ZN => n4104);
   U2892 : OAI221_X1 port map( B1 => n5171, B2 => n5633, C1 => n2275, C2 => 
                           n5470, A => n4085, ZN => n4080);
   U2893 : AOI22_X1 port map( A1 => n5638, A2 => registers_2_18_port, B1 => 
                           n5640, B2 => registers_29_18_port, ZN => n4085);
   U2894 : OAI221_X1 port map( B1 => n5172, B2 => n5634, C1 => n2276, C2 => 
                           n5471, A => n4066, ZN => n4061);
   U2895 : AOI22_X1 port map( A1 => n5639, A2 => registers_2_19_port, B1 => 
                           n5641, B2 => registers_29_19_port, ZN => n4066);
   U2896 : OAI221_X1 port map( B1 => n5173, B2 => n5633, C1 => n2277, C2 => 
                           n5469, A => n4047, ZN => n4042);
   U2897 : AOI22_X1 port map( A1 => n5637, A2 => registers_2_20_port, B1 => 
                           n2734, B2 => registers_29_20_port, ZN => n4047);
   U2898 : OAI221_X1 port map( B1 => n5174, B2 => n5634, C1 => n2278, C2 => 
                           n5469, A => n4028, ZN => n4023);
   U2899 : AOI22_X1 port map( A1 => n5637, A2 => registers_2_21_port, B1 => 
                           n5640, B2 => registers_29_21_port, ZN => n4028);
   U2900 : OAI221_X1 port map( B1 => n5175, B2 => n5636, C1 => n2279, C2 => 
                           n5470, A => n4009, ZN => n2917);
   U2901 : AOI22_X1 port map( A1 => n5638, A2 => registers_2_22_port, B1 => 
                           n5641, B2 => registers_29_22_port, ZN => n4009);
   U2902 : OAI221_X1 port map( B1 => n5176, B2 => n5635, C1 => n2280, C2 => 
                           n5470, A => n2903, ZN => n2898);
   U2903 : AOI22_X1 port map( A1 => n5638, A2 => registers_2_23_port, B1 => 
                           n2734, B2 => registers_29_23_port, ZN => n2903);
   U2904 : OAI221_X1 port map( B1 => n5177, B2 => n5635, C1 => n2281, C2 => 
                           n5471, A => n2884, ZN => n2879);
   U2905 : AOI22_X1 port map( A1 => n5639, A2 => registers_2_24_port, B1 => 
                           n5640, B2 => registers_29_24_port, ZN => n2884);
   U2906 : OAI221_X1 port map( B1 => n5178, B2 => n5636, C1 => n2282, C2 => 
                           n5469, A => n2865, ZN => n2860);
   U2907 : AOI22_X1 port map( A1 => n5637, A2 => registers_2_25_port, B1 => 
                           n5641, B2 => registers_29_25_port, ZN => n2865);
   U2908 : OAI221_X1 port map( B1 => n5179, B2 => n5635, C1 => n2119, C2 => 
                           n5471, A => n2846, ZN => n2841);
   U2909 : AOI22_X1 port map( A1 => n5639, A2 => registers_2_26_port, B1 => 
                           n2734, B2 => registers_29_26_port, ZN => n2846);
   U2910 : OAI221_X1 port map( B1 => n2388, B2 => n5636, C1 => n2120, C2 => 
                           n5470, A => n2827, ZN => n2822);
   U2911 : AOI22_X1 port map( A1 => n5638, A2 => registers_2_27_port, B1 => 
                           n5640, B2 => registers_29_27_port, ZN => n2827);
   U2912 : OAI221_X1 port map( B1 => n5180, B2 => n5631, C1 => n2283, C2 => 
                           n5471, A => n2808, ZN => n2803);
   U2913 : AOI22_X1 port map( A1 => n5639, A2 => registers_2_28_port, B1 => 
                           n5641, B2 => registers_29_28_port, ZN => n2808);
   U2914 : OAI221_X1 port map( B1 => n5181, B2 => n5634, C1 => n2284, C2 => 
                           n5469, A => n2789, ZN => n2784);
   U2915 : AOI22_X1 port map( A1 => n5637, A2 => registers_2_29_port, B1 => 
                           n2734, B2 => registers_29_29_port, ZN => n2789);
   U2916 : OAI221_X1 port map( B1 => n5182, B2 => n5630, C1 => n2285, C2 => 
                           n5469, A => n2770, ZN => n2765);
   U2917 : AOI22_X1 port map( A1 => n5637, A2 => registers_2_30_port, B1 => 
                           n5640, B2 => registers_29_30_port, ZN => n2770);
   U2918 : OAI221_X1 port map( B1 => n5183, B2 => n5633, C1 => n2287, C2 => 
                           n5470, A => n2732, ZN => n2717);
   U2919 : AOI22_X1 port map( A1 => n5638, A2 => registers_2_31_port, B1 => 
                           n5641, B2 => registers_29_31_port, ZN => n2732);
   U2920 : AOI22_X1 port map( A1 => n5638, A2 => registers_2_0_port, B1 => 
                           n5640, B2 => registers_29_0_port, ZN => n4462);
   U2921 : AOI22_X1 port map( A1 => n5614, A2 => registers_14_0_port, B1 => 
                           n5623, B2 => registers_11_0_port, ZN => n4463);
   U2922 : AOI22_X1 port map( A1 => n5619, A2 => registers_14_1_port, B1 => 
                           n5627, B2 => registers_11_1_port, ZN => n4409);
   U2923 : AOI22_X1 port map( A1 => n5620, A2 => registers_14_2_port, B1 => 
                           n5623, B2 => registers_11_2_port, ZN => n4390);
   U2924 : AOI22_X1 port map( A1 => n5615, A2 => registers_14_3_port, B1 => 
                           n5624, B2 => registers_11_3_port, ZN => n4371);
   U2925 : AOI22_X1 port map( A1 => n5615, A2 => registers_14_4_port, B1 => 
                           n5624, B2 => registers_11_4_port, ZN => n4352);
   U2926 : AOI22_X1 port map( A1 => n5618, A2 => registers_14_5_port, B1 => 
                           n5624, B2 => registers_11_5_port, ZN => n4333);
   U2927 : AOI22_X1 port map( A1 => n5616, A2 => registers_14_6_port, B1 => 
                           n5625, B2 => registers_11_6_port, ZN => n4314);
   U2928 : AOI22_X1 port map( A1 => n5616, A2 => registers_14_7_port, B1 => 
                           n5623, B2 => registers_11_7_port, ZN => n4295);
   U2929 : AOI22_X1 port map( A1 => n5616, A2 => registers_14_8_port, B1 => 
                           n5623, B2 => registers_11_8_port, ZN => n4276);
   U2930 : AOI22_X1 port map( A1 => n5618, A2 => registers_14_9_port, B1 => 
                           n5626, B2 => registers_11_9_port, ZN => n4257);
   U2931 : AOI22_X1 port map( A1 => n5617, A2 => registers_14_10_port, B1 => 
                           n5625, B2 => registers_11_10_port, ZN => n4238);
   U2932 : AOI22_X1 port map( A1 => n5618, A2 => registers_14_11_port, B1 => 
                           n5626, B2 => registers_11_11_port, ZN => n4219);
   U2933 : AOI22_X1 port map( A1 => n5619, A2 => registers_14_12_port, B1 => 
                           n5627, B2 => registers_11_12_port, ZN => n4200);
   U2934 : AOI22_X1 port map( A1 => n5619, A2 => registers_14_13_port, B1 => 
                           n5627, B2 => registers_11_13_port, ZN => n4181);
   U2935 : AOI22_X1 port map( A1 => n5617, A2 => registers_14_14_port, B1 => 
                           n5625, B2 => registers_11_14_port, ZN => n4162);
   U2936 : AOI22_X1 port map( A1 => n5618, A2 => registers_14_15_port, B1 => 
                           n5626, B2 => registers_11_15_port, ZN => n4143);
   U2937 : AOI22_X1 port map( A1 => n5619, A2 => registers_14_16_port, B1 => 
                           n5627, B2 => registers_11_16_port, ZN => n4124);
   U2938 : AOI22_X1 port map( A1 => n5619, A2 => registers_14_17_port, B1 => 
                           n5627, B2 => registers_11_17_port, ZN => n4105);
   U2939 : AOI22_X1 port map( A1 => n5620, A2 => registers_14_18_port, B1 => 
                           n5628, B2 => registers_11_18_port, ZN => n4086);
   U2940 : AOI22_X1 port map( A1 => n5620, A2 => registers_14_19_port, B1 => 
                           n5628, B2 => registers_11_19_port, ZN => n4067);
   U2941 : AOI22_X1 port map( A1 => n5620, A2 => registers_14_20_port, B1 => 
                           n5628, B2 => registers_11_20_port, ZN => n4048);
   U2942 : AOI22_X1 port map( A1 => n5620, A2 => registers_14_21_port, B1 => 
                           n5628, B2 => registers_11_21_port, ZN => n4029);
   U2943 : AOI22_X1 port map( A1 => n5614, A2 => registers_14_22_port, B1 => 
                           n5623, B2 => registers_11_22_port, ZN => n4010);
   U2944 : AOI22_X1 port map( A1 => n5614, A2 => registers_14_23_port, B1 => 
                           n5627, B2 => registers_11_23_port, ZN => n2904);
   U2945 : AOI22_X1 port map( A1 => n5619, A2 => registers_14_24_port, B1 => 
                           n5628, B2 => registers_11_24_port, ZN => n2885);
   U2946 : AOI22_X1 port map( A1 => n5615, A2 => registers_14_25_port, B1 => 
                           n5624, B2 => registers_11_25_port, ZN => n2866);
   U2947 : AOI22_X1 port map( A1 => n5615, A2 => registers_14_26_port, B1 => 
                           n5626, B2 => registers_11_26_port, ZN => n2847);
   U2948 : AOI22_X1 port map( A1 => n5618, A2 => registers_14_27_port, B1 => 
                           n5626, B2 => registers_11_27_port, ZN => n2828);
   U2949 : AOI22_X1 port map( A1 => n5616, A2 => registers_14_28_port, B1 => 
                           n5625, B2 => registers_11_28_port, ZN => n2809);
   U2950 : AOI22_X1 port map( A1 => n5614, A2 => registers_14_29_port, B1 => 
                           n5626, B2 => registers_11_29_port, ZN => n2790);
   U2951 : AOI22_X1 port map( A1 => n5617, A2 => registers_14_30_port, B1 => 
                           n5628, B2 => registers_11_30_port, ZN => n2771);
   U2952 : AOI22_X1 port map( A1 => n5617, A2 => registers_14_31_port, B1 => 
                           n5625, B2 => registers_11_31_port, ZN => n2737);
   U2953 : INV_X1 port map( A => rd2_addr(1), ZN => n4458);
   U2954 : INV_X1 port map( A => rd2_addr(2), ZN => n4441);
   U2955 : INV_X1 port map( A => rd1_addr(2), ZN => n5095);
   U2956 : INV_X1 port map( A => rd2_addr(4), ZN => n4459);
   U2957 : INV_X1 port map( A => rd1_addr(4), ZN => n5096);
   U2958 : AND3_X1 port map( A1 => n6156, A2 => en, A3 => rd1_en, ZN => n5490);
   U2959 : AND3_X1 port map( A1 => n6156, A2 => en, A3 => rd1_en, ZN => n4476);
   U2960 : AND3_X1 port map( A1 => n6156, A2 => en, A3 => rd1_en, ZN => n5489);
   U2961 : NOR3_X1 port map( A1 => n4461, A2 => rd2_addr(0), A3 => n4459, ZN =>
                           n4442);
   U2962 : NOR3_X1 port map( A1 => n5096, A2 => rd1_addr(0), A3 => n5097, ZN =>
                           n5079);
   U2963 : NOR3_X1 port map( A1 => n4434, A2 => rd2_addr(4), A3 => n4461, ZN =>
                           n4426);
   U2964 : AND3_X1 port map( A1 => rd2_addr(2), A2 => n4458, A3 => n4442, ZN =>
                           n5644);
   U2965 : AND3_X1 port map( A1 => rd2_addr(2), A2 => n4458, A3 => n4442, ZN =>
                           n5645);
   U2966 : AND3_X1 port map( A1 => rd2_addr(2), A2 => n4458, A3 => n4438, ZN =>
                           n5640);
   U2967 : AND3_X1 port map( A1 => rd2_addr(2), A2 => n4458, A3 => n4438, ZN =>
                           n5641);
   U2968 : AND3_X1 port map( A1 => rd2_addr(2), A2 => n4458, A3 => n4442, ZN =>
                           n2728);
   U2969 : AND3_X1 port map( A1 => rd2_addr(2), A2 => n4458, A3 => n4438, ZN =>
                           n2734);
   U2970 : INV_X1 port map( A => rd1_addr(1), ZN => n5090);
   U2971 : NOR2_X1 port map( A1 => rd2_addr(3), A2 => rd2_addr(4), ZN => n4433)
                           ;
   U2972 : NOR2_X1 port map( A1 => rd1_addr(3), A2 => rd1_addr(4), ZN => n5086)
                           ;
   U2973 : INV_X1 port map( A => rd2_addr(0), ZN => n4434);
   U2974 : INV_X1 port map( A => rd1_addr(0), ZN => n5087);
   U2975 : AND2_X1 port map( A1 => n4433, A2 => rd2_addr(0), ZN => n4435);
   U2976 : AND2_X1 port map( A1 => n5086, A2 => rd1_addr(0), ZN => n5085);
   U2977 : INV_X1 port map( A => rd1_addr(3), ZN => n5097);
   U2978 : INV_X1 port map( A => rd2_addr(3), ZN => n4461);
   U2979 : INV_X1 port map( A => wr_en, ZN => n2182);
   U2980 : NAND3_X1 port map( A1 => n5081, A2 => n5504, A3 => n5078, ZN => 
                           n5438);
   U2981 : NAND3_X1 port map( A1 => n5081, A2 => n5504, A3 => n5078, ZN => 
                           n5439);
   U2982 : NAND3_X1 port map( A1 => n5078, A2 => n5506, A3 => n5088, ZN => 
                           n5443);
   U2983 : NAND3_X1 port map( A1 => n5078, A2 => n5506, A3 => n5088, ZN => 
                           n5444);
   U2984 : NAND3_X1 port map( A1 => n5081, A2 => n5504, A3 => n5067, ZN => 
                           n5448);
   U2985 : NAND3_X1 port map( A1 => n5081, A2 => n5504, A3 => n5067, ZN => 
                           n5449);
   U2986 : NAND3_X1 port map( A1 => n5078, A2 => n5505, A3 => n5069, ZN => 
                           n5456);
   U2987 : NAND3_X1 port map( A1 => n5078, A2 => n5505, A3 => n5069, ZN => 
                           n5457);
   U2988 : NAND3_X1 port map( A1 => n5067, A2 => n5505, A3 => n5079, ZN => 
                           n5461);
   U2989 : NAND3_X1 port map( A1 => n5067, A2 => n5505, A3 => n5079, ZN => 
                           n5462);
   U2990 : NAND3_X1 port map( A1 => n4433, A2 => n4434, A3 => n4425, ZN => 
                           n5484);
   U2991 : NAND3_X1 port map( A1 => n4433, A2 => n4434, A3 => n4425, ZN => 
                           n5485);
   U2992 : INV_X1 port map( A => n4509, ZN => n5515);
   U2993 : INV_X1 port map( A => n4509, ZN => n5516);
   U2994 : INV_X1 port map( A => n5515, ZN => n5517);
   U2995 : INV_X1 port map( A => n5515, ZN => n5518);
   U2996 : INV_X1 port map( A => n5516, ZN => n5519);
   U2997 : INV_X1 port map( A => n5515, ZN => n5520);
   U2998 : INV_X1 port map( A => n5516, ZN => n5521);
   U2999 : INV_X1 port map( A => n5516, ZN => n5522);
   U3000 : INV_X1 port map( A => n5543, ZN => n5544);
   U3001 : INV_X1 port map( A => n5543, ZN => n5545);
   U3002 : INV_X1 port map( A => n5543, ZN => n5546);
   U3003 : INV_X1 port map( A => n5543, ZN => n5547);
   U3004 : INV_X1 port map( A => n5543, ZN => n5548);
   U3005 : INV_X1 port map( A => n5543, ZN => n5549);
   U3006 : INV_X1 port map( A => n5543, ZN => n5550);
   U3007 : INV_X1 port map( A => n4494, ZN => n5553);
   U3008 : INV_X1 port map( A => n4494, ZN => n5554);
   U3009 : INV_X1 port map( A => n5553, ZN => n5555);
   U3010 : INV_X1 port map( A => n5553, ZN => n5556);
   U3011 : INV_X1 port map( A => n5554, ZN => n5557);
   U3012 : INV_X1 port map( A => n5553, ZN => n5558);
   U3013 : INV_X1 port map( A => n5554, ZN => n5559);
   U3014 : INV_X1 port map( A => n5554, ZN => n5560);
   U3015 : INV_X1 port map( A => n5598, ZN => n5599);
   U3016 : INV_X1 port map( A => n5598, ZN => n5600);
   U3017 : INV_X1 port map( A => n5598, ZN => n5601);
   U3018 : INV_X1 port map( A => n5598, ZN => n5602);
   U3019 : INV_X1 port map( A => n5598, ZN => n5603);
   U3020 : INV_X1 port map( A => n5598, ZN => n5604);
   U3021 : INV_X1 port map( A => n5598, ZN => n5605);
   U3022 : INV_X1 port map( A => n2738, ZN => n5613);
   U3023 : INV_X1 port map( A => n5613, ZN => n5614);
   U3024 : INV_X1 port map( A => n5613, ZN => n5615);
   U3025 : INV_X1 port map( A => n5613, ZN => n5616);
   U3026 : INV_X1 port map( A => n5613, ZN => n5617);
   U3027 : INV_X1 port map( A => n5613, ZN => n5618);
   U3028 : INV_X1 port map( A => n5613, ZN => n5619);
   U3029 : INV_X1 port map( A => n5613, ZN => n5620);
   U3030 : INV_X1 port map( A => n2739, ZN => n5621);
   U3031 : INV_X1 port map( A => n2739, ZN => n5622);
   U3032 : INV_X1 port map( A => n5621, ZN => n5623);
   U3033 : INV_X1 port map( A => n5621, ZN => n5624);
   U3034 : INV_X1 port map( A => n5621, ZN => n5625);
   U3035 : INV_X1 port map( A => n5622, ZN => n5626);
   U3036 : INV_X1 port map( A => n5622, ZN => n5627);
   U3037 : INV_X1 port map( A => n5622, ZN => n5628);
   U3038 : INV_X1 port map( A => n5629, ZN => n5630);
   U3039 : INV_X1 port map( A => n5629, ZN => n5631);
   U3040 : INV_X1 port map( A => n5629, ZN => n5632);
   U3041 : INV_X1 port map( A => n5629, ZN => n5633);
   U3042 : INV_X1 port map( A => n5629, ZN => n5634);
   U3043 : INV_X1 port map( A => n5629, ZN => n5635);
   U3044 : INV_X1 port map( A => n5629, ZN => n5636);
   U3045 : INV_X1 port map( A => n5668, ZN => n5670);
   U3046 : INV_X1 port map( A => n5668, ZN => n5671);
   U3047 : INV_X1 port map( A => n5669, ZN => n5672);
   U3048 : INV_X1 port map( A => n5668, ZN => n5673);
   U3049 : INV_X1 port map( A => n5668, ZN => n5674);
   U3050 : INV_X1 port map( A => n5669, ZN => n5675);
   U3051 : INV_X1 port map( A => n5669, ZN => n5676);
   U3052 : INV_X1 port map( A => n2703, ZN => n5688);
   U3053 : INV_X1 port map( A => n5688, ZN => n5689);
   U3054 : INV_X1 port map( A => n5688, ZN => n5690);
   U3055 : INV_X1 port map( A => n5688, ZN => n5691);
   U3056 : INV_X1 port map( A => n5688, ZN => n5692);
   U3057 : INV_X1 port map( A => n5688, ZN => n5693);
   U3058 : INV_X1 port map( A => n5688, ZN => n5694);
   U3059 : INV_X1 port map( A => n5688, ZN => n5695);
   U3060 : INV_X1 port map( A => n5700, ZN => n5701);
   U3061 : INV_X1 port map( A => n5699, ZN => n5702);
   U3062 : INV_X1 port map( A => n5699, ZN => n5703);
   U3063 : INV_X1 port map( A => n5700, ZN => n5704);
   U3064 : INV_X1 port map( A => n5700, ZN => n5705);
   U3065 : INV_X1 port map( A => n5700, ZN => n5706);
   U3066 : INV_X1 port map( A => n5700, ZN => n5707);
   U3067 : INV_X1 port map( A => n5709, ZN => n5710);
   U3068 : INV_X1 port map( A => n5708, ZN => n5711);
   U3069 : INV_X1 port map( A => n5708, ZN => n5712);
   U3070 : INV_X1 port map( A => n5709, ZN => n5713);
   U3071 : INV_X1 port map( A => n5709, ZN => n5714);
   U3072 : INV_X1 port map( A => n5709, ZN => n5715);
   U3073 : INV_X1 port map( A => n5709, ZN => n5716);
   U3074 : INV_X1 port map( A => n5718, ZN => n5719);
   U3075 : INV_X1 port map( A => n5717, ZN => n5720);
   U3076 : INV_X1 port map( A => n5717, ZN => n5721);
   U3077 : INV_X1 port map( A => n5718, ZN => n5722);
   U3078 : INV_X1 port map( A => n5718, ZN => n5723);
   U3079 : INV_X1 port map( A => n5718, ZN => n5724);
   U3080 : INV_X1 port map( A => n5718, ZN => n5725);
   U3081 : INV_X1 port map( A => n5727, ZN => n5728);
   U3082 : INV_X1 port map( A => n5727, ZN => n5729);
   U3083 : INV_X1 port map( A => n5726, ZN => n5730);
   U3084 : INV_X1 port map( A => n5726, ZN => n5731);
   U3085 : INV_X1 port map( A => n5727, ZN => n5732);
   U3086 : INV_X1 port map( A => n5727, ZN => n5733);
   U3087 : INV_X1 port map( A => n5727, ZN => n5734);
   U3088 : INV_X1 port map( A => n5735, ZN => n5737);
   U3089 : INV_X1 port map( A => n5735, ZN => n5738);
   U3090 : INV_X1 port map( A => n5735, ZN => n5739);
   U3091 : INV_X1 port map( A => n5735, ZN => n5740);
   U3092 : INV_X1 port map( A => n5735, ZN => n5741);
   U3093 : INV_X1 port map( A => n5735, ZN => n5742);
   U3094 : INV_X1 port map( A => n5736, ZN => n5743);
   U3095 : INV_X1 port map( A => n5745, ZN => n5746);
   U3096 : INV_X1 port map( A => n5744, ZN => n5747);
   U3097 : INV_X1 port map( A => n5744, ZN => n5748);
   U3098 : INV_X1 port map( A => n5745, ZN => n5749);
   U3099 : INV_X1 port map( A => n5745, ZN => n5750);
   U3100 : INV_X1 port map( A => n5745, ZN => n5751);
   U3101 : INV_X1 port map( A => n5745, ZN => n5752);
   U3102 : INV_X1 port map( A => n5754, ZN => n5755);
   U3103 : INV_X1 port map( A => n5753, ZN => n5756);
   U3104 : INV_X1 port map( A => n5753, ZN => n5757);
   U3105 : INV_X1 port map( A => n5754, ZN => n5758);
   U3106 : INV_X1 port map( A => n5754, ZN => n5759);
   U3107 : INV_X1 port map( A => n5754, ZN => n5760);
   U3108 : INV_X1 port map( A => n5754, ZN => n5761);
   U3109 : INV_X1 port map( A => n5763, ZN => n5764);
   U3110 : INV_X1 port map( A => n5763, ZN => n5765);
   U3111 : INV_X1 port map( A => n5762, ZN => n5766);
   U3112 : INV_X1 port map( A => n5762, ZN => n5767);
   U3113 : INV_X1 port map( A => n5763, ZN => n5768);
   U3114 : INV_X1 port map( A => n5763, ZN => n5769);
   U3115 : INV_X1 port map( A => n5763, ZN => n5770);
   U3116 : INV_X1 port map( A => n5772, ZN => n5773);
   U3117 : INV_X1 port map( A => n5771, ZN => n5774);
   U3118 : INV_X1 port map( A => n5771, ZN => n5775);
   U3119 : INV_X1 port map( A => n5772, ZN => n5776);
   U3120 : INV_X1 port map( A => n5772, ZN => n5777);
   U3121 : INV_X1 port map( A => n5772, ZN => n5778);
   U3122 : INV_X1 port map( A => n5772, ZN => n5779);
   U3123 : INV_X1 port map( A => n5781, ZN => n5782);
   U3124 : INV_X1 port map( A => n5780, ZN => n5783);
   U3125 : INV_X1 port map( A => n5780, ZN => n5784);
   U3126 : INV_X1 port map( A => n5781, ZN => n5785);
   U3127 : INV_X1 port map( A => n5781, ZN => n5786);
   U3128 : INV_X1 port map( A => n5781, ZN => n5787);
   U3129 : INV_X1 port map( A => n5781, ZN => n5788);
   U3130 : INV_X1 port map( A => n5790, ZN => n5791);
   U3131 : INV_X1 port map( A => n5789, ZN => n5792);
   U3132 : INV_X1 port map( A => n5789, ZN => n5793);
   U3133 : INV_X1 port map( A => n5790, ZN => n5794);
   U3134 : INV_X1 port map( A => n5790, ZN => n5795);
   U3135 : INV_X1 port map( A => n5790, ZN => n5796);
   U3136 : INV_X1 port map( A => n5790, ZN => n5797);
   U3137 : INV_X1 port map( A => n5799, ZN => n5800);
   U3138 : INV_X1 port map( A => n5799, ZN => n5801);
   U3139 : INV_X1 port map( A => n5798, ZN => n5802);
   U3140 : INV_X1 port map( A => n5798, ZN => n5803);
   U3141 : INV_X1 port map( A => n5799, ZN => n5804);
   U3142 : INV_X1 port map( A => n5799, ZN => n5805);
   U3143 : INV_X1 port map( A => n5799, ZN => n5806);
   U3144 : INV_X1 port map( A => n5807, ZN => n5809);
   U3145 : INV_X1 port map( A => n5807, ZN => n5810);
   U3146 : INV_X1 port map( A => n5807, ZN => n5811);
   U3147 : INV_X1 port map( A => n5807, ZN => n5812);
   U3148 : INV_X1 port map( A => n5807, ZN => n5813);
   U3149 : INV_X1 port map( A => n5807, ZN => n5814);
   U3150 : INV_X1 port map( A => n5808, ZN => n5815);
   U3151 : INV_X1 port map( A => n5816, ZN => n5818);
   U3152 : INV_X1 port map( A => n5816, ZN => n5819);
   U3153 : INV_X1 port map( A => n5816, ZN => n5820);
   U3154 : INV_X1 port map( A => n5816, ZN => n5821);
   U3155 : INV_X1 port map( A => n5816, ZN => n5822);
   U3156 : INV_X1 port map( A => n5816, ZN => n5823);
   U3157 : INV_X1 port map( A => n5817, ZN => n5824);
   U3158 : INV_X1 port map( A => n5826, ZN => n5827);
   U3159 : INV_X1 port map( A => n5825, ZN => n5828);
   U3160 : INV_X1 port map( A => n5825, ZN => n5829);
   U3161 : INV_X1 port map( A => n5826, ZN => n5830);
   U3162 : INV_X1 port map( A => n5826, ZN => n5831);
   U3163 : INV_X1 port map( A => n5826, ZN => n5832);
   U3164 : INV_X1 port map( A => n5826, ZN => n5833);
   U3165 : INV_X1 port map( A => n5834, ZN => n5836);
   U3166 : INV_X1 port map( A => n5834, ZN => n5837);
   U3167 : INV_X1 port map( A => n5834, ZN => n5838);
   U3168 : INV_X1 port map( A => n5835, ZN => n5839);
   U3169 : INV_X1 port map( A => n5835, ZN => n5840);
   U3170 : INV_X1 port map( A => n5835, ZN => n5841);
   U3171 : INV_X1 port map( A => n5835, ZN => n5842);
   U3172 : INV_X1 port map( A => n5843, ZN => n5845);
   U3173 : INV_X1 port map( A => n5843, ZN => n5846);
   U3174 : INV_X1 port map( A => n5843, ZN => n5847);
   U3175 : INV_X1 port map( A => n5843, ZN => n5848);
   U3176 : INV_X1 port map( A => n5843, ZN => n5849);
   U3177 : INV_X1 port map( A => n5843, ZN => n5850);
   U3178 : INV_X1 port map( A => n5844, ZN => n5851);
   U3179 : INV_X1 port map( A => n5853, ZN => n5854);
   U3180 : INV_X1 port map( A => n5853, ZN => n5855);
   U3181 : INV_X1 port map( A => n5853, ZN => n5856);
   U3182 : INV_X1 port map( A => n5852, ZN => n5857);
   U3183 : INV_X1 port map( A => n5852, ZN => n5858);
   U3184 : INV_X1 port map( A => n5853, ZN => n5859);
   U3185 : INV_X1 port map( A => n5853, ZN => n5860);
   U3186 : INV_X1 port map( A => n5861, ZN => n5863);
   U3187 : INV_X1 port map( A => n5861, ZN => n5864);
   U3188 : INV_X1 port map( A => n5861, ZN => n5865);
   U3189 : INV_X1 port map( A => n5861, ZN => n5866);
   U3190 : INV_X1 port map( A => n5861, ZN => n5867);
   U3191 : INV_X1 port map( A => n5861, ZN => n5868);
   U3192 : INV_X1 port map( A => n5862, ZN => n5869);
   U3193 : INV_X1 port map( A => n5871, ZN => n5872);
   U3194 : INV_X1 port map( A => n5870, ZN => n5873);
   U3195 : INV_X1 port map( A => n5870, ZN => n5874);
   U3196 : INV_X1 port map( A => n5871, ZN => n5875);
   U3197 : INV_X1 port map( A => n5871, ZN => n5876);
   U3198 : INV_X1 port map( A => n5871, ZN => n5877);
   U3199 : INV_X1 port map( A => n5871, ZN => n5878);
   U3200 : INV_X1 port map( A => n5879, ZN => n5881);
   U3201 : INV_X1 port map( A => n5879, ZN => n5882);
   U3202 : INV_X1 port map( A => n5879, ZN => n5883);
   U3203 : INV_X1 port map( A => n5879, ZN => n5884);
   U3204 : INV_X1 port map( A => n5879, ZN => n5885);
   U3205 : INV_X1 port map( A => n5880, ZN => n5886);
   U3206 : INV_X1 port map( A => n5880, ZN => n5887);
   U3207 : INV_X1 port map( A => n5889, ZN => n5890);
   U3208 : INV_X1 port map( A => n5888, ZN => n5891);
   U3209 : INV_X1 port map( A => n5888, ZN => n5892);
   U3210 : INV_X1 port map( A => n5889, ZN => n5893);
   U3211 : INV_X1 port map( A => n5889, ZN => n5894);
   U3212 : INV_X1 port map( A => n5889, ZN => n5895);
   U3213 : INV_X1 port map( A => n5889, ZN => n5896);
   U3214 : INV_X1 port map( A => n5897, ZN => n5899);
   U3215 : INV_X1 port map( A => n5897, ZN => n5900);
   U3216 : INV_X1 port map( A => n5897, ZN => n5901);
   U3217 : INV_X1 port map( A => n5898, ZN => n5902);
   U3218 : INV_X1 port map( A => n5898, ZN => n5903);
   U3219 : INV_X1 port map( A => n5897, ZN => n5904);
   U3220 : INV_X1 port map( A => n5897, ZN => n5905);
   U3221 : INV_X1 port map( A => n5906, ZN => n5908);
   U3222 : INV_X1 port map( A => n5906, ZN => n5909);
   U3223 : INV_X1 port map( A => n5906, ZN => n5910);
   U3224 : INV_X1 port map( A => n5906, ZN => n5911);
   U3225 : INV_X1 port map( A => n5906, ZN => n5912);
   U3226 : INV_X1 port map( A => n5907, ZN => n5913);
   U3227 : INV_X1 port map( A => n5907, ZN => n5914);
   U3228 : INV_X1 port map( A => n5915, ZN => n5917);
   U3229 : INV_X1 port map( A => n5915, ZN => n5918);
   U3230 : INV_X1 port map( A => n5915, ZN => n5919);
   U3231 : INV_X1 port map( A => n5915, ZN => n5920);
   U3232 : INV_X1 port map( A => n5915, ZN => n5921);
   U3233 : INV_X1 port map( A => n5916, ZN => n5922);
   U3234 : INV_X1 port map( A => n5916, ZN => n5923);
   U3235 : INV_X1 port map( A => n5924, ZN => n5926);
   U3236 : INV_X1 port map( A => n5924, ZN => n5927);
   U3237 : INV_X1 port map( A => n5422, ZN => n5928);
   U3238 : INV_X1 port map( A => n5925, ZN => n5929);
   U3239 : INV_X1 port map( A => n5925, ZN => n5930);
   U3240 : INV_X1 port map( A => n5925, ZN => n5931);
   U3241 : INV_X1 port map( A => n5925, ZN => n5932);
   U3242 : INV_X1 port map( A => n5934, ZN => n5935);
   U3243 : INV_X1 port map( A => n5934, ZN => n5936);
   U3244 : INV_X1 port map( A => n5933, ZN => n5937);
   U3245 : INV_X1 port map( A => n5933, ZN => n5938);
   U3246 : INV_X1 port map( A => n5934, ZN => n5939);
   U3247 : INV_X1 port map( A => n5934, ZN => n5940);
   U3248 : INV_X1 port map( A => n5934, ZN => n5941);
   U3249 : CLKBUF_X1 port map( A => n6170, Z => n6074);
   U3250 : CLKBUF_X1 port map( A => n6170, Z => n6075);
   U3251 : CLKBUF_X1 port map( A => n6170, Z => n6076);
   U3252 : CLKBUF_X1 port map( A => n6170, Z => n6077);
   U3253 : CLKBUF_X1 port map( A => n6170, Z => n6078);
   U3254 : CLKBUF_X1 port map( A => n6169, Z => n6079);
   U3255 : CLKBUF_X1 port map( A => n6169, Z => n6080);
   U3256 : CLKBUF_X1 port map( A => n6169, Z => n6081);
   U3257 : CLKBUF_X1 port map( A => n6169, Z => n6082);
   U3258 : CLKBUF_X1 port map( A => n6169, Z => n6083);
   U3259 : CLKBUF_X1 port map( A => n6169, Z => n6084);
   U3260 : CLKBUF_X1 port map( A => n6168, Z => n6085);
   U3261 : CLKBUF_X1 port map( A => n6168, Z => n6086);
   U3262 : CLKBUF_X1 port map( A => n6168, Z => n6087);
   U3263 : CLKBUF_X1 port map( A => n6168, Z => n6088);
   U3264 : CLKBUF_X1 port map( A => n6168, Z => n6089);
   U3265 : CLKBUF_X1 port map( A => n6168, Z => n6090);
   U3266 : CLKBUF_X1 port map( A => n6167, Z => n6091);
   U3267 : CLKBUF_X1 port map( A => n6167, Z => n6092);
   U3268 : CLKBUF_X1 port map( A => n6167, Z => n6093);
   U3269 : CLKBUF_X1 port map( A => n6167, Z => n6094);
   U3270 : CLKBUF_X1 port map( A => n6167, Z => n6095);
   U3271 : CLKBUF_X1 port map( A => n6167, Z => n6096);
   U3272 : CLKBUF_X1 port map( A => n6166, Z => n6097);
   U3273 : CLKBUF_X1 port map( A => n6166, Z => n6098);
   U3274 : CLKBUF_X1 port map( A => n6166, Z => n6099);
   U3275 : CLKBUF_X1 port map( A => n6166, Z => n6100);
   U3276 : CLKBUF_X1 port map( A => n6166, Z => n6101);
   U3277 : CLKBUF_X1 port map( A => n6166, Z => n6102);
   U3278 : CLKBUF_X1 port map( A => n6165, Z => n6103);
   U3279 : CLKBUF_X1 port map( A => n6165, Z => n6104);
   U3280 : CLKBUF_X1 port map( A => n6165, Z => n6105);
   U3281 : CLKBUF_X1 port map( A => n6165, Z => n6106);
   U3282 : CLKBUF_X1 port map( A => n6165, Z => n6107);
   U3283 : CLKBUF_X1 port map( A => n6165, Z => n6108);
   U3284 : CLKBUF_X1 port map( A => n6164, Z => n6109);
   U3285 : CLKBUF_X1 port map( A => n6164, Z => n6110);
   U3286 : CLKBUF_X1 port map( A => n6164, Z => n6111);
   U3287 : CLKBUF_X1 port map( A => n6164, Z => n6112);
   U3288 : CLKBUF_X1 port map( A => n6164, Z => n6113);
   U3289 : CLKBUF_X1 port map( A => n6164, Z => n6114);
   U3290 : CLKBUF_X1 port map( A => n6163, Z => n6115);
   U3291 : CLKBUF_X1 port map( A => n6163, Z => n6116);
   U3292 : CLKBUF_X1 port map( A => n6163, Z => n6117);
   U3293 : CLKBUF_X1 port map( A => n6163, Z => n6118);
   U3294 : CLKBUF_X1 port map( A => n6163, Z => n6119);
   U3295 : CLKBUF_X1 port map( A => n6163, Z => n6120);
   U3296 : CLKBUF_X1 port map( A => n6162, Z => n6121);
   U3297 : CLKBUF_X1 port map( A => n6162, Z => n6122);
   U3298 : CLKBUF_X1 port map( A => n6162, Z => n6123);
   U3299 : CLKBUF_X1 port map( A => n6162, Z => n6124);
   U3300 : CLKBUF_X1 port map( A => n6162, Z => n6125);
   U3301 : CLKBUF_X1 port map( A => n6162, Z => n6126);
   U3302 : CLKBUF_X1 port map( A => n6161, Z => n6127);
   U3303 : CLKBUF_X1 port map( A => n6161, Z => n6128);
   U3304 : CLKBUF_X1 port map( A => n6161, Z => n6129);
   U3305 : CLKBUF_X1 port map( A => n6161, Z => n6130);
   U3306 : CLKBUF_X1 port map( A => n6161, Z => n6131);
   U3307 : CLKBUF_X1 port map( A => n6161, Z => n6132);
   U3308 : CLKBUF_X1 port map( A => n6160, Z => n6133);
   U3309 : CLKBUF_X1 port map( A => n6160, Z => n6134);
   U3310 : CLKBUF_X1 port map( A => n6160, Z => n6135);
   U3311 : CLKBUF_X1 port map( A => n6160, Z => n6136);
   U3312 : CLKBUF_X1 port map( A => n6160, Z => n6137);
   U3313 : CLKBUF_X1 port map( A => n6160, Z => n6138);
   U3314 : CLKBUF_X1 port map( A => n6159, Z => n6139);
   U3315 : CLKBUF_X1 port map( A => n6159, Z => n6140);
   U3316 : CLKBUF_X1 port map( A => n6159, Z => n6141);
   U3317 : CLKBUF_X1 port map( A => n6159, Z => n6142);
   U3318 : CLKBUF_X1 port map( A => n6159, Z => n6143);
   U3319 : CLKBUF_X1 port map( A => n6159, Z => n6144);
   U3320 : CLKBUF_X1 port map( A => n6158, Z => n6145);
   U3321 : CLKBUF_X1 port map( A => n6158, Z => n6146);
   U3322 : CLKBUF_X1 port map( A => n6158, Z => n6147);
   U3323 : CLKBUF_X1 port map( A => n6158, Z => n6148);
   U3324 : CLKBUF_X1 port map( A => n6158, Z => n6149);
   U3325 : CLKBUF_X1 port map( A => n6158, Z => n6150);
   U3326 : CLKBUF_X1 port map( A => n6157, Z => n6151);
   U3327 : CLKBUF_X1 port map( A => n6157, Z => n6152);
   U3328 : CLKBUF_X1 port map( A => n6157, Z => n6153);
   U3329 : CLKBUF_X1 port map( A => n6157, Z => n6154);
   U3330 : CLKBUF_X1 port map( A => n6157, Z => n6155);

end SYN_register_file_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Extender_SRC_SIZE26_DEST_SIZE32 is

   port( s : in std_logic;  i : in std_logic_vector (25 downto 0);  o : out 
         std_logic_vector (31 downto 0));

end Extender_SRC_SIZE26_DEST_SIZE32;

architecture SYN_extender_arch of Extender_SRC_SIZE26_DEST_SIZE32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal o_31 : std_logic;

begin
   o <= ( o_31, o_31, o_31, o_31, o_31, o_31, i(25), i(24), i(23), i(22), i(21)
      , i(20), i(19), i(18), i(17), i(16), i(15), i(14), i(13), i(12), i(11), 
      i(10), i(9), i(8), i(7), i(6), i(5), i(4), i(3), i(2), i(1), i(0) );
   
   U1 : AND2_X1 port map( A1 => s, A2 => i(25), ZN => o_31);

end SYN_extender_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Extender_SRC_SIZE16_DEST_SIZE32 is

   port( s : in std_logic;  i : in std_logic_vector (15 downto 0);  o : out 
         std_logic_vector (31 downto 0));

end Extender_SRC_SIZE16_DEST_SIZE32;

architecture SYN_extender_arch of Extender_SRC_SIZE16_DEST_SIZE32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal o_31 : std_logic;

begin
   o <= ( o_31, o_31, o_31, o_31, o_31, o_31, o_31, o_31, o_31, o_31, o_31, 
      o_31, o_31, o_31, o_31, o_31, i(15), i(14), i(13), i(12), i(11), i(10), 
      i(9), i(8), i(7), i(6), i(5), i(4), i(3), i(2), i(1), i(0) );
   
   U1 : AND2_X1 port map( A1 => s, A2 => i(15), ZN => o_31);

end SYN_extender_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE5 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (4 downto 0);  
         dout : out std_logic_vector (4 downto 0));

end Mux_DATA_SIZE5;

architecture SYN_mux_arch of Mux_DATA_SIZE5 is

   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n7, n8, n9, n10, n11, n12 : std_logic;

begin
   
   U1 : INV_X1 port map( A => sel, ZN => n8);
   U2 : INV_X1 port map( A => n12, ZN => dout(0));
   U3 : AOI22_X1 port map( A1 => din0(0), A2 => n8, B1 => din1(0), B2 => sel, 
                           ZN => n12);
   U4 : INV_X1 port map( A => n11, ZN => dout(1));
   U5 : AOI22_X1 port map( A1 => din0(1), A2 => n8, B1 => din1(1), B2 => sel, 
                           ZN => n11);
   U6 : INV_X1 port map( A => n10, ZN => dout(2));
   U7 : AOI22_X1 port map( A1 => din0(2), A2 => n8, B1 => din1(2), B2 => sel, 
                           ZN => n10);
   U8 : INV_X1 port map( A => n9, ZN => dout(3));
   U9 : AOI22_X1 port map( A1 => din0(3), A2 => n8, B1 => din1(3), B2 => sel, 
                           ZN => n9);
   U10 : INV_X1 port map( A => n7, ZN => dout(4));
   U11 : AOI22_X1 port map( A1 => din0(4), A2 => n8, B1 => sel, B2 => din1(4), 
                           ZN => n7);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE32_12 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 0);
         dout : out std_logic_vector (31 downto 0));

end Reg_DATA_SIZE32_12;

architecture SYN_reg_arch of Reg_DATA_SIZE32_12 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, net108873, net108874, net108875, net108876, net108877, 
      net108878, net108879, net108880, net108881, net108882, net108883, 
      net108884, net108885, net108886, net108887, net108888, net108889, 
      net108890, net108891, net108892, net108893, net108894, net108895, 
      net108896, net108897, net108898, net108899, net108900, net108901, 
      net108902, net108903, net108904, n33, n34, n35, n36, n37, n38, n39, n40, 
      n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55
      , n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, 
      n70, n71, n72, n73, n74, n75, n76, n77 : std_logic;

begin
   
   dout_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => n77, Q => 
                           dout(27), QN => net108900);
   dout_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => n76, Q => 
                           dout(26), QN => net108899);
   dout_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => n76, Q => 
                           dout(25), QN => net108898);
   dout_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => n77, Q => 
                           dout(24), QN => net108897);
   dout_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => n76, Q => 
                           dout(23), QN => net108896);
   dout_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => n76, Q => 
                           dout(22), QN => net108895);
   dout_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => n76, Q => 
                           dout(21), QN => net108894);
   dout_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => n76, Q => 
                           dout(20), QN => net108893);
   dout_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => n75, Q => 
                           dout(19), QN => net108892);
   dout_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => n76, Q => 
                           dout(18), QN => net108891);
   dout_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => n75, Q => 
                           dout(17), QN => net108890);
   dout_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => n75, Q => 
                           dout(16), QN => net108889);
   dout_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => n76, Q => 
                           dout(15), QN => net108888);
   dout_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => n75, Q => 
                           dout(12), QN => net108885);
   dout_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => n75, Q => 
                           dout(11), QN => net108884);
   dout_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => n75, Q => 
                           dout(10), QN => net108883);
   dout_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => n76, Q => 
                           dout(8), QN => net108881);
   dout_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => n76, Q => 
                           dout(7), QN => net108880);
   dout_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => n75, Q => 
                           dout(6), QN => net108879);
   dout_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => n76, Q => 
                           dout(5), QN => net108878);
   dout_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => n75, Q => 
                           dout(3), QN => net108876);
   dout_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => n75, Q => 
                           dout(2), QN => net108875);
   dout_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => n75, Q => 
                           dout(1), QN => net108874);
   dout_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => n77, Q => 
                           dout(0), QN => net108873);
   dout_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => n76, Q => 
                           dout(4), QN => net108877);
   dout_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => n75, Q => 
                           dout(14), QN => net108887);
   dout_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => n75, Q => 
                           dout(13), QN => net108886);
   dout_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => n77, Q => 
                           dout(31), QN => net108904);
   dout_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => n77, Q => 
                           dout(9), QN => net108882);
   dout_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => n77, Q => 
                           dout(30), QN => net108903);
   dout_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => n77, Q => 
                           dout(28), QN => net108901);
   dout_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => n77, Q => 
                           dout(29), QN => net108902);
   U2 : BUF_X1 port map( A => en, Z => n69);
   U3 : BUF_X1 port map( A => en, Z => n70);
   U4 : BUF_X1 port map( A => rst, Z => n75);
   U5 : BUF_X1 port map( A => rst, Z => n76);
   U6 : BUF_X1 port map( A => rst, Z => n77);
   U7 : OAI21_X1 port map( B1 => net108883, B2 => n73, A => n50, ZN => n22);
   U8 : NAND2_X1 port map( A1 => din(10), A2 => n70, ZN => n50);
   U9 : OAI21_X1 port map( B1 => net108887, B2 => n73, A => n55, ZN => n18);
   U10 : NAND2_X1 port map( A1 => din(14), A2 => n70, ZN => n55);
   U11 : OAI21_X1 port map( B1 => net108886, B2 => n73, A => n54, ZN => n19);
   U12 : NAND2_X1 port map( A1 => din(13), A2 => n70, ZN => n54);
   U13 : OAI21_X1 port map( B1 => net108882, B2 => n73, A => n49, ZN => n23);
   U14 : NAND2_X1 port map( A1 => din(9), A2 => n71, ZN => n49);
   U15 : OAI21_X1 port map( B1 => net108885, B2 => n73, A => n52, ZN => n20);
   U16 : NAND2_X1 port map( A1 => din(12), A2 => n70, ZN => n52);
   U17 : OAI21_X1 port map( B1 => net108892, B2 => n73, A => n60, ZN => n13);
   U18 : NAND2_X1 port map( A1 => din(19), A2 => n69, ZN => n60);
   U19 : OAI21_X1 port map( B1 => net108900, B2 => n71, A => n37, ZN => n5);
   U20 : NAND2_X1 port map( A1 => din(27), A2 => n69, ZN => n37);
   U21 : OAI21_X1 port map( B1 => net108898, B2 => n71, A => n35, ZN => n7);
   U22 : NAND2_X1 port map( A1 => din(25), A2 => n69, ZN => n35);
   U23 : OAI21_X1 port map( B1 => net108897, B2 => n71, A => n34, ZN => n8);
   U24 : NAND2_X1 port map( A1 => din(24), A2 => n69, ZN => n34);
   U25 : OAI21_X1 port map( B1 => net108874, B2 => n71, A => n40, ZN => n31);
   U26 : NAND2_X1 port map( A1 => din(1), A2 => n70, ZN => n40);
   U27 : OAI21_X1 port map( B1 => net108877, B2 => n72, A => n44, ZN => n28);
   U28 : NAND2_X1 port map( A1 => din(4), A2 => n71, ZN => n44);
   U29 : OAI21_X1 port map( B1 => net108896, B2 => n72, A => n33, ZN => n9);
   U30 : NAND2_X1 port map( A1 => n74, A2 => din(23), ZN => n33);
   U31 : OAI21_X1 port map( B1 => net108881, B2 => n72, A => n48, ZN => n24);
   U32 : NAND2_X1 port map( A1 => din(8), A2 => n71, ZN => n48);
   U33 : OAI21_X1 port map( B1 => net108880, B2 => n72, A => n47, ZN => n25);
   U34 : NAND2_X1 port map( A1 => din(7), A2 => n71, ZN => n47);
   U35 : OAI21_X1 port map( B1 => net108878, B2 => n72, A => n45, ZN => n27);
   U36 : NAND2_X1 port map( A1 => din(5), A2 => n71, ZN => n45);
   U37 : OAI21_X1 port map( B1 => net108879, B2 => n72, A => n46, ZN => n26);
   U38 : NAND2_X1 port map( A1 => din(6), A2 => n71, ZN => n46);
   U39 : OAI21_X1 port map( B1 => net108893, B2 => n74, A => n61, ZN => n12);
   U40 : NAND2_X1 port map( A1 => din(20), A2 => n69, ZN => n61);
   U41 : OAI21_X1 port map( B1 => net108894, B2 => n74, A => n62, ZN => n11);
   U42 : NAND2_X1 port map( A1 => din(21), A2 => n69, ZN => n62);
   U43 : OAI21_X1 port map( B1 => net108895, B2 => n74, A => n63, ZN => n10);
   U44 : NAND2_X1 port map( A1 => din(22), A2 => n69, ZN => n63);
   U45 : OAI21_X1 port map( B1 => net108899, B2 => n72, A => n36, ZN => n6);
   U46 : NAND2_X1 port map( A1 => din(26), A2 => n69, ZN => n36);
   U47 : OAI21_X1 port map( B1 => net108891, B2 => n73, A => n59, ZN => n14);
   U48 : NAND2_X1 port map( A1 => din(18), A2 => n69, ZN => n59);
   U49 : OAI21_X1 port map( B1 => net108890, B2 => n73, A => n58, ZN => n15);
   U50 : NAND2_X1 port map( A1 => din(17), A2 => n69, ZN => n58);
   U51 : OAI21_X1 port map( B1 => net108889, B2 => n73, A => n57, ZN => n16);
   U52 : NAND2_X1 port map( A1 => din(16), A2 => n69, ZN => n57);
   U53 : OAI21_X1 port map( B1 => net108884, B2 => n73, A => n51, ZN => n21);
   U54 : NAND2_X1 port map( A1 => din(11), A2 => n70, ZN => n51);
   U55 : OAI21_X1 port map( B1 => net108888, B2 => n73, A => n56, ZN => n17);
   U56 : NAND2_X1 port map( A1 => din(15), A2 => n70, ZN => n56);
   U57 : OAI21_X1 port map( B1 => net108873, B2 => n72, A => n39, ZN => n32);
   U58 : NAND2_X1 port map( A1 => din(0), A2 => n70, ZN => n39);
   U59 : OAI21_X1 port map( B1 => net108875, B2 => n72, A => n41, ZN => n30);
   U60 : NAND2_X1 port map( A1 => din(2), A2 => n70, ZN => n41);
   U61 : OAI21_X1 port map( B1 => net108876, B2 => n72, A => n43, ZN => n29);
   U62 : NAND2_X1 port map( A1 => din(3), A2 => n70, ZN => n43);
   U63 : OR2_X1 port map( A1 => net108901, A2 => n71, ZN => n65);
   U64 : NAND2_X1 port map( A1 => n38, A2 => n65, ZN => n4);
   U65 : BUF_X1 port map( A => en, Z => n71);
   U66 : OR2_X1 port map( A1 => net108903, A2 => n73, ZN => n66);
   U67 : NAND2_X1 port map( A1 => n53, A2 => n66, ZN => n2);
   U68 : BUF_X1 port map( A => en, Z => n73);
   U69 : OR2_X1 port map( A1 => net108902, A2 => n72, ZN => n67);
   U70 : NAND2_X1 port map( A1 => n42, A2 => n67, ZN => n3);
   U71 : OR2_X1 port map( A1 => net108904, A2 => n72, ZN => n68);
   U72 : NAND2_X1 port map( A1 => n64, A2 => n68, ZN => n1);
   U73 : BUF_X1 port map( A => en, Z => n72);
   U74 : NAND2_X1 port map( A1 => din(28), A2 => n70, ZN => n38);
   U75 : NAND2_X1 port map( A1 => din(29), A2 => n71, ZN => n42);
   U76 : NAND2_X1 port map( A1 => din(30), A2 => n70, ZN => n53);
   U77 : NAND2_X1 port map( A1 => din(31), A2 => n69, ZN => n64);
   U78 : CLKBUF_X1 port map( A => en, Z => n74);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE32_0 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 0);
         dout : out std_logic_vector (31 downto 0));

end Reg_DATA_SIZE32_0;

architecture SYN_reg_arch of Reg_DATA_SIZE32_0 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
      n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93
      , n94, n95, n96, net108097, net108098, net108099, net108100, net108101, 
      net108102, net108103, net108104, net108105, net108106, net108107, 
      net108108, net108109, net108110, net108111, net108112, net108113, 
      net108114, net108115, net108116, net108117, net108118, net108119, 
      net108120, net108121, net108122, net108123, net108124, net108125, 
      net108126, net108127, net108128, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
      n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25
      , n26, n27, n28, n29, n30, n31, n32, n33, n34, n36, n37, n38, n39, n40, 
      n41, n42, n43, n44 : std_logic;

begin
   
   dout_reg_31_inst : DFFR_X1 port map( D => n96, CK => clk, RN => n42, Q => 
                           dout(31), QN => net108128);
   dout_reg_30_inst : DFFR_X1 port map( D => n95, CK => clk, RN => n42, Q => 
                           dout(30), QN => net108127);
   dout_reg_29_inst : DFFR_X1 port map( D => n94, CK => clk, RN => n42, Q => 
                           dout(29), QN => net108126);
   dout_reg_28_inst : DFFR_X1 port map( D => n93, CK => clk, RN => n42, Q => 
                           dout(28), QN => net108125);
   dout_reg_27_inst : DFFR_X1 port map( D => n92, CK => clk, RN => n42, Q => 
                           dout(27), QN => net108124);
   dout_reg_26_inst : DFFR_X1 port map( D => n91, CK => clk, RN => n42, Q => 
                           dout(26), QN => net108123);
   dout_reg_25_inst : DFFR_X1 port map( D => n90, CK => clk, RN => n42, Q => 
                           dout(25), QN => net108122);
   dout_reg_24_inst : DFFR_X1 port map( D => n89, CK => clk, RN => n42, Q => 
                           dout(24), QN => net108121);
   dout_reg_23_inst : DFFR_X1 port map( D => n88, CK => clk, RN => n42, Q => 
                           dout(23), QN => net108120);
   dout_reg_22_inst : DFFR_X1 port map( D => n87, CK => clk, RN => n42, Q => 
                           dout(22), QN => net108119);
   dout_reg_21_inst : DFFR_X1 port map( D => n86, CK => clk, RN => n42, Q => 
                           dout(21), QN => net108118);
   dout_reg_20_inst : DFFR_X1 port map( D => n85, CK => clk, RN => n42, Q => 
                           dout(20), QN => net108117);
   dout_reg_19_inst : DFFR_X1 port map( D => n84, CK => clk, RN => n43, Q => 
                           dout(19), QN => net108116);
   dout_reg_18_inst : DFFR_X1 port map( D => n83, CK => clk, RN => n43, Q => 
                           dout(18), QN => net108115);
   dout_reg_17_inst : DFFR_X1 port map( D => n82, CK => clk, RN => n43, Q => 
                           dout(17), QN => net108114);
   dout_reg_16_inst : DFFR_X1 port map( D => n81, CK => clk, RN => n43, Q => 
                           dout(16), QN => net108113);
   dout_reg_15_inst : DFFR_X1 port map( D => n80, CK => clk, RN => n43, Q => 
                           dout(15), QN => net108112);
   dout_reg_14_inst : DFFR_X1 port map( D => n79, CK => clk, RN => n43, Q => 
                           dout(14), QN => net108111);
   dout_reg_13_inst : DFFR_X1 port map( D => n78, CK => clk, RN => n43, Q => 
                           dout(13), QN => net108110);
   dout_reg_12_inst : DFFR_X1 port map( D => n77, CK => clk, RN => n43, Q => 
                           dout(12), QN => net108109);
   dout_reg_11_inst : DFFR_X1 port map( D => n76, CK => clk, RN => n43, Q => 
                           dout(11), QN => net108108);
   dout_reg_10_inst : DFFR_X1 port map( D => n75, CK => clk, RN => n43, Q => 
                           dout(10), QN => net108107);
   dout_reg_9_inst : DFFR_X1 port map( D => n74, CK => clk, RN => n43, Q => 
                           dout(9), QN => net108106);
   dout_reg_8_inst : DFFR_X1 port map( D => n73, CK => clk, RN => n43, Q => 
                           dout(8), QN => net108105);
   dout_reg_7_inst : DFFR_X1 port map( D => n72, CK => clk, RN => n44, Q => 
                           dout(7), QN => net108104);
   dout_reg_6_inst : DFFR_X1 port map( D => n71, CK => clk, RN => n44, Q => n33
                           , QN => net108103);
   dout_reg_5_inst : DFFR_X1 port map( D => n70, CK => clk, RN => n44, Q => 
                           dout(5), QN => net108102);
   dout_reg_4_inst : DFFR_X1 port map( D => n69, CK => clk, RN => n44, Q => 
                           dout(4), QN => net108101);
   dout_reg_3_inst : DFFR_X1 port map( D => n68, CK => clk, RN => n44, Q => 
                           dout(3), QN => net108100);
   dout_reg_2_inst : DFFR_X1 port map( D => n67, CK => clk, RN => n44, Q => 
                           dout(2), QN => net108099);
   dout_reg_1_inst : DFFR_X1 port map( D => n66, CK => clk, RN => n44, Q => 
                           dout(1), QN => net108098);
   dout_reg_0_inst : DFFR_X1 port map( D => n65, CK => clk, RN => n44, Q => 
                           dout(0), QN => net108097);
   U2 : INV_X1 port map( A => n33, ZN => n34);
   U3 : INV_X2 port map( A => net108103, ZN => dout(6));
   U4 : BUF_X1 port map( A => en, Z => n37);
   U5 : BUF_X1 port map( A => en, Z => n38);
   U6 : BUF_X1 port map( A => en, Z => n39);
   U7 : BUF_X1 port map( A => en, Z => n40);
   U8 : BUF_X1 port map( A => en, Z => n36);
   U9 : BUF_X1 port map( A => rst, Z => n43);
   U10 : BUF_X1 port map( A => rst, Z => n42);
   U11 : BUF_X1 port map( A => rst, Z => n44);
   U12 : NAND2_X1 port map( A1 => din(5), A2 => n36, ZN => n27);
   U13 : NAND2_X1 port map( A1 => din(6), A2 => n36, ZN => n26);
   U14 : NAND2_X1 port map( A1 => din(2), A2 => n36, ZN => n30);
   U15 : NAND2_X1 port map( A1 => din(3), A2 => n36, ZN => n29);
   U16 : OAI21_X1 port map( B1 => net108127, B2 => n38, A => n2, ZN => n95);
   U17 : OAI21_X1 port map( B1 => net108126, B2 => n38, A => n3, ZN => n94);
   U18 : OAI21_X1 port map( B1 => net108123, B2 => n38, A => n6, ZN => n91);
   U19 : NAND2_X1 port map( A1 => din(26), A2 => n37, ZN => n6);
   U20 : OAI21_X1 port map( B1 => net108121, B2 => n38, A => n8, ZN => n89);
   U21 : NAND2_X1 port map( A1 => din(24), A2 => n37, ZN => n8);
   U22 : OAI21_X1 port map( B1 => net108124, B2 => n38, A => n5, ZN => n92);
   U23 : NAND2_X1 port map( A1 => din(27), A2 => n36, ZN => n5);
   U24 : OAI21_X1 port map( B1 => net108125, B2 => n39, A => n4, ZN => n93);
   U25 : OAI21_X1 port map( B1 => net108117, B2 => n39, A => n12, ZN => n85);
   U26 : NAND2_X1 port map( A1 => din(20), A2 => n38, ZN => n12);
   U27 : OAI21_X1 port map( B1 => net108118, B2 => n39, A => n11, ZN => n86);
   U28 : NAND2_X1 port map( A1 => din(21), A2 => n37, ZN => n11);
   U29 : OAI21_X1 port map( B1 => net108119, B2 => n39, A => n10, ZN => n87);
   U30 : NAND2_X1 port map( A1 => din(22), A2 => n38, ZN => n10);
   U31 : OAI21_X1 port map( B1 => net108120, B2 => n39, A => n9, ZN => n88);
   U32 : NAND2_X1 port map( A1 => din(23), A2 => n37, ZN => n9);
   U33 : OAI21_X1 port map( B1 => net108122, B2 => n39, A => n7, ZN => n90);
   U34 : NAND2_X1 port map( A1 => din(25), A2 => n37, ZN => n7);
   U35 : OAI21_X1 port map( B1 => net108113, B2 => n39, A => n16, ZN => n81);
   U36 : NAND2_X1 port map( A1 => din(16), A2 => n38, ZN => n16);
   U37 : OAI21_X1 port map( B1 => net108114, B2 => n39, A => n15, ZN => n82);
   U38 : NAND2_X1 port map( A1 => din(17), A2 => n38, ZN => n15);
   U39 : OAI21_X1 port map( B1 => net108115, B2 => n39, A => n14, ZN => n83);
   U40 : NAND2_X1 port map( A1 => din(18), A2 => n38, ZN => n14);
   U41 : OAI21_X1 port map( B1 => net108116, B2 => n39, A => n13, ZN => n84);
   U42 : NAND2_X1 port map( A1 => din(19), A2 => n38, ZN => n13);
   U43 : OAI21_X1 port map( B1 => net108128, B2 => n39, A => n1, ZN => n96);
   U44 : NAND2_X1 port map( A1 => n41, A2 => din(31), ZN => n1);
   U45 : OAI21_X1 port map( B1 => net108101, B2 => n40, A => n28, ZN => n69);
   U46 : NAND2_X1 port map( A1 => din(4), A2 => n36, ZN => n28);
   U47 : OAI21_X1 port map( B1 => net108104, B2 => n40, A => n25, ZN => n72);
   U48 : NAND2_X1 port map( A1 => din(7), A2 => n36, ZN => n25);
   U49 : OAI21_X1 port map( B1 => net108105, B2 => n40, A => n24, ZN => n73);
   U50 : NAND2_X1 port map( A1 => din(8), A2 => n37, ZN => n24);
   U51 : OAI21_X1 port map( B1 => net108106, B2 => n40, A => n23, ZN => n74);
   U52 : NAND2_X1 port map( A1 => din(9), A2 => n37, ZN => n23);
   U53 : OAI21_X1 port map( B1 => net108107, B2 => n40, A => n22, ZN => n75);
   U54 : NAND2_X1 port map( A1 => din(10), A2 => n37, ZN => n22);
   U55 : OAI21_X1 port map( B1 => net108108, B2 => n40, A => n21, ZN => n76);
   U56 : NAND2_X1 port map( A1 => din(11), A2 => n37, ZN => n21);
   U57 : OAI21_X1 port map( B1 => net108109, B2 => n40, A => n20, ZN => n77);
   U58 : NAND2_X1 port map( A1 => din(12), A2 => n37, ZN => n20);
   U59 : OAI21_X1 port map( B1 => net108110, B2 => n40, A => n19, ZN => n78);
   U60 : NAND2_X1 port map( A1 => din(13), A2 => n37, ZN => n19);
   U61 : OAI21_X1 port map( B1 => net108111, B2 => n40, A => n18, ZN => n79);
   U62 : NAND2_X1 port map( A1 => din(14), A2 => n37, ZN => n18);
   U63 : OAI21_X1 port map( B1 => net108112, B2 => n40, A => n17, ZN => n80);
   U64 : NAND2_X1 port map( A1 => din(15), A2 => n38, ZN => n17);
   U65 : OAI21_X1 port map( B1 => net108097, B2 => n39, A => n32, ZN => n65);
   U66 : OAI21_X1 port map( B1 => net108098, B2 => n41, A => n31, ZN => n66);
   U67 : NAND2_X1 port map( A1 => din(1), A2 => n36, ZN => n31);
   U68 : NAND2_X1 port map( A1 => din(29), A2 => n36, ZN => n3);
   U69 : NAND2_X1 port map( A1 => din(30), A2 => n36, ZN => n2);
   U70 : OAI21_X1 port map( B1 => net108100, B2 => n41, A => n29, ZN => n68);
   U71 : OAI21_X1 port map( B1 => n34, B2 => n40, A => n26, ZN => n71);
   U72 : NAND2_X1 port map( A1 => din(28), A2 => n36, ZN => n4);
   U73 : OAI21_X1 port map( B1 => net108102, B2 => n40, A => n27, ZN => n70);
   U74 : OAI21_X1 port map( B1 => net108099, B2 => n41, A => n30, ZN => n67);
   U75 : NAND2_X1 port map( A1 => din(0), A2 => n36, ZN => n32);
   U76 : CLKBUF_X1 port map( A => en, Z => n41);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE32_0 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0);  
         dout : out std_logic_vector (31 downto 0));

end Mux_DATA_SIZE32_0;

architecture SYN_mux_arch of Mux_DATA_SIZE32_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n34, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, net134004, net134002, net134000, net133998, net133996, 
      net133994, net133992, net133990, net133988, net134014, net134012, n66, n1
      , n2, n3 : std_logic;

begin
   
   U1 : INV_X2 port map( A => n44, ZN => dout(2));
   U2 : INV_X1 port map( A => n39, ZN => dout(5));
   U3 : INV_X1 port map( A => n34, ZN => dout(9));
   U4 : INV_X1 port map( A => n57, ZN => dout(18));
   U5 : BUF_X1 port map( A => n3, Z => n2);
   U6 : AOI22_X1 port map( A1 => din0(0), A2 => net133990, B1 => din1(0), B2 =>
                           n1, ZN => n66);
   U7 : INV_X1 port map( A => n66, ZN => dout(0));
   U8 : CLKBUF_X1 port map( A => n3, Z => n1);
   U9 : AOI22_X1 port map( A1 => din0(11), A2 => net133988, B1 => din1(11), B2 
                           => n1, ZN => n64);
   U10 : AOI22_X1 port map( A1 => din0(10), A2 => net133988, B1 => din1(10), B2
                           => n1, ZN => n65);
   U11 : AOI22_X1 port map( A1 => din0(9), A2 => net133990, B1 => n1, B2 => 
                           din1(9), ZN => n34);
   U12 : BUF_X1 port map( A => sel, Z => n3);
   U13 : CLKBUF_X1 port map( A => n3, Z => net134004);
   U14 : INV_X1 port map( A => n2, ZN => net133988);
   U15 : INV_X1 port map( A => n2, ZN => net133990);
   U16 : CLKBUF_X1 port map( A => sel, Z => net134014);
   U17 : CLKBUF_X1 port map( A => sel, Z => net134012);
   U18 : INV_X1 port map( A => n58, ZN => dout(17));
   U19 : INV_X1 port map( A => n55, ZN => dout(1));
   U20 : INV_X1 port map( A => n63, ZN => dout(12));
   U21 : INV_X1 port map( A => n40, ZN => dout(4));
   U22 : CLKBUF_X1 port map( A => net134014, Z => net134002);
   U23 : BUF_X1 port map( A => net134012, Z => net133994);
   U24 : CLKBUF_X1 port map( A => net134012, Z => net133992);
   U25 : BUF_X1 port map( A => net134014, Z => net134000);
   U26 : CLKBUF_X1 port map( A => net134014, Z => net133998);
   U27 : CLKBUF_X1 port map( A => net134012, Z => net133996);
   U28 : INV_X1 port map( A => n56, ZN => dout(19));
   U29 : AOI22_X1 port map( A1 => din0(19), A2 => net133990, B1 => din1(19), B2
                           => net134002, ZN => n56);
   U30 : INV_X1 port map( A => n50, ZN => dout(24));
   U31 : AOI22_X1 port map( A1 => din0(24), A2 => net133988, B1 => din1(24), B2
                           => net133998, ZN => n50);
   U32 : INV_X1 port map( A => n54, ZN => dout(20));
   U33 : AOI22_X1 port map( A1 => din0(20), A2 => net133988, B1 => din1(20), B2
                           => net134000, ZN => n54);
   U34 : INV_X1 port map( A => n49, ZN => dout(25));
   U35 : AOI22_X1 port map( A1 => din0(25), A2 => net133988, B1 => din1(25), B2
                           => net133998, ZN => n49);
   U36 : INV_X1 port map( A => n48, ZN => dout(26));
   U37 : AOI22_X1 port map( A1 => din0(26), A2 => net133988, B1 => din1(26), B2
                           => net133996, ZN => n48);
   U38 : INV_X1 port map( A => n53, ZN => dout(21));
   U39 : AOI22_X1 port map( A1 => din0(21), A2 => net133988, B1 => din1(21), B2
                           => net134000, ZN => n53);
   U40 : INV_X1 port map( A => n52, ZN => dout(22));
   U41 : AOI22_X1 port map( A1 => din0(22), A2 => net133988, B1 => din1(22), B2
                           => net133998, ZN => n52);
   U42 : AOI22_X1 port map( A1 => din0(2), A2 => net133988, B1 => din1(2), B2 
                           => net133994, ZN => n44);
   U43 : INV_X1 port map( A => n51, ZN => dout(23));
   U44 : AOI22_X1 port map( A1 => din0(23), A2 => net133988, B1 => din1(23), B2
                           => net133998, ZN => n51);
   U45 : INV_X1 port map( A => n65, ZN => dout(10));
   U46 : INV_X1 port map( A => n60, ZN => dout(15));
   U47 : AOI22_X1 port map( A1 => din0(15), A2 => net133988, B1 => din1(15), B2
                           => net134004, ZN => n60);
   U48 : AOI22_X1 port map( A1 => din0(12), A2 => net133988, B1 => din1(12), B2
                           => net134004, ZN => n63);
   U49 : INV_X1 port map( A => n42, ZN => dout(31));
   U50 : AOI22_X1 port map( A1 => din0(31), A2 => net133990, B1 => din1(31), B2
                           => net133994, ZN => n42);
   U51 : AOI22_X1 port map( A1 => din0(5), A2 => net133990, B1 => din1(5), B2 
                           => net133992, ZN => n39);
   U52 : INV_X1 port map( A => n47, ZN => dout(27));
   U53 : INV_X1 port map( A => n36, ZN => dout(8));
   U54 : AOI22_X1 port map( A1 => din0(8), A2 => net133990, B1 => din1(8), B2 
                           => net133992, ZN => n36);
   U55 : INV_X1 port map( A => n62, ZN => dout(13));
   U56 : INV_X1 port map( A => n59, ZN => dout(16));
   U57 : AOI22_X1 port map( A1 => din0(16), A2 => net133988, B1 => din1(16), B2
                           => net134002, ZN => n59);
   U58 : INV_X1 port map( A => n41, ZN => dout(3));
   U59 : AOI22_X1 port map( A1 => din0(3), A2 => net133990, B1 => din1(3), B2 
                           => net133994, ZN => n41);
   U60 : AOI22_X1 port map( A1 => din0(4), A2 => net133990, B1 => din1(4), B2 
                           => net133994, ZN => n40);
   U61 : INV_X1 port map( A => n61, ZN => dout(14));
   U62 : AOI22_X1 port map( A1 => din0(14), A2 => net133988, B1 => din1(14), B2
                           => net134004, ZN => n61);
   U63 : AOI22_X1 port map( A1 => din0(17), A2 => net133988, B1 => din1(17), B2
                           => net134002, ZN => n58);
   U64 : AOI22_X1 port map( A1 => din0(18), A2 => net133988, B1 => din1(18), B2
                           => net134002, ZN => n57);
   U65 : INV_X1 port map( A => n37, ZN => dout(7));
   U66 : AOI22_X1 port map( A1 => din0(7), A2 => net133990, B1 => din1(7), B2 
                           => net133992, ZN => n37);
   U67 : INV_X1 port map( A => n38, ZN => dout(6));
   U68 : AOI22_X1 port map( A1 => din0(6), A2 => net133990, B1 => din1(6), B2 
                           => net133992, ZN => n38);
   U69 : AOI22_X1 port map( A1 => din0(1), A2 => net133988, B1 => din1(1), B2 
                           => net134000, ZN => n55);
   U70 : INV_X1 port map( A => n43, ZN => dout(30));
   U71 : INV_X1 port map( A => n45, ZN => dout(29));
   U72 : AOI22_X1 port map( A1 => din0(29), A2 => net133988, B1 => din1(29), B2
                           => net133996, ZN => n45);
   U73 : AOI22_X1 port map( A1 => din0(30), A2 => net133988, B1 => din1(30), B2
                           => net134000, ZN => n43);
   U74 : AOI22_X1 port map( A1 => din0(13), A2 => net133988, B1 => din1(13), B2
                           => net134004, ZN => n62);
   U75 : AOI22_X1 port map( A1 => din0(27), A2 => net133988, B1 => din1(27), B2
                           => net133996, ZN => n47);
   U76 : INV_X1 port map( A => n64, ZN => dout(11));
   U77 : AOI22_X1 port map( A1 => din0(28), A2 => net133988, B1 => din1(28), B2
                           => net133996, ZN => n46);
   U78 : INV_X1 port map( A => n46, ZN => dout(28));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Adder_DATA_SIZE32_0 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end Adder_DATA_SIZE32_0;

architecture SYN_adder_arch of Adder_DATA_SIZE32_0 is

   component P4Adder_DATA_SIZE32_SPARSITY4_0
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;

begin
   
   ADDER0 : P4Adder_DATA_SIZE32_SPARSITY4_0 port map( cin => cin, a(31) => 
                           a(31), a(30) => a(30), a(29) => a(29), a(28) => 
                           a(28), a(27) => a(27), a(26) => a(26), a(25) => 
                           a(25), a(24) => a(24), a(23) => a(23), a(22) => 
                           a(22), a(21) => a(21), a(20) => a(20), a(19) => 
                           a(19), a(18) => a(18), a(17) => a(17), a(16) => 
                           a(16), a(15) => a(15), a(14) => a(14), a(13) => 
                           a(13), a(12) => a(12), a(11) => a(11), a(10) => 
                           a(10), a(9) => a(9), a(8) => a(8), a(7) => a(7), 
                           a(6) => a(6), a(5) => a(5), a(4) => a(4), a(3) => 
                           a(3), a(2) => a(2), a(1) => a(1), a(0) => a(0), 
                           b(31) => b(31), b(30) => b(30), b(29) => b(29), 
                           b(28) => b(28), b(27) => b(27), b(26) => b(26), 
                           b(25) => b(25), b(24) => b(24), b(23) => b(23), 
                           b(22) => b(22), b(21) => b(21), b(20) => b(20), 
                           b(19) => b(19), b(18) => b(18), b(17) => b(17), 
                           b(16) => b(16), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           s(31) => s(31), s(30) => s(30), s(29) => s(29), 
                           s(28) => s(28), s(27) => s(27), s(26) => s(26), 
                           s(25) => s(25), s(24) => s(24), s(23) => s(23), 
                           s(22) => s(22), s(21) => s(21), s(20) => s(20), 
                           s(19) => s(19), s(18) => s(18), s(17) => s(17), 
                           s(16) => s(16), s(15) => s(15), s(14) => s(14), 
                           s(13) => s(13), s(12) => s(12), s(11) => s(11), 
                           s(10) => s(10), s(9) => s(9), s(8) => s(8), s(7) => 
                           s(7), s(6) => s(6), s(5) => s(5), s(4) => s(4), s(3)
                           => s(3), s(2) => s(2), s(1) => s(1), s(0) => s(0), 
                           cout => cout);

end SYN_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Branch_DATA_SIZE32_OPCD_SIZE6_ADDR_SIZE32 is

   port( rst, clk : in std_logic;  reg_a, ld_a : in std_logic_vector (31 downto
         0);  opcd : in std_logic_vector (5 downto 0);  addr : in 
         std_logic_vector (31 downto 0);  sig_bal : in std_logic;  sig_bpw, 
         sig_brt : out std_logic);

end Branch_DATA_SIZE32_OPCD_SIZE6_ADDR_SIZE32;

architecture SYN_branch_arch of Branch_DATA_SIZE32_OPCD_SIZE6_ADDR_SIZE32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X2
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal bht_0_26_port, bht_0_25_port, bht_0_24_port, bht_0_23_port, 
      bht_0_22_port, bht_0_21_port, bht_0_20_port, bht_0_19_port, bht_0_18_port
      , bht_0_17_port, bht_0_16_port, bht_0_15_port, bht_0_14_port, 
      bht_0_13_port, bht_0_12_port, bht_0_11_port, bht_0_10_port, bht_0_9_port,
      bht_0_8_port, bht_0_7_port, bht_0_6_port, bht_0_5_port, bht_0_4_port, 
      bht_0_3_port, bht_0_2_port, bht_0_1_port, bht_0_0_port, bht_1_26_port, 
      bht_1_25_port, bht_1_24_port, bht_1_23_port, bht_1_22_port, bht_1_21_port
      , bht_1_20_port, bht_1_19_port, bht_1_18_port, bht_1_17_port, 
      bht_1_16_port, bht_1_15_port, bht_1_14_port, bht_1_13_port, bht_1_12_port
      , bht_1_11_port, bht_1_10_port, bht_1_9_port, bht_1_8_port, bht_1_7_port,
      bht_1_6_port, bht_1_5_port, bht_1_4_port, bht_1_3_port, bht_1_2_port, 
      bht_1_1_port, bht_1_0_port, bht_2_26_port, bht_2_25_port, bht_2_24_port, 
      bht_2_23_port, bht_2_22_port, bht_2_21_port, bht_2_20_port, bht_2_19_port
      , bht_2_18_port, bht_2_17_port, bht_2_16_port, bht_2_15_port, 
      bht_2_14_port, bht_2_13_port, bht_2_12_port, bht_2_11_port, bht_2_10_port
      , bht_2_9_port, bht_2_8_port, bht_2_7_port, bht_2_6_port, bht_2_5_port, 
      bht_2_4_port, bht_2_3_port, bht_2_2_port, bht_2_1_port, bht_2_0_port, 
      bht_3_26_port, bht_3_25_port, bht_3_24_port, bht_3_23_port, bht_3_22_port
      , bht_3_21_port, bht_3_20_port, bht_3_19_port, bht_3_18_port, 
      bht_3_17_port, bht_3_16_port, bht_3_15_port, bht_3_14_port, bht_3_13_port
      , bht_3_12_port, bht_3_11_port, bht_3_10_port, bht_3_9_port, bht_3_8_port
      , bht_3_7_port, bht_3_6_port, bht_3_5_port, bht_3_4_port, bht_3_3_port, 
      bht_3_2_port, bht_3_1_port, bht_3_0_port, bht_4_26_port, bht_4_25_port, 
      bht_4_24_port, bht_4_23_port, bht_4_22_port, bht_4_21_port, bht_4_20_port
      , bht_4_19_port, bht_4_18_port, bht_4_17_port, bht_4_16_port, 
      bht_4_15_port, bht_4_14_port, bht_4_13_port, bht_4_12_port, bht_4_11_port
      , bht_4_10_port, bht_4_9_port, bht_4_8_port, bht_4_7_port, bht_4_6_port, 
      bht_4_5_port, bht_4_4_port, bht_4_3_port, bht_4_2_port, bht_4_1_port, 
      bht_4_0_port, bht_5_26_port, bht_5_25_port, bht_5_24_port, bht_5_23_port,
      bht_5_22_port, bht_5_21_port, bht_5_20_port, bht_5_19_port, bht_5_18_port
      , bht_5_17_port, bht_5_16_port, bht_5_15_port, bht_5_14_port, 
      bht_5_13_port, bht_5_12_port, bht_5_11_port, bht_5_10_port, bht_5_9_port,
      bht_5_8_port, bht_5_7_port, bht_5_6_port, bht_5_5_port, bht_5_4_port, 
      bht_5_3_port, bht_5_2_port, bht_5_1_port, bht_5_0_port, bht_6_26_port, 
      bht_6_25_port, bht_6_24_port, bht_6_23_port, bht_6_22_port, bht_6_21_port
      , bht_6_20_port, bht_6_19_port, bht_6_18_port, bht_6_17_port, 
      bht_6_16_port, bht_6_15_port, bht_6_14_port, bht_6_13_port, bht_6_12_port
      , bht_6_11_port, bht_6_10_port, bht_6_9_port, bht_6_8_port, bht_6_7_port,
      bht_6_6_port, bht_6_5_port, bht_6_4_port, bht_6_3_port, bht_6_2_port, 
      bht_6_1_port, bht_6_0_port, bht_7_26_port, bht_7_25_port, bht_7_24_port, 
      bht_7_23_port, bht_7_22_port, bht_7_21_port, bht_7_20_port, bht_7_19_port
      , bht_7_18_port, bht_7_17_port, bht_7_16_port, bht_7_15_port, 
      bht_7_14_port, bht_7_13_port, bht_7_12_port, bht_7_11_port, bht_7_10_port
      , bht_7_9_port, bht_7_8_port, bht_7_7_port, bht_7_6_port, bht_7_5_port, 
      bht_7_4_port, bht_7_3_port, bht_7_2_port, bht_7_1_port, bht_7_0_port, 
      bht_8_26_port, bht_8_25_port, bht_8_24_port, bht_8_23_port, bht_8_22_port
      , bht_8_21_port, bht_8_20_port, bht_8_19_port, bht_8_18_port, 
      bht_8_17_port, bht_8_16_port, bht_8_15_port, bht_8_14_port, bht_8_13_port
      , bht_8_12_port, bht_8_11_port, bht_8_10_port, bht_8_9_port, bht_8_8_port
      , bht_8_7_port, bht_8_6_port, bht_8_5_port, bht_8_4_port, bht_8_3_port, 
      bht_8_2_port, bht_8_1_port, bht_8_0_port, bht_9_26_port, bht_9_25_port, 
      bht_9_24_port, bht_9_23_port, bht_9_22_port, bht_9_21_port, bht_9_20_port
      , bht_9_19_port, bht_9_18_port, bht_9_17_port, bht_9_16_port, 
      bht_9_15_port, bht_9_14_port, bht_9_13_port, bht_9_12_port, bht_9_11_port
      , bht_9_10_port, bht_9_9_port, bht_9_8_port, bht_9_7_port, bht_9_6_port, 
      bht_9_5_port, bht_9_4_port, bht_9_3_port, bht_9_2_port, bht_9_1_port, 
      bht_9_0_port, bht_10_26_port, bht_10_25_port, bht_10_24_port, 
      bht_10_23_port, bht_10_22_port, bht_10_21_port, bht_10_20_port, 
      bht_10_19_port, bht_10_18_port, bht_10_17_port, bht_10_16_port, 
      bht_10_15_port, bht_10_14_port, bht_10_13_port, bht_10_12_port, 
      bht_10_11_port, bht_10_10_port, bht_10_9_port, bht_10_8_port, 
      bht_10_7_port, bht_10_6_port, bht_10_5_port, bht_10_4_port, bht_10_3_port
      , bht_10_2_port, bht_10_1_port, bht_10_0_port, bht_11_26_port, 
      bht_11_25_port, bht_11_24_port, bht_11_23_port, bht_11_22_port, 
      bht_11_21_port, bht_11_20_port, bht_11_19_port, bht_11_18_port, 
      bht_11_17_port, bht_11_16_port, bht_11_15_port, bht_11_14_port, 
      bht_11_13_port, bht_11_12_port, bht_11_11_port, bht_11_10_port, 
      bht_11_9_port, bht_11_8_port, bht_11_7_port, bht_11_6_port, bht_11_5_port
      , bht_11_4_port, bht_11_3_port, bht_11_2_port, bht_11_1_port, 
      bht_11_0_port, bht_12_26_port, bht_12_25_port, bht_12_24_port, 
      bht_12_23_port, bht_12_22_port, bht_12_21_port, bht_12_20_port, 
      bht_12_19_port, bht_12_18_port, bht_12_17_port, bht_12_16_port, 
      bht_12_15_port, bht_12_14_port, bht_12_13_port, bht_12_12_port, 
      bht_12_11_port, bht_12_10_port, bht_12_9_port, bht_12_8_port, 
      bht_12_7_port, bht_12_6_port, bht_12_5_port, bht_12_4_port, bht_12_3_port
      , bht_12_2_port, bht_12_1_port, bht_12_0_port, bht_13_26_port, 
      bht_13_25_port, bht_13_24_port, bht_13_23_port, bht_13_22_port, 
      bht_13_21_port, bht_13_20_port, bht_13_19_port, bht_13_18_port, 
      bht_13_17_port, bht_13_16_port, bht_13_15_port, bht_13_14_port, 
      bht_13_13_port, bht_13_12_port, bht_13_11_port, bht_13_10_port, 
      bht_13_9_port, bht_13_8_port, bht_13_7_port, bht_13_6_port, bht_13_5_port
      , bht_13_4_port, bht_13_3_port, bht_13_2_port, bht_13_1_port, 
      bht_13_0_port, bht_14_26_port, bht_14_25_port, bht_14_24_port, 
      bht_14_23_port, bht_14_22_port, bht_14_21_port, bht_14_20_port, 
      bht_14_19_port, bht_14_18_port, bht_14_17_port, bht_14_16_port, 
      bht_14_15_port, bht_14_14_port, bht_14_13_port, bht_14_12_port, 
      bht_14_11_port, bht_14_10_port, bht_14_9_port, bht_14_8_port, 
      bht_14_7_port, bht_14_6_port, bht_14_5_port, bht_14_4_port, bht_14_3_port
      , bht_14_2_port, bht_14_1_port, bht_14_0_port, bht_15_26_port, 
      bht_15_25_port, bht_15_24_port, bht_15_23_port, bht_15_22_port, 
      bht_15_21_port, bht_15_20_port, bht_15_19_port, bht_15_18_port, 
      bht_15_17_port, bht_15_16_port, bht_15_15_port, bht_15_14_port, 
      bht_15_13_port, bht_15_12_port, bht_15_11_port, bht_15_10_port, 
      bht_15_9_port, bht_15_8_port, bht_15_7_port, bht_15_6_port, bht_15_5_port
      , bht_15_4_port, bht_15_3_port, bht_15_2_port, bht_15_1_port, 
      bht_15_0_port, bht_16_26_port, bht_16_25_port, bht_16_24_port, 
      bht_16_23_port, bht_16_22_port, bht_16_21_port, bht_16_20_port, 
      bht_16_19_port, bht_16_18_port, bht_16_17_port, bht_16_16_port, 
      bht_16_15_port, bht_16_14_port, bht_16_13_port, bht_16_12_port, 
      bht_16_11_port, bht_16_10_port, bht_16_9_port, bht_16_8_port, 
      bht_16_7_port, bht_16_6_port, bht_16_5_port, bht_16_4_port, bht_16_3_port
      , bht_16_2_port, bht_16_1_port, bht_16_0_port, bht_17_26_port, 
      bht_17_25_port, bht_17_24_port, bht_17_23_port, bht_17_22_port, 
      bht_17_21_port, bht_17_20_port, bht_17_19_port, bht_17_18_port, 
      bht_17_17_port, bht_17_16_port, bht_17_15_port, bht_17_14_port, 
      bht_17_13_port, bht_17_12_port, bht_17_11_port, bht_17_10_port, 
      bht_17_9_port, bht_17_8_port, bht_17_7_port, bht_17_6_port, bht_17_5_port
      , bht_17_4_port, bht_17_3_port, bht_17_2_port, bht_17_1_port, 
      bht_17_0_port, bht_18_26_port, bht_18_25_port, bht_18_24_port, 
      bht_18_23_port, bht_18_22_port, bht_18_21_port, bht_18_20_port, 
      bht_18_19_port, bht_18_18_port, bht_18_17_port, bht_18_16_port, 
      bht_18_15_port, bht_18_14_port, bht_18_13_port, bht_18_12_port, 
      bht_18_11_port, bht_18_10_port, bht_18_9_port, bht_18_8_port, 
      bht_18_7_port, bht_18_6_port, bht_18_5_port, bht_18_4_port, bht_18_3_port
      , bht_18_2_port, bht_18_1_port, bht_18_0_port, bht_19_26_port, 
      bht_19_25_port, bht_19_24_port, bht_19_23_port, bht_19_22_port, 
      bht_19_21_port, bht_19_20_port, bht_19_19_port, bht_19_18_port, 
      bht_19_17_port, bht_19_16_port, bht_19_15_port, bht_19_14_port, 
      bht_19_13_port, bht_19_12_port, bht_19_11_port, bht_19_10_port, 
      bht_19_9_port, bht_19_8_port, bht_19_7_port, bht_19_6_port, bht_19_5_port
      , bht_19_4_port, bht_19_3_port, bht_19_2_port, bht_19_1_port, 
      bht_19_0_port, bht_20_26_port, bht_20_25_port, bht_20_24_port, 
      bht_20_23_port, bht_20_22_port, bht_20_21_port, bht_20_20_port, 
      bht_20_19_port, bht_20_18_port, bht_20_17_port, bht_20_16_port, 
      bht_20_15_port, bht_20_14_port, bht_20_13_port, bht_20_12_port, 
      bht_20_11_port, bht_20_10_port, bht_20_9_port, bht_20_8_port, 
      bht_20_7_port, bht_20_6_port, bht_20_5_port, bht_20_4_port, bht_20_3_port
      , bht_20_2_port, bht_20_1_port, bht_20_0_port, bht_21_26_port, 
      bht_21_25_port, bht_21_24_port, bht_21_23_port, bht_21_22_port, 
      bht_21_21_port, bht_21_20_port, bht_21_19_port, bht_21_18_port, 
      bht_21_17_port, bht_21_16_port, bht_21_15_port, bht_21_14_port, 
      bht_21_13_port, bht_21_12_port, bht_21_11_port, bht_21_10_port, 
      bht_21_9_port, bht_21_8_port, bht_21_7_port, bht_21_6_port, bht_21_5_port
      , bht_21_4_port, bht_21_3_port, bht_21_2_port, bht_21_1_port, 
      bht_21_0_port, bht_22_26_port, bht_22_25_port, bht_22_24_port, 
      bht_22_23_port, bht_22_22_port, bht_22_21_port, bht_22_20_port, 
      bht_22_19_port, bht_22_18_port, bht_22_17_port, bht_22_16_port, 
      bht_22_15_port, bht_22_14_port, bht_22_13_port, bht_22_12_port, 
      bht_22_11_port, bht_22_10_port, bht_22_9_port, bht_22_8_port, 
      bht_22_7_port, bht_22_6_port, bht_22_5_port, bht_22_4_port, bht_22_3_port
      , bht_22_2_port, bht_22_1_port, bht_22_0_port, bht_23_26_port, 
      bht_23_25_port, bht_23_24_port, bht_23_23_port, bht_23_22_port, 
      bht_23_21_port, bht_23_20_port, bht_23_19_port, bht_23_18_port, 
      bht_23_17_port, bht_23_16_port, bht_23_15_port, bht_23_14_port, 
      bht_23_13_port, bht_23_12_port, bht_23_11_port, bht_23_10_port, 
      bht_23_9_port, bht_23_8_port, bht_23_7_port, bht_23_6_port, bht_23_5_port
      , bht_23_4_port, bht_23_3_port, bht_23_2_port, bht_23_1_port, 
      bht_23_0_port, bht_24_26_port, bht_24_25_port, bht_24_24_port, 
      bht_24_23_port, bht_24_22_port, bht_24_21_port, bht_24_20_port, 
      bht_24_19_port, bht_24_18_port, bht_24_17_port, bht_24_16_port, 
      bht_24_15_port, bht_24_14_port, bht_24_13_port, bht_24_12_port, 
      bht_24_11_port, bht_24_10_port, bht_24_9_port, bht_24_8_port, 
      bht_24_7_port, bht_24_6_port, bht_24_5_port, bht_24_4_port, bht_24_3_port
      , bht_24_2_port, bht_24_1_port, bht_24_0_port, bht_25_26_port, 
      bht_25_25_port, bht_25_24_port, bht_25_23_port, bht_25_22_port, 
      bht_25_21_port, bht_25_20_port, bht_25_19_port, bht_25_18_port, 
      bht_25_17_port, bht_25_16_port, bht_25_15_port, bht_25_14_port, 
      bht_25_13_port, bht_25_12_port, bht_25_11_port, bht_25_10_port, 
      bht_25_9_port, bht_25_8_port, bht_25_7_port, bht_25_6_port, bht_25_5_port
      , bht_25_4_port, bht_25_3_port, bht_25_2_port, bht_25_1_port, 
      bht_25_0_port, bht_26_26_port, bht_26_25_port, bht_26_24_port, 
      bht_26_23_port, bht_26_22_port, bht_26_21_port, bht_26_20_port, 
      bht_26_19_port, bht_26_18_port, bht_26_17_port, bht_26_16_port, 
      bht_26_15_port, bht_26_14_port, bht_26_13_port, bht_26_12_port, 
      bht_26_11_port, bht_26_10_port, bht_26_9_port, bht_26_8_port, 
      bht_26_7_port, bht_26_6_port, bht_26_5_port, bht_26_4_port, bht_26_3_port
      , bht_26_2_port, bht_26_1_port, bht_26_0_port, bht_27_26_port, 
      bht_27_25_port, bht_27_24_port, bht_27_23_port, bht_27_22_port, 
      bht_27_21_port, bht_27_20_port, bht_27_19_port, bht_27_18_port, 
      bht_27_17_port, bht_27_16_port, bht_27_15_port, bht_27_14_port, 
      bht_27_13_port, bht_27_12_port, bht_27_11_port, bht_27_10_port, 
      bht_27_9_port, bht_27_8_port, bht_27_7_port, bht_27_6_port, bht_27_5_port
      , bht_27_4_port, bht_27_3_port, bht_27_2_port, bht_27_1_port, 
      bht_27_0_port, bht_28_26_port, bht_28_25_port, bht_28_24_port, 
      bht_28_23_port, bht_28_22_port, bht_28_21_port, bht_28_20_port, 
      bht_28_19_port, bht_28_18_port, bht_28_17_port, bht_28_16_port, 
      bht_28_15_port, bht_28_14_port, bht_28_13_port, bht_28_12_port, 
      bht_28_11_port, bht_28_10_port, bht_28_9_port, bht_28_8_port, 
      bht_28_7_port, bht_28_6_port, bht_28_5_port, bht_28_4_port, bht_28_3_port
      , bht_28_2_port, bht_28_1_port, bht_28_0_port, bht_29_26_port, 
      bht_29_25_port, bht_29_24_port, bht_29_23_port, bht_29_22_port, 
      bht_29_21_port, bht_29_20_port, bht_29_19_port, bht_29_18_port, 
      bht_29_17_port, bht_29_16_port, bht_29_15_port, bht_29_14_port, 
      bht_29_13_port, bht_29_12_port, bht_29_11_port, bht_29_10_port, 
      bht_29_9_port, bht_29_8_port, bht_29_7_port, bht_29_6_port, bht_29_5_port
      , bht_29_4_port, bht_29_3_port, bht_29_2_port, bht_29_1_port, 
      bht_29_0_port, bht_30_26_port, bht_30_25_port, bht_30_24_port, 
      bht_30_23_port, bht_30_22_port, bht_30_21_port, bht_30_20_port, 
      bht_30_19_port, bht_30_18_port, bht_30_17_port, bht_30_16_port, 
      bht_30_15_port, bht_30_14_port, bht_30_13_port, bht_30_12_port, 
      bht_30_11_port, bht_30_10_port, bht_30_9_port, bht_30_8_port, 
      bht_30_7_port, bht_30_6_port, bht_30_5_port, bht_30_4_port, bht_30_3_port
      , bht_30_2_port, bht_30_1_port, bht_30_0_port, bht_31_26_port, 
      bht_31_25_port, bht_31_24_port, bht_31_23_port, bht_31_22_port, 
      bht_31_21_port, bht_31_20_port, bht_31_19_port, bht_31_18_port, 
      bht_31_17_port, bht_31_16_port, bht_31_15_port, bht_31_14_port, 
      bht_31_13_port, bht_31_12_port, bht_31_11_port, bht_31_10_port, 
      bht_31_9_port, bht_31_8_port, bht_31_7_port, bht_31_6_port, bht_31_5_port
      , bht_31_4_port, bht_31_3_port, bht_31_2_port, bht_31_1_port, 
      bht_31_0_port, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134
      , N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146,
      N147, N148, N149, N150, N151, index_r_4_port, index_r_3_port, 
      index_r_2_port, index_r_1_port, index_r_0_port, entry_r_26_port, 
      entry_r_25_port, entry_r_24_port, entry_r_23_port, entry_r_22_port, 
      entry_r_21_port, entry_r_20_port, entry_r_19_port, entry_r_18_port, 
      entry_r_17_port, entry_r_16_port, entry_r_15_port, entry_r_14_port, 
      entry_r_13_port, entry_r_12_port, entry_r_11_port, entry_r_10_port, 
      entry_r_9_port, entry_r_8_port, entry_r_7_port, entry_r_6_port, 
      entry_r_5_port, entry_r_4_port, entry_r_3_port, entry_r_2_port, 
      entry_r_1_port, entry_r_0_port, N188, sig_bal_delay, opcd_delay_5_port, 
      opcd_delay_4_port, opcd_delay_3_port, opcd_delay_2_port, sig_brt_delay, 
      N2110, N2164, N2218, N2272, N2326, N2380, N2434, N2488, N2542, N2596, 
      N2650, N2704, N2758, N2812, N2866, N2920, N2974, N3028, N3082, N3136, 
      N3190, N3244, N3298, N3352, N3406, N3460, N3514, N3568, N3622, N3676, 
      N3730, N3733, N3735, N3737, N3739, N3741, N3743, N3745, N3747, N3749, 
      N3751, N3753, N3755, N3757, N3759, N3761, N3763, N3765, N3767, N3769, 
      N3771, N3773, N3775, N3777, N3779, N3781, N3783, N3784, N3785, n200, n214
      , n219, n4, n5, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , net108064, net108065, net108066, net108067, net108068, net108069, 
      net108070, net108071, net108072, net108073, net108074, net108075, 
      net108076, net108077, net108078, net108079, net108080, net108081, 
      net108082, net108083, net108084, net108085, net108086, net108087, 
      net108088, net108089, net108090, net108091, net108092, net108093, 
      net108094, net108095, net108096, n91, n94, n97, n98, n100, n101, n103, 
      n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, 
      n116, n117, n118, n120, n121, n122, n123, n124, n125_port, n126_port, 
      n127_port, n130_port, n131_port, n132_port, n137_port, n139_port, 
      n140_port, n141_port, n142_port, n143_port, n144_port, n145_port, 
      n146_port, n147_port, n148_port, n149_port, n150_port, n151_port, n152, 
      n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, 
      n165, n166, n167, n168, n169, n170, n171, n172, n174, n175, n176, n177, 
      n178, n179, n180, n181, n182, n183, n184, n185, n186, n188_port, n189, 
      n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n201, n203, 
      n204, n205, n206, n208, n209, n210, n211, n212, n213, n215, n216, n217, 
      n218, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n278, n279, 
      n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, 
      n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, 
      n304, n305, n306, n311, n312, n313, n314, n315, n316, n317, n318, n319, 
      n320, n321, n322, n323, n324, n325, n326, n331, n332, n333, n334, n335, 
      n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n351, 
      n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, 
      n364, n365, n366, n372, n373, n374, n375, n376, n377, n378, n379, n380, 
      n381, n382, n383, n384, n385, n386, n387, n392, n393, n394, n395, n396, 
      n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n412, 
      n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, 
      n425, n426, n427, n432, n433, n434, n435, n436, n437, n438, n439, n440, 
      n441, n442, n443, n444, n445, n446, n447, n452, n453, n454, n455, n456, 
      n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, 
      n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, 
      n481, n482, n483, n484, n485, n486, n487, n489, n494, n495, n496, n497, 
      n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, 
      n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, 
      n529, n530, n531, n532, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n558, n559, n560, 
      n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, 
      n573, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, 
      n589, n590, n591, n592, n593, n595, n600, n601, n602, n603, n604, n605, 
      n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, 
      n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, 
      n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, 
      n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, 
      n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, 
      n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n680, n681, 
      n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, 
      n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, 
      n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n720, n721, 
      n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, 
      n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, 
      n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n761, 
      n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, 
      n774, n775, n776, n781, n782, n783, n784, n785, n786, n787, n788, n789, 
      n790, n791, n792, n793, n794, n795, n796, n801, n802, n803, n804, n805, 
      n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, 
      n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, 
      n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, 
      n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n797, n798, 
      n799, n800, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, 
      n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, 
      n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, 
      n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, 
      n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, 
      n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, 
      n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, 
      n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, 
      n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, 
      n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, 
      n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, 
      n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, 
      n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, 
      n1005, n1006, n1007, n1008, n1009, n1010, sig_brt_port, n1012, n1013, 
      n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, 
      n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, 
      n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, 
      n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, 
      n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, 
      n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, 
      n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, 
      n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, 
      n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, 
      n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, 
      n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, 
      n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, 
      n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, 
      n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, 
      n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, 
      n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, 
      n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, 
      n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, 
      n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, 
      n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, 
      n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, 
      n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, 
      n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, 
      n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, 
      n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, 
      n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, 
      n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, 
      n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, 
      n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, 
      n1304, n1305, n1306, n1307, n1308 : std_logic;

begin
   sig_brt <= sig_brt_port;
   
   index_r_reg_4_inst : DLH_X1 port map( G => n1292, D => addr(6), Q => 
                           index_r_4_port);
   index_r_reg_3_inst : DLH_X1 port map( G => n1292, D => n987, Q => 
                           index_r_3_port);
   index_r_reg_2_inst : DLH_X1 port map( G => n1292, D => addr(4), Q => 
                           index_r_2_port);
   index_r_reg_1_inst : DLH_X1 port map( G => n1292, D => addr(3), Q => 
                           index_r_1_port);
   index_r_reg_0_inst : DLH_X1 port map( G => n1292, D => n888, Q => 
                           index_r_0_port);
   sig_bal_delay_reg : DFFR_X1 port map( D => n1294, CK => clk, RN => rst, Q =>
                           sig_bal_delay, QN => n856);
   opcd_delay_reg_5_inst : DFFR_X1 port map( D => opcd(5), CK => clk, RN => rst
                           , Q => opcd_delay_5_port, QN => net108096);
   opcd_delay_reg_4_inst : DFFR_X1 port map( D => opcd(4), CK => clk, RN => rst
                           , Q => opcd_delay_4_port, QN => net108095);
   opcd_delay_reg_3_inst : DFFR_X1 port map( D => opcd(3), CK => clk, RN => rst
                           , Q => opcd_delay_3_port, QN => net108094);
   opcd_delay_reg_2_inst : DFFR_X1 port map( D => opcd(2), CK => clk, RN => rst
                           , Q => opcd_delay_2_port, QN => net108093);
   opcd_delay_reg_1_inst : DFFR_X1 port map( D => opcd(1), CK => clk, RN => rst
                           , Q => net108092, QN => n214);
   opcd_delay_reg_0_inst : DFFR_X1 port map( D => opcd(0), CK => clk, RN => rst
                           , Q => net108091, QN => n219);
   index_r_delay_reg_4_inst : DFFR_X1 port map( D => index_r_4_port, CK => clk,
                           RN => rst, Q => n4, QN => n859);
   index_r_delay_reg_3_inst : DFFR_X1 port map( D => index_r_3_port, CK => clk,
                           RN => rst, Q => n8, QN => n855);
   index_r_delay_reg_2_inst : DFFR_X1 port map( D => index_r_2_port, CK => clk,
                           RN => rst, Q => n853, QN => n34);
   index_r_delay_reg_1_inst : DFFR_X1 port map( D => index_r_1_port, CK => clk,
                           RN => rst, Q => n5, QN => n858);
   index_r_delay_reg_0_inst : DFFR_X1 port map( D => index_r_0_port, CK => clk,
                           RN => rst, Q => n800, QN => n200);
   bht_reg_31_25_inst : DLH_X1 port map( G => n1290, D => n1120, Q => 
                           bht_31_25_port);
   entry_r_reg_26_inst : DLH_X1 port map( G => n962, D => N151, Q => 
                           entry_r_26_port);
   entry_r_delay_reg_26_inst : DFFR_X1 port map( D => entry_r_26_port, CK => 
                           clk, RN => rst, Q => net108090, QN => n33);
   bht_reg_0_26_inst : DLH_X1 port map( G => n1119, D => n1114, Q => 
                           bht_0_26_port);
   bht_reg_2_26_inst : DLH_X1 port map( G => n1203, D => n1114, Q => 
                           bht_2_26_port);
   bht_reg_4_26_inst : DLH_X1 port map( G => n1209, D => n1114, Q => 
                           bht_4_26_port);
   bht_reg_6_26_inst : DLH_X1 port map( G => n1215, D => n1114, Q => 
                           bht_6_26_port);
   bht_reg_8_26_inst : DLH_X1 port map( G => n1221, D => n1114, Q => 
                           bht_8_26_port);
   bht_reg_10_26_inst : DLH_X1 port map( G => n1227, D => n1114, Q => 
                           bht_10_26_port);
   bht_reg_12_26_inst : DLH_X1 port map( G => n1233, D => n1114, Q => 
                           bht_12_26_port);
   bht_reg_14_26_inst : DLH_X1 port map( G => n1239, D => n1114, Q => 
                           bht_14_26_port);
   bht_reg_16_26_inst : DLH_X1 port map( G => n1245, D => n1114, Q => 
                           bht_16_26_port);
   bht_reg_18_26_inst : DLH_X1 port map( G => n1251, D => n1114, Q => 
                           bht_18_26_port);
   bht_reg_20_26_inst : DLH_X1 port map( G => n1257, D => n1114, Q => 
                           bht_20_26_port);
   bht_reg_22_26_inst : DLH_X1 port map( G => n1263, D => n1115, Q => 
                           bht_22_26_port);
   bht_reg_24_26_inst : DLH_X1 port map( G => n1269, D => n1115, Q => 
                           bht_24_26_port);
   bht_reg_26_26_inst : DLH_X1 port map( G => n1275, D => n1115, Q => 
                           bht_26_26_port);
   bht_reg_28_26_inst : DLH_X1 port map( G => n1281, D => n1115, Q => 
                           bht_28_26_port);
   bht_reg_30_26_inst : DLH_X1 port map( G => n1287, D => n1115, Q => 
                           bht_30_26_port);
   bht_reg_31_26_inst : DLH_X1 port map( G => n1290, D => n1115, Q => 
                           bht_31_26_port);
   bht_reg_29_26_inst : DLH_X1 port map( G => n1284, D => n1115, Q => 
                           bht_29_26_port);
   bht_reg_27_26_inst : DLH_X1 port map( G => n1278, D => n1115, Q => 
                           bht_27_26_port);
   bht_reg_25_26_inst : DLH_X1 port map( G => n1272, D => n1115, Q => 
                           bht_25_26_port);
   bht_reg_23_26_inst : DLH_X1 port map( G => n1266, D => n1115, Q => 
                           bht_23_26_port);
   bht_reg_21_26_inst : DLH_X1 port map( G => n1260, D => n1115, Q => 
                           bht_21_26_port);
   bht_reg_19_26_inst : DLH_X1 port map( G => n1254, D => n1116, Q => 
                           bht_19_26_port);
   bht_reg_17_26_inst : DLH_X1 port map( G => n1248, D => n1116, Q => 
                           bht_17_26_port);
   bht_reg_15_26_inst : DLH_X1 port map( G => n1242, D => n1116, Q => 
                           bht_15_26_port);
   bht_reg_13_26_inst : DLH_X1 port map( G => n1236, D => n1116, Q => 
                           bht_13_26_port);
   bht_reg_11_26_inst : DLH_X1 port map( G => n1230, D => n1116, Q => 
                           bht_11_26_port);
   bht_reg_9_26_inst : DLH_X1 port map( G => n1224, D => n1116, Q => 
                           bht_9_26_port);
   bht_reg_7_26_inst : DLH_X1 port map( G => n1218, D => n1116, Q => 
                           bht_7_26_port);
   bht_reg_5_26_inst : DLH_X1 port map( G => n1212, D => n1116, Q => 
                           bht_5_26_port);
   bht_reg_3_26_inst : DLH_X1 port map( G => n1206, D => n1116, Q => 
                           bht_3_26_port);
   bht_reg_1_26_inst : DLH_X1 port map( G => n1200, D => n1116, Q => 
                           bht_1_26_port);
   entry_r_reg_24_inst : DLH_X1 port map( G => n962, D => N149, Q => 
                           entry_r_24_port);
   entry_r_delay_reg_24_inst : DFFR_X1 port map( D => entry_r_24_port, CK => 
                           clk, RN => rst, Q => net108089, QN => n32);
   bht_reg_0_24_inst : DLH_X1 port map( G => n1119, D => n1123, Q => 
                           bht_0_24_port);
   bht_reg_2_24_inst : DLH_X1 port map( G => n1203, D => n1123, Q => 
                           bht_2_24_port);
   bht_reg_4_24_inst : DLH_X1 port map( G => n1209, D => n1123, Q => 
                           bht_4_24_port);
   bht_reg_6_24_inst : DLH_X1 port map( G => n1215, D => n1123, Q => 
                           bht_6_24_port);
   bht_reg_8_24_inst : DLH_X1 port map( G => n1221, D => n1123, Q => 
                           bht_8_24_port);
   bht_reg_10_24_inst : DLH_X1 port map( G => n1227, D => n1123, Q => 
                           bht_10_24_port);
   bht_reg_12_24_inst : DLH_X1 port map( G => n1233, D => n1123, Q => 
                           bht_12_24_port);
   bht_reg_14_24_inst : DLH_X1 port map( G => n1239, D => n1123, Q => 
                           bht_14_24_port);
   bht_reg_16_24_inst : DLH_X1 port map( G => n1245, D => n1123, Q => 
                           bht_16_24_port);
   bht_reg_18_24_inst : DLH_X1 port map( G => n1251, D => n1123, Q => 
                           bht_18_24_port);
   bht_reg_20_24_inst : DLH_X1 port map( G => n1257, D => n1123, Q => 
                           bht_20_24_port);
   bht_reg_22_24_inst : DLH_X1 port map( G => n1263, D => n1124, Q => 
                           bht_22_24_port);
   bht_reg_24_24_inst : DLH_X1 port map( G => n1269, D => n1124, Q => 
                           bht_24_24_port);
   bht_reg_26_24_inst : DLH_X1 port map( G => n1275, D => n1124, Q => 
                           bht_26_24_port);
   bht_reg_28_24_inst : DLH_X1 port map( G => n1281, D => n1124, Q => 
                           bht_28_24_port);
   bht_reg_30_24_inst : DLH_X1 port map( G => n1287, D => n1124, Q => 
                           bht_30_24_port);
   bht_reg_31_24_inst : DLH_X1 port map( G => n1290, D => n1124, Q => 
                           bht_31_24_port);
   bht_reg_29_24_inst : DLH_X1 port map( G => n1284, D => n1124, Q => 
                           bht_29_24_port);
   bht_reg_27_24_inst : DLH_X1 port map( G => n1278, D => n1124, Q => 
                           bht_27_24_port);
   bht_reg_25_24_inst : DLH_X1 port map( G => n1272, D => n1124, Q => 
                           bht_25_24_port);
   bht_reg_23_24_inst : DLH_X1 port map( G => n1266, D => n1124, Q => 
                           bht_23_24_port);
   bht_reg_21_24_inst : DLH_X1 port map( G => n1260, D => n1124, Q => 
                           bht_21_24_port);
   bht_reg_19_24_inst : DLH_X1 port map( G => n1254, D => n1125, Q => 
                           bht_19_24_port);
   bht_reg_17_24_inst : DLH_X1 port map( G => n1248, D => n1125, Q => 
                           bht_17_24_port);
   bht_reg_15_24_inst : DLH_X1 port map( G => n1242, D => n1125, Q => 
                           bht_15_24_port);
   bht_reg_13_24_inst : DLH_X1 port map( G => n1236, D => n1125, Q => 
                           bht_13_24_port);
   bht_reg_11_24_inst : DLH_X1 port map( G => n1230, D => n1125, Q => 
                           bht_11_24_port);
   bht_reg_9_24_inst : DLH_X1 port map( G => n1224, D => n1125, Q => 
                           bht_9_24_port);
   bht_reg_7_24_inst : DLH_X1 port map( G => n1218, D => n1125, Q => 
                           bht_7_24_port);
   bht_reg_5_24_inst : DLH_X1 port map( G => n1212, D => n1125, Q => 
                           bht_5_24_port);
   bht_reg_3_24_inst : DLH_X1 port map( G => n1206, D => n1125, Q => 
                           bht_3_24_port);
   bht_reg_1_24_inst : DLH_X1 port map( G => n1200, D => n1125, Q => 
                           bht_1_24_port);
   entry_r_reg_23_inst : DLH_X1 port map( G => n962, D => N148, Q => 
                           entry_r_23_port);
   entry_r_delay_reg_23_inst : DFFR_X1 port map( D => entry_r_23_port, CK => 
                           clk, RN => rst, Q => net108088, QN => n31);
   bht_reg_0_23_inst : DLH_X1 port map( G => n1119, D => n1126, Q => 
                           bht_0_23_port);
   bht_reg_2_23_inst : DLH_X1 port map( G => n1203, D => n1126, Q => 
                           bht_2_23_port);
   bht_reg_4_23_inst : DLH_X1 port map( G => n1209, D => n1126, Q => 
                           bht_4_23_port);
   bht_reg_6_23_inst : DLH_X1 port map( G => n1215, D => n1126, Q => 
                           bht_6_23_port);
   bht_reg_8_23_inst : DLH_X1 port map( G => n1221, D => n1126, Q => 
                           bht_8_23_port);
   bht_reg_10_23_inst : DLH_X1 port map( G => n1227, D => n1126, Q => 
                           bht_10_23_port);
   bht_reg_12_23_inst : DLH_X1 port map( G => n1233, D => n1126, Q => 
                           bht_12_23_port);
   bht_reg_14_23_inst : DLH_X1 port map( G => n1239, D => n1126, Q => 
                           bht_14_23_port);
   bht_reg_16_23_inst : DLH_X1 port map( G => n1245, D => n1126, Q => 
                           bht_16_23_port);
   bht_reg_18_23_inst : DLH_X1 port map( G => n1251, D => n1126, Q => 
                           bht_18_23_port);
   bht_reg_20_23_inst : DLH_X1 port map( G => n1257, D => n1126, Q => 
                           bht_20_23_port);
   bht_reg_22_23_inst : DLH_X1 port map( G => n1263, D => n1127, Q => 
                           bht_22_23_port);
   bht_reg_24_23_inst : DLH_X1 port map( G => n1269, D => n1127, Q => 
                           bht_24_23_port);
   bht_reg_26_23_inst : DLH_X1 port map( G => n1275, D => n1127, Q => 
                           bht_26_23_port);
   bht_reg_28_23_inst : DLH_X1 port map( G => n1281, D => n1127, Q => 
                           bht_28_23_port);
   bht_reg_30_23_inst : DLH_X1 port map( G => n1287, D => n1127, Q => 
                           bht_30_23_port);
   bht_reg_31_23_inst : DLH_X1 port map( G => n1290, D => n1127, Q => 
                           bht_31_23_port);
   bht_reg_29_23_inst : DLH_X1 port map( G => n1284, D => n1127, Q => 
                           bht_29_23_port);
   bht_reg_27_23_inst : DLH_X1 port map( G => n1278, D => n1127, Q => 
                           bht_27_23_port);
   bht_reg_25_23_inst : DLH_X1 port map( G => n1272, D => n1127, Q => 
                           bht_25_23_port);
   bht_reg_23_23_inst : DLH_X1 port map( G => n1266, D => n1127, Q => 
                           bht_23_23_port);
   bht_reg_21_23_inst : DLH_X1 port map( G => n1260, D => n1127, Q => 
                           bht_21_23_port);
   bht_reg_19_23_inst : DLH_X1 port map( G => n1254, D => n1128, Q => 
                           bht_19_23_port);
   bht_reg_17_23_inst : DLH_X1 port map( G => n1248, D => n1128, Q => 
                           bht_17_23_port);
   bht_reg_15_23_inst : DLH_X1 port map( G => n1242, D => n1128, Q => 
                           bht_15_23_port);
   bht_reg_13_23_inst : DLH_X1 port map( G => n1236, D => n1128, Q => 
                           bht_13_23_port);
   bht_reg_11_23_inst : DLH_X1 port map( G => n1230, D => n1128, Q => 
                           bht_11_23_port);
   bht_reg_9_23_inst : DLH_X1 port map( G => n1224, D => n1128, Q => 
                           bht_9_23_port);
   bht_reg_7_23_inst : DLH_X1 port map( G => n1218, D => n1128, Q => 
                           bht_7_23_port);
   bht_reg_5_23_inst : DLH_X1 port map( G => n1212, D => n1128, Q => 
                           bht_5_23_port);
   bht_reg_3_23_inst : DLH_X1 port map( G => n1206, D => n1128, Q => 
                           bht_3_23_port);
   bht_reg_1_23_inst : DLH_X1 port map( G => n1200, D => n1128, Q => 
                           bht_1_23_port);
   entry_r_reg_22_inst : DLH_X1 port map( G => n962, D => N147, Q => 
                           entry_r_22_port);
   entry_r_delay_reg_22_inst : DFFR_X1 port map( D => entry_r_22_port, CK => 
                           clk, RN => rst, Q => net108087, QN => n30);
   bht_reg_0_22_inst : DLH_X1 port map( G => n1119, D => n1129, Q => 
                           bht_0_22_port);
   bht_reg_2_22_inst : DLH_X1 port map( G => n1203, D => n1129, Q => 
                           bht_2_22_port);
   bht_reg_4_22_inst : DLH_X1 port map( G => n1209, D => n1129, Q => 
                           bht_4_22_port);
   bht_reg_6_22_inst : DLH_X1 port map( G => n1215, D => n1129, Q => 
                           bht_6_22_port);
   bht_reg_8_22_inst : DLH_X1 port map( G => n1221, D => n1129, Q => 
                           bht_8_22_port);
   bht_reg_10_22_inst : DLH_X1 port map( G => n1227, D => n1129, Q => 
                           bht_10_22_port);
   bht_reg_12_22_inst : DLH_X1 port map( G => n1233, D => n1129, Q => 
                           bht_12_22_port);
   bht_reg_14_22_inst : DLH_X1 port map( G => n1239, D => n1129, Q => 
                           bht_14_22_port);
   bht_reg_16_22_inst : DLH_X1 port map( G => n1245, D => n1129, Q => 
                           bht_16_22_port);
   bht_reg_18_22_inst : DLH_X1 port map( G => n1251, D => n1129, Q => 
                           bht_18_22_port);
   bht_reg_20_22_inst : DLH_X1 port map( G => n1257, D => n1129, Q => 
                           bht_20_22_port);
   bht_reg_22_22_inst : DLH_X1 port map( G => n1263, D => n1130, Q => 
                           bht_22_22_port);
   bht_reg_24_22_inst : DLH_X1 port map( G => n1269, D => n1130, Q => 
                           bht_24_22_port);
   bht_reg_26_22_inst : DLH_X1 port map( G => n1275, D => n1130, Q => 
                           bht_26_22_port);
   bht_reg_28_22_inst : DLH_X1 port map( G => n1281, D => n1130, Q => 
                           bht_28_22_port);
   bht_reg_30_22_inst : DLH_X1 port map( G => n1287, D => n1130, Q => 
                           bht_30_22_port);
   bht_reg_31_22_inst : DLH_X1 port map( G => n1290, D => n1130, Q => 
                           bht_31_22_port);
   bht_reg_29_22_inst : DLH_X1 port map( G => n1284, D => n1130, Q => 
                           bht_29_22_port);
   bht_reg_27_22_inst : DLH_X1 port map( G => n1278, D => n1130, Q => 
                           bht_27_22_port);
   bht_reg_25_22_inst : DLH_X1 port map( G => n1272, D => n1130, Q => 
                           bht_25_22_port);
   bht_reg_23_22_inst : DLH_X1 port map( G => n1266, D => n1130, Q => 
                           bht_23_22_port);
   bht_reg_21_22_inst : DLH_X1 port map( G => n1260, D => n1130, Q => 
                           bht_21_22_port);
   bht_reg_19_22_inst : DLH_X1 port map( G => n1254, D => n1131, Q => 
                           bht_19_22_port);
   bht_reg_17_22_inst : DLH_X1 port map( G => n1248, D => n1131, Q => 
                           bht_17_22_port);
   bht_reg_15_22_inst : DLH_X1 port map( G => n1242, D => n1131, Q => 
                           bht_15_22_port);
   bht_reg_13_22_inst : DLH_X1 port map( G => n1236, D => n1131, Q => 
                           bht_13_22_port);
   bht_reg_11_22_inst : DLH_X1 port map( G => n1230, D => n1131, Q => 
                           bht_11_22_port);
   bht_reg_9_22_inst : DLH_X1 port map( G => n1224, D => n1131, Q => 
                           bht_9_22_port);
   bht_reg_7_22_inst : DLH_X1 port map( G => n1218, D => n1131, Q => 
                           bht_7_22_port);
   bht_reg_5_22_inst : DLH_X1 port map( G => n1212, D => n1131, Q => 
                           bht_5_22_port);
   bht_reg_3_22_inst : DLH_X1 port map( G => n1206, D => n1131, Q => 
                           bht_3_22_port);
   bht_reg_1_22_inst : DLH_X1 port map( G => n1200, D => n1131, Q => 
                           bht_1_22_port);
   entry_r_reg_21_inst : DLH_X1 port map( G => n962, D => N146, Q => 
                           entry_r_21_port);
   entry_r_delay_reg_21_inst : DFFR_X1 port map( D => entry_r_21_port, CK => 
                           clk, RN => rst, Q => net108086, QN => n29);
   bht_reg_0_21_inst : DLH_X1 port map( G => n1118, D => n1132, Q => 
                           bht_0_21_port);
   bht_reg_2_21_inst : DLH_X1 port map( G => n1202, D => n1132, Q => 
                           bht_2_21_port);
   bht_reg_4_21_inst : DLH_X1 port map( G => n1208, D => n1132, Q => 
                           bht_4_21_port);
   bht_reg_6_21_inst : DLH_X1 port map( G => n1214, D => n1132, Q => 
                           bht_6_21_port);
   bht_reg_8_21_inst : DLH_X1 port map( G => n1220, D => n1132, Q => 
                           bht_8_21_port);
   bht_reg_10_21_inst : DLH_X1 port map( G => n1226, D => n1132, Q => 
                           bht_10_21_port);
   bht_reg_12_21_inst : DLH_X1 port map( G => n1232, D => n1132, Q => 
                           bht_12_21_port);
   bht_reg_14_21_inst : DLH_X1 port map( G => n1238, D => n1132, Q => 
                           bht_14_21_port);
   bht_reg_16_21_inst : DLH_X1 port map( G => n1244, D => n1132, Q => 
                           bht_16_21_port);
   bht_reg_18_21_inst : DLH_X1 port map( G => n1250, D => n1132, Q => 
                           bht_18_21_port);
   bht_reg_20_21_inst : DLH_X1 port map( G => n1256, D => n1132, Q => 
                           bht_20_21_port);
   bht_reg_22_21_inst : DLH_X1 port map( G => n1262, D => n1133, Q => 
                           bht_22_21_port);
   bht_reg_24_21_inst : DLH_X1 port map( G => n1268, D => n1133, Q => 
                           bht_24_21_port);
   bht_reg_26_21_inst : DLH_X1 port map( G => n1274, D => n1133, Q => 
                           bht_26_21_port);
   bht_reg_28_21_inst : DLH_X1 port map( G => n1280, D => n1133, Q => 
                           bht_28_21_port);
   bht_reg_30_21_inst : DLH_X1 port map( G => n1286, D => n1133, Q => 
                           bht_30_21_port);
   bht_reg_31_21_inst : DLH_X1 port map( G => n1289, D => n1133, Q => 
                           bht_31_21_port);
   bht_reg_29_21_inst : DLH_X1 port map( G => n1283, D => n1133, Q => 
                           bht_29_21_port);
   bht_reg_27_21_inst : DLH_X1 port map( G => n1277, D => n1133, Q => 
                           bht_27_21_port);
   bht_reg_25_21_inst : DLH_X1 port map( G => n1271, D => n1133, Q => 
                           bht_25_21_port);
   bht_reg_23_21_inst : DLH_X1 port map( G => n1265, D => n1133, Q => 
                           bht_23_21_port);
   bht_reg_21_21_inst : DLH_X1 port map( G => n1259, D => n1133, Q => 
                           bht_21_21_port);
   bht_reg_19_21_inst : DLH_X1 port map( G => n1253, D => n1134, Q => 
                           bht_19_21_port);
   bht_reg_17_21_inst : DLH_X1 port map( G => n1247, D => n1134, Q => 
                           bht_17_21_port);
   bht_reg_15_21_inst : DLH_X1 port map( G => n1241, D => n1134, Q => 
                           bht_15_21_port);
   bht_reg_13_21_inst : DLH_X1 port map( G => n1235, D => n1134, Q => 
                           bht_13_21_port);
   bht_reg_11_21_inst : DLH_X1 port map( G => n1229, D => n1134, Q => 
                           bht_11_21_port);
   bht_reg_9_21_inst : DLH_X1 port map( G => n1223, D => n1134, Q => 
                           bht_9_21_port);
   bht_reg_7_21_inst : DLH_X1 port map( G => n1217, D => n1134, Q => 
                           bht_7_21_port);
   bht_reg_5_21_inst : DLH_X1 port map( G => n1211, D => n1134, Q => 
                           bht_5_21_port);
   bht_reg_3_21_inst : DLH_X1 port map( G => n1205, D => n1134, Q => 
                           bht_3_21_port);
   bht_reg_1_21_inst : DLH_X1 port map( G => n1199, D => n1134, Q => 
                           bht_1_21_port);
   entry_r_reg_20_inst : DLH_X1 port map( G => n962, D => N145, Q => 
                           entry_r_20_port);
   entry_r_delay_reg_20_inst : DFFR_X1 port map( D => entry_r_20_port, CK => 
                           clk, RN => rst, Q => net108085, QN => n28);
   bht_reg_0_20_inst : DLH_X1 port map( G => n1118, D => n1135, Q => 
                           bht_0_20_port);
   bht_reg_2_20_inst : DLH_X1 port map( G => n1202, D => n1135, Q => 
                           bht_2_20_port);
   bht_reg_4_20_inst : DLH_X1 port map( G => n1208, D => n1135, Q => 
                           bht_4_20_port);
   bht_reg_6_20_inst : DLH_X1 port map( G => n1214, D => n1135, Q => 
                           bht_6_20_port);
   bht_reg_8_20_inst : DLH_X1 port map( G => n1220, D => n1135, Q => 
                           bht_8_20_port);
   bht_reg_10_20_inst : DLH_X1 port map( G => n1226, D => n1135, Q => 
                           bht_10_20_port);
   bht_reg_12_20_inst : DLH_X1 port map( G => n1232, D => n1135, Q => 
                           bht_12_20_port);
   bht_reg_14_20_inst : DLH_X1 port map( G => n1238, D => n1135, Q => 
                           bht_14_20_port);
   bht_reg_16_20_inst : DLH_X1 port map( G => n1244, D => n1135, Q => 
                           bht_16_20_port);
   bht_reg_18_20_inst : DLH_X1 port map( G => n1250, D => n1135, Q => 
                           bht_18_20_port);
   bht_reg_20_20_inst : DLH_X1 port map( G => n1256, D => n1135, Q => 
                           bht_20_20_port);
   bht_reg_22_20_inst : DLH_X1 port map( G => n1262, D => n1136, Q => 
                           bht_22_20_port);
   bht_reg_24_20_inst : DLH_X1 port map( G => n1268, D => n1136, Q => 
                           bht_24_20_port);
   bht_reg_26_20_inst : DLH_X1 port map( G => n1274, D => n1136, Q => 
                           bht_26_20_port);
   bht_reg_28_20_inst : DLH_X1 port map( G => n1280, D => n1136, Q => 
                           bht_28_20_port);
   bht_reg_30_20_inst : DLH_X1 port map( G => n1286, D => n1136, Q => 
                           bht_30_20_port);
   bht_reg_31_20_inst : DLH_X1 port map( G => n1289, D => n1136, Q => 
                           bht_31_20_port);
   bht_reg_29_20_inst : DLH_X1 port map( G => n1283, D => n1136, Q => 
                           bht_29_20_port);
   bht_reg_27_20_inst : DLH_X1 port map( G => n1277, D => n1136, Q => 
                           bht_27_20_port);
   bht_reg_25_20_inst : DLH_X1 port map( G => n1271, D => n1136, Q => 
                           bht_25_20_port);
   bht_reg_23_20_inst : DLH_X1 port map( G => n1265, D => n1136, Q => 
                           bht_23_20_port);
   bht_reg_21_20_inst : DLH_X1 port map( G => n1259, D => n1136, Q => 
                           bht_21_20_port);
   bht_reg_19_20_inst : DLH_X1 port map( G => n1253, D => n1137, Q => 
                           bht_19_20_port);
   bht_reg_17_20_inst : DLH_X1 port map( G => n1247, D => n1137, Q => 
                           bht_17_20_port);
   bht_reg_15_20_inst : DLH_X1 port map( G => n1241, D => n1137, Q => 
                           bht_15_20_port);
   bht_reg_13_20_inst : DLH_X1 port map( G => n1235, D => n1137, Q => 
                           bht_13_20_port);
   bht_reg_11_20_inst : DLH_X1 port map( G => n1229, D => n1137, Q => 
                           bht_11_20_port);
   bht_reg_9_20_inst : DLH_X1 port map( G => n1223, D => n1137, Q => 
                           bht_9_20_port);
   bht_reg_7_20_inst : DLH_X1 port map( G => n1217, D => n1137, Q => 
                           bht_7_20_port);
   bht_reg_5_20_inst : DLH_X1 port map( G => n1211, D => n1137, Q => 
                           bht_5_20_port);
   bht_reg_3_20_inst : DLH_X1 port map( G => n1205, D => n1137, Q => 
                           bht_3_20_port);
   bht_reg_1_20_inst : DLH_X1 port map( G => n1199, D => n1137, Q => 
                           bht_1_20_port);
   entry_r_reg_19_inst : DLH_X1 port map( G => n962, D => N144, Q => 
                           entry_r_19_port);
   entry_r_delay_reg_19_inst : DFFR_X1 port map( D => entry_r_19_port, CK => 
                           clk, RN => rst, Q => net108084, QN => n27);
   bht_reg_0_19_inst : DLH_X1 port map( G => n1118, D => n1138, Q => 
                           bht_0_19_port);
   bht_reg_2_19_inst : DLH_X1 port map( G => n1202, D => n1138, Q => 
                           bht_2_19_port);
   bht_reg_4_19_inst : DLH_X1 port map( G => n1208, D => n1138, Q => 
                           bht_4_19_port);
   bht_reg_6_19_inst : DLH_X1 port map( G => n1214, D => n1138, Q => 
                           bht_6_19_port);
   bht_reg_8_19_inst : DLH_X1 port map( G => n1220, D => n1138, Q => 
                           bht_8_19_port);
   bht_reg_10_19_inst : DLH_X1 port map( G => n1226, D => n1138, Q => 
                           bht_10_19_port);
   bht_reg_12_19_inst : DLH_X1 port map( G => n1232, D => n1138, Q => 
                           bht_12_19_port);
   bht_reg_14_19_inst : DLH_X1 port map( G => n1238, D => n1138, Q => 
                           bht_14_19_port);
   bht_reg_16_19_inst : DLH_X1 port map( G => n1244, D => n1138, Q => 
                           bht_16_19_port);
   bht_reg_18_19_inst : DLH_X1 port map( G => n1250, D => n1138, Q => 
                           bht_18_19_port);
   bht_reg_20_19_inst : DLH_X1 port map( G => n1256, D => n1138, Q => 
                           bht_20_19_port);
   bht_reg_22_19_inst : DLH_X1 port map( G => n1262, D => n1139, Q => 
                           bht_22_19_port);
   bht_reg_24_19_inst : DLH_X1 port map( G => n1268, D => n1139, Q => 
                           bht_24_19_port);
   bht_reg_26_19_inst : DLH_X1 port map( G => n1274, D => n1139, Q => 
                           bht_26_19_port);
   bht_reg_28_19_inst : DLH_X1 port map( G => n1280, D => n1139, Q => 
                           bht_28_19_port);
   bht_reg_30_19_inst : DLH_X1 port map( G => n1286, D => n1139, Q => 
                           bht_30_19_port);
   bht_reg_31_19_inst : DLH_X1 port map( G => n1289, D => n1139, Q => 
                           bht_31_19_port);
   bht_reg_29_19_inst : DLH_X1 port map( G => n1283, D => n1139, Q => 
                           bht_29_19_port);
   bht_reg_27_19_inst : DLH_X1 port map( G => n1277, D => n1139, Q => 
                           bht_27_19_port);
   bht_reg_25_19_inst : DLH_X1 port map( G => n1271, D => n1139, Q => 
                           bht_25_19_port);
   bht_reg_23_19_inst : DLH_X1 port map( G => n1265, D => n1139, Q => 
                           bht_23_19_port);
   bht_reg_21_19_inst : DLH_X1 port map( G => n1259, D => n1139, Q => 
                           bht_21_19_port);
   bht_reg_19_19_inst : DLH_X1 port map( G => n1253, D => n1140, Q => 
                           bht_19_19_port);
   bht_reg_17_19_inst : DLH_X1 port map( G => n1247, D => n1140, Q => 
                           bht_17_19_port);
   bht_reg_15_19_inst : DLH_X1 port map( G => n1241, D => n1140, Q => 
                           bht_15_19_port);
   bht_reg_13_19_inst : DLH_X1 port map( G => n1235, D => n1140, Q => 
                           bht_13_19_port);
   bht_reg_11_19_inst : DLH_X1 port map( G => n1229, D => n1140, Q => 
                           bht_11_19_port);
   bht_reg_9_19_inst : DLH_X1 port map( G => n1223, D => n1140, Q => 
                           bht_9_19_port);
   bht_reg_7_19_inst : DLH_X1 port map( G => n1217, D => n1140, Q => 
                           bht_7_19_port);
   bht_reg_5_19_inst : DLH_X1 port map( G => n1211, D => n1140, Q => 
                           bht_5_19_port);
   bht_reg_3_19_inst : DLH_X1 port map( G => n1205, D => n1140, Q => 
                           bht_3_19_port);
   bht_reg_1_19_inst : DLH_X1 port map( G => n1199, D => n1140, Q => 
                           bht_1_19_port);
   entry_r_reg_18_inst : DLH_X1 port map( G => n962, D => N143, Q => 
                           entry_r_18_port);
   entry_r_delay_reg_18_inst : DFFR_X1 port map( D => entry_r_18_port, CK => 
                           clk, RN => rst, Q => net108083, QN => n26);
   bht_reg_0_18_inst : DLH_X1 port map( G => n1118, D => n1141, Q => 
                           bht_0_18_port);
   bht_reg_2_18_inst : DLH_X1 port map( G => n1202, D => n1141, Q => 
                           bht_2_18_port);
   bht_reg_4_18_inst : DLH_X1 port map( G => n1208, D => n1141, Q => 
                           bht_4_18_port);
   bht_reg_6_18_inst : DLH_X1 port map( G => n1214, D => n1141, Q => 
                           bht_6_18_port);
   bht_reg_8_18_inst : DLH_X1 port map( G => n1220, D => n1141, Q => 
                           bht_8_18_port);
   bht_reg_10_18_inst : DLH_X1 port map( G => n1226, D => n1141, Q => 
                           bht_10_18_port);
   bht_reg_12_18_inst : DLH_X1 port map( G => n1232, D => n1141, Q => 
                           bht_12_18_port);
   bht_reg_14_18_inst : DLH_X1 port map( G => n1238, D => n1141, Q => 
                           bht_14_18_port);
   bht_reg_16_18_inst : DLH_X1 port map( G => n1244, D => n1141, Q => 
                           bht_16_18_port);
   bht_reg_18_18_inst : DLH_X1 port map( G => n1250, D => n1141, Q => 
                           bht_18_18_port);
   bht_reg_20_18_inst : DLH_X1 port map( G => n1256, D => n1141, Q => 
                           bht_20_18_port);
   bht_reg_22_18_inst : DLH_X1 port map( G => n1262, D => n1142, Q => 
                           bht_22_18_port);
   bht_reg_24_18_inst : DLH_X1 port map( G => n1268, D => n1142, Q => 
                           bht_24_18_port);
   bht_reg_26_18_inst : DLH_X1 port map( G => n1274, D => n1142, Q => 
                           bht_26_18_port);
   bht_reg_28_18_inst : DLH_X1 port map( G => n1280, D => n1142, Q => 
                           bht_28_18_port);
   bht_reg_30_18_inst : DLH_X1 port map( G => n1286, D => n1142, Q => 
                           bht_30_18_port);
   bht_reg_31_18_inst : DLH_X1 port map( G => n1289, D => n1142, Q => 
                           bht_31_18_port);
   bht_reg_29_18_inst : DLH_X1 port map( G => n1283, D => n1142, Q => 
                           bht_29_18_port);
   bht_reg_27_18_inst : DLH_X1 port map( G => n1277, D => n1142, Q => 
                           bht_27_18_port);
   bht_reg_25_18_inst : DLH_X1 port map( G => n1271, D => n1142, Q => 
                           bht_25_18_port);
   bht_reg_23_18_inst : DLH_X1 port map( G => n1265, D => n1142, Q => 
                           bht_23_18_port);
   bht_reg_21_18_inst : DLH_X1 port map( G => n1259, D => n1142, Q => 
                           bht_21_18_port);
   bht_reg_19_18_inst : DLH_X1 port map( G => n1253, D => n1143, Q => 
                           bht_19_18_port);
   bht_reg_17_18_inst : DLH_X1 port map( G => n1247, D => n1143, Q => 
                           bht_17_18_port);
   bht_reg_15_18_inst : DLH_X1 port map( G => n1241, D => n1143, Q => 
                           bht_15_18_port);
   bht_reg_13_18_inst : DLH_X1 port map( G => n1235, D => n1143, Q => 
                           bht_13_18_port);
   bht_reg_11_18_inst : DLH_X1 port map( G => n1229, D => n1143, Q => 
                           bht_11_18_port);
   bht_reg_9_18_inst : DLH_X1 port map( G => n1223, D => n1143, Q => 
                           bht_9_18_port);
   bht_reg_7_18_inst : DLH_X1 port map( G => n1217, D => n1143, Q => 
                           bht_7_18_port);
   bht_reg_5_18_inst : DLH_X1 port map( G => n1211, D => n1143, Q => 
                           bht_5_18_port);
   bht_reg_3_18_inst : DLH_X1 port map( G => n1205, D => n1143, Q => 
                           bht_3_18_port);
   bht_reg_1_18_inst : DLH_X1 port map( G => n1199, D => n1143, Q => 
                           bht_1_18_port);
   entry_r_reg_17_inst : DLH_X1 port map( G => n962, D => N142, Q => 
                           entry_r_17_port);
   entry_r_delay_reg_17_inst : DFFR_X1 port map( D => entry_r_17_port, CK => 
                           clk, RN => rst, Q => net108082, QN => n25);
   bht_reg_0_17_inst : DLH_X1 port map( G => n1118, D => n1144, Q => 
                           bht_0_17_port);
   bht_reg_2_17_inst : DLH_X1 port map( G => n1202, D => n1144, Q => 
                           bht_2_17_port);
   bht_reg_4_17_inst : DLH_X1 port map( G => n1208, D => n1144, Q => 
                           bht_4_17_port);
   bht_reg_6_17_inst : DLH_X1 port map( G => n1214, D => n1144, Q => 
                           bht_6_17_port);
   bht_reg_8_17_inst : DLH_X1 port map( G => n1220, D => n1144, Q => 
                           bht_8_17_port);
   bht_reg_10_17_inst : DLH_X1 port map( G => n1226, D => n1144, Q => 
                           bht_10_17_port);
   bht_reg_12_17_inst : DLH_X1 port map( G => n1232, D => n1144, Q => 
                           bht_12_17_port);
   bht_reg_14_17_inst : DLH_X1 port map( G => n1238, D => n1144, Q => 
                           bht_14_17_port);
   bht_reg_16_17_inst : DLH_X1 port map( G => n1244, D => n1144, Q => 
                           bht_16_17_port);
   bht_reg_18_17_inst : DLH_X1 port map( G => n1250, D => n1144, Q => 
                           bht_18_17_port);
   bht_reg_20_17_inst : DLH_X1 port map( G => n1256, D => n1144, Q => 
                           bht_20_17_port);
   bht_reg_22_17_inst : DLH_X1 port map( G => n1262, D => n1145, Q => 
                           bht_22_17_port);
   bht_reg_24_17_inst : DLH_X1 port map( G => n1268, D => n1145, Q => 
                           bht_24_17_port);
   bht_reg_26_17_inst : DLH_X1 port map( G => n1274, D => n1145, Q => 
                           bht_26_17_port);
   bht_reg_28_17_inst : DLH_X1 port map( G => n1280, D => n1145, Q => 
                           bht_28_17_port);
   bht_reg_30_17_inst : DLH_X1 port map( G => n1286, D => n1145, Q => 
                           bht_30_17_port);
   bht_reg_31_17_inst : DLH_X1 port map( G => n1289, D => n1145, Q => 
                           bht_31_17_port);
   bht_reg_29_17_inst : DLH_X1 port map( G => n1283, D => n1145, Q => 
                           bht_29_17_port);
   bht_reg_27_17_inst : DLH_X1 port map( G => n1277, D => n1145, Q => 
                           bht_27_17_port);
   bht_reg_25_17_inst : DLH_X1 port map( G => n1271, D => n1145, Q => 
                           bht_25_17_port);
   bht_reg_23_17_inst : DLH_X1 port map( G => n1265, D => n1145, Q => 
                           bht_23_17_port);
   bht_reg_21_17_inst : DLH_X1 port map( G => n1259, D => n1145, Q => 
                           bht_21_17_port);
   bht_reg_19_17_inst : DLH_X1 port map( G => n1253, D => n1146, Q => 
                           bht_19_17_port);
   bht_reg_17_17_inst : DLH_X1 port map( G => n1247, D => n1146, Q => 
                           bht_17_17_port);
   bht_reg_15_17_inst : DLH_X1 port map( G => n1241, D => n1146, Q => 
                           bht_15_17_port);
   bht_reg_13_17_inst : DLH_X1 port map( G => n1235, D => n1146, Q => 
                           bht_13_17_port);
   bht_reg_11_17_inst : DLH_X1 port map( G => n1229, D => n1146, Q => 
                           bht_11_17_port);
   bht_reg_9_17_inst : DLH_X1 port map( G => n1223, D => n1146, Q => 
                           bht_9_17_port);
   bht_reg_7_17_inst : DLH_X1 port map( G => n1217, D => n1146, Q => 
                           bht_7_17_port);
   bht_reg_5_17_inst : DLH_X1 port map( G => n1211, D => n1146, Q => 
                           bht_5_17_port);
   bht_reg_3_17_inst : DLH_X1 port map( G => n1205, D => n1146, Q => 
                           bht_3_17_port);
   bht_reg_1_17_inst : DLH_X1 port map( G => n1199, D => n1146, Q => 
                           bht_1_17_port);
   entry_r_reg_16_inst : DLH_X1 port map( G => n962, D => N141, Q => 
                           entry_r_16_port);
   entry_r_delay_reg_16_inst : DFFR_X1 port map( D => entry_r_16_port, CK => 
                           clk, RN => rst, Q => net108081, QN => n24);
   bht_reg_0_16_inst : DLH_X1 port map( G => n1118, D => n1147, Q => 
                           bht_0_16_port);
   bht_reg_2_16_inst : DLH_X1 port map( G => n1202, D => n1147, Q => 
                           bht_2_16_port);
   bht_reg_4_16_inst : DLH_X1 port map( G => n1208, D => n1147, Q => 
                           bht_4_16_port);
   bht_reg_6_16_inst : DLH_X1 port map( G => n1214, D => n1147, Q => 
                           bht_6_16_port);
   bht_reg_8_16_inst : DLH_X1 port map( G => n1220, D => n1147, Q => 
                           bht_8_16_port);
   bht_reg_10_16_inst : DLH_X1 port map( G => n1226, D => n1147, Q => 
                           bht_10_16_port);
   bht_reg_12_16_inst : DLH_X1 port map( G => n1232, D => n1147, Q => 
                           bht_12_16_port);
   bht_reg_14_16_inst : DLH_X1 port map( G => n1238, D => n1147, Q => 
                           bht_14_16_port);
   bht_reg_16_16_inst : DLH_X1 port map( G => n1244, D => n1147, Q => 
                           bht_16_16_port);
   bht_reg_18_16_inst : DLH_X1 port map( G => n1250, D => n1147, Q => 
                           bht_18_16_port);
   bht_reg_20_16_inst : DLH_X1 port map( G => n1256, D => n1147, Q => 
                           bht_20_16_port);
   bht_reg_22_16_inst : DLH_X1 port map( G => n1262, D => n1148, Q => 
                           bht_22_16_port);
   bht_reg_24_16_inst : DLH_X1 port map( G => n1268, D => n1148, Q => 
                           bht_24_16_port);
   bht_reg_26_16_inst : DLH_X1 port map( G => n1274, D => n1148, Q => 
                           bht_26_16_port);
   bht_reg_28_16_inst : DLH_X1 port map( G => n1280, D => n1148, Q => 
                           bht_28_16_port);
   bht_reg_30_16_inst : DLH_X1 port map( G => n1286, D => n1148, Q => 
                           bht_30_16_port);
   bht_reg_31_16_inst : DLH_X1 port map( G => n1289, D => n1148, Q => 
                           bht_31_16_port);
   bht_reg_29_16_inst : DLH_X1 port map( G => n1283, D => n1148, Q => 
                           bht_29_16_port);
   bht_reg_27_16_inst : DLH_X1 port map( G => n1277, D => n1148, Q => 
                           bht_27_16_port);
   bht_reg_25_16_inst : DLH_X1 port map( G => n1271, D => n1148, Q => 
                           bht_25_16_port);
   bht_reg_23_16_inst : DLH_X1 port map( G => n1265, D => n1148, Q => 
                           bht_23_16_port);
   bht_reg_21_16_inst : DLH_X1 port map( G => n1259, D => n1148, Q => 
                           bht_21_16_port);
   bht_reg_19_16_inst : DLH_X1 port map( G => n1253, D => n1149, Q => 
                           bht_19_16_port);
   bht_reg_17_16_inst : DLH_X1 port map( G => n1247, D => n1149, Q => 
                           bht_17_16_port);
   bht_reg_15_16_inst : DLH_X1 port map( G => n1241, D => n1149, Q => 
                           bht_15_16_port);
   bht_reg_13_16_inst : DLH_X1 port map( G => n1235, D => n1149, Q => 
                           bht_13_16_port);
   bht_reg_11_16_inst : DLH_X1 port map( G => n1229, D => n1149, Q => 
                           bht_11_16_port);
   bht_reg_9_16_inst : DLH_X1 port map( G => n1223, D => n1149, Q => 
                           bht_9_16_port);
   bht_reg_7_16_inst : DLH_X1 port map( G => n1217, D => n1149, Q => 
                           bht_7_16_port);
   bht_reg_5_16_inst : DLH_X1 port map( G => n1211, D => n1149, Q => 
                           bht_5_16_port);
   bht_reg_3_16_inst : DLH_X1 port map( G => n1205, D => n1149, Q => 
                           bht_3_16_port);
   bht_reg_1_16_inst : DLH_X1 port map( G => n1199, D => n1149, Q => 
                           bht_1_16_port);
   entry_r_reg_15_inst : DLH_X1 port map( G => n961, D => N140, Q => 
                           entry_r_15_port);
   entry_r_delay_reg_15_inst : DFFR_X1 port map( D => entry_r_15_port, CK => 
                           clk, RN => rst, Q => net108080, QN => n23);
   bht_reg_0_15_inst : DLH_X1 port map( G => n1118, D => n1150, Q => 
                           bht_0_15_port);
   bht_reg_2_15_inst : DLH_X1 port map( G => n1202, D => n1150, Q => 
                           bht_2_15_port);
   bht_reg_4_15_inst : DLH_X1 port map( G => n1208, D => n1150, Q => 
                           bht_4_15_port);
   bht_reg_6_15_inst : DLH_X1 port map( G => n1214, D => n1150, Q => 
                           bht_6_15_port);
   bht_reg_8_15_inst : DLH_X1 port map( G => n1220, D => n1150, Q => 
                           bht_8_15_port);
   bht_reg_10_15_inst : DLH_X1 port map( G => n1226, D => n1150, Q => 
                           bht_10_15_port);
   bht_reg_12_15_inst : DLH_X1 port map( G => n1232, D => n1150, Q => 
                           bht_12_15_port);
   bht_reg_14_15_inst : DLH_X1 port map( G => n1238, D => n1150, Q => 
                           bht_14_15_port);
   bht_reg_16_15_inst : DLH_X1 port map( G => n1244, D => n1150, Q => 
                           bht_16_15_port);
   bht_reg_18_15_inst : DLH_X1 port map( G => n1250, D => n1150, Q => 
                           bht_18_15_port);
   bht_reg_20_15_inst : DLH_X1 port map( G => n1256, D => n1150, Q => 
                           bht_20_15_port);
   bht_reg_22_15_inst : DLH_X1 port map( G => n1262, D => n1151, Q => 
                           bht_22_15_port);
   bht_reg_24_15_inst : DLH_X1 port map( G => n1268, D => n1151, Q => 
                           bht_24_15_port);
   bht_reg_26_15_inst : DLH_X1 port map( G => n1274, D => n1151, Q => 
                           bht_26_15_port);
   bht_reg_28_15_inst : DLH_X1 port map( G => n1280, D => n1151, Q => 
                           bht_28_15_port);
   bht_reg_30_15_inst : DLH_X1 port map( G => n1286, D => n1151, Q => 
                           bht_30_15_port);
   bht_reg_31_15_inst : DLH_X1 port map( G => n1289, D => n1151, Q => 
                           bht_31_15_port);
   bht_reg_29_15_inst : DLH_X1 port map( G => n1283, D => n1151, Q => 
                           bht_29_15_port);
   bht_reg_27_15_inst : DLH_X1 port map( G => n1277, D => n1151, Q => 
                           bht_27_15_port);
   bht_reg_25_15_inst : DLH_X1 port map( G => n1271, D => n1151, Q => 
                           bht_25_15_port);
   bht_reg_23_15_inst : DLH_X1 port map( G => n1265, D => n1151, Q => 
                           bht_23_15_port);
   bht_reg_21_15_inst : DLH_X1 port map( G => n1259, D => n1151, Q => 
                           bht_21_15_port);
   bht_reg_19_15_inst : DLH_X1 port map( G => n1253, D => n1152, Q => 
                           bht_19_15_port);
   bht_reg_17_15_inst : DLH_X1 port map( G => n1247, D => n1152, Q => 
                           bht_17_15_port);
   bht_reg_15_15_inst : DLH_X1 port map( G => n1241, D => n1152, Q => 
                           bht_15_15_port);
   bht_reg_13_15_inst : DLH_X1 port map( G => n1235, D => n1152, Q => 
                           bht_13_15_port);
   bht_reg_11_15_inst : DLH_X1 port map( G => n1229, D => n1152, Q => 
                           bht_11_15_port);
   bht_reg_9_15_inst : DLH_X1 port map( G => n1223, D => n1152, Q => 
                           bht_9_15_port);
   bht_reg_7_15_inst : DLH_X1 port map( G => n1217, D => n1152, Q => 
                           bht_7_15_port);
   bht_reg_5_15_inst : DLH_X1 port map( G => n1211, D => n1152, Q => 
                           bht_5_15_port);
   bht_reg_3_15_inst : DLH_X1 port map( G => n1205, D => n1152, Q => 
                           bht_3_15_port);
   bht_reg_1_15_inst : DLH_X1 port map( G => n1199, D => n1152, Q => 
                           bht_1_15_port);
   entry_r_reg_14_inst : DLH_X1 port map( G => n961, D => N139, Q => 
                           entry_r_14_port);
   entry_r_delay_reg_14_inst : DFFR_X1 port map( D => entry_r_14_port, CK => 
                           clk, RN => rst, Q => net108079, QN => n22);
   bht_reg_0_14_inst : DLH_X1 port map( G => n1118, D => n1153, Q => 
                           bht_0_14_port);
   bht_reg_2_14_inst : DLH_X1 port map( G => n1202, D => n1153, Q => 
                           bht_2_14_port);
   bht_reg_4_14_inst : DLH_X1 port map( G => n1208, D => n1153, Q => 
                           bht_4_14_port);
   bht_reg_6_14_inst : DLH_X1 port map( G => n1214, D => n1153, Q => 
                           bht_6_14_port);
   bht_reg_8_14_inst : DLH_X1 port map( G => n1220, D => n1153, Q => 
                           bht_8_14_port);
   bht_reg_10_14_inst : DLH_X1 port map( G => n1226, D => n1153, Q => 
                           bht_10_14_port);
   bht_reg_12_14_inst : DLH_X1 port map( G => n1232, D => n1153, Q => 
                           bht_12_14_port);
   bht_reg_14_14_inst : DLH_X1 port map( G => n1238, D => n1153, Q => 
                           bht_14_14_port);
   bht_reg_16_14_inst : DLH_X1 port map( G => n1244, D => n1153, Q => 
                           bht_16_14_port);
   bht_reg_18_14_inst : DLH_X1 port map( G => n1250, D => n1153, Q => 
                           bht_18_14_port);
   bht_reg_20_14_inst : DLH_X1 port map( G => n1256, D => n1153, Q => 
                           bht_20_14_port);
   bht_reg_22_14_inst : DLH_X1 port map( G => n1262, D => n1154, Q => 
                           bht_22_14_port);
   bht_reg_24_14_inst : DLH_X1 port map( G => n1268, D => n1154, Q => 
                           bht_24_14_port);
   bht_reg_26_14_inst : DLH_X1 port map( G => n1274, D => n1154, Q => 
                           bht_26_14_port);
   bht_reg_28_14_inst : DLH_X1 port map( G => n1280, D => n1154, Q => 
                           bht_28_14_port);
   bht_reg_30_14_inst : DLH_X1 port map( G => n1286, D => n1154, Q => 
                           bht_30_14_port);
   bht_reg_31_14_inst : DLH_X1 port map( G => n1289, D => n1154, Q => 
                           bht_31_14_port);
   bht_reg_29_14_inst : DLH_X1 port map( G => n1283, D => n1154, Q => 
                           bht_29_14_port);
   bht_reg_27_14_inst : DLH_X1 port map( G => n1277, D => n1154, Q => 
                           bht_27_14_port);
   bht_reg_25_14_inst : DLH_X1 port map( G => n1271, D => n1154, Q => 
                           bht_25_14_port);
   bht_reg_23_14_inst : DLH_X1 port map( G => n1265, D => n1154, Q => 
                           bht_23_14_port);
   bht_reg_21_14_inst : DLH_X1 port map( G => n1259, D => n1154, Q => 
                           bht_21_14_port);
   bht_reg_19_14_inst : DLH_X1 port map( G => n1253, D => n1155, Q => 
                           bht_19_14_port);
   bht_reg_17_14_inst : DLH_X1 port map( G => n1247, D => n1155, Q => 
                           bht_17_14_port);
   bht_reg_15_14_inst : DLH_X1 port map( G => n1241, D => n1155, Q => 
                           bht_15_14_port);
   bht_reg_13_14_inst : DLH_X1 port map( G => n1235, D => n1155, Q => 
                           bht_13_14_port);
   bht_reg_11_14_inst : DLH_X1 port map( G => n1229, D => n1155, Q => 
                           bht_11_14_port);
   bht_reg_9_14_inst : DLH_X1 port map( G => n1223, D => n1155, Q => 
                           bht_9_14_port);
   bht_reg_7_14_inst : DLH_X1 port map( G => n1217, D => n1155, Q => 
                           bht_7_14_port);
   bht_reg_5_14_inst : DLH_X1 port map( G => n1211, D => n1155, Q => 
                           bht_5_14_port);
   bht_reg_3_14_inst : DLH_X1 port map( G => n1205, D => n1155, Q => 
                           bht_3_14_port);
   bht_reg_1_14_inst : DLH_X1 port map( G => n1199, D => n1155, Q => 
                           bht_1_14_port);
   entry_r_reg_13_inst : DLH_X1 port map( G => n961, D => N138, Q => 
                           entry_r_13_port);
   entry_r_delay_reg_13_inst : DFFR_X1 port map( D => entry_r_13_port, CK => 
                           clk, RN => rst, Q => net108078, QN => n21);
   bht_reg_0_13_inst : DLH_X1 port map( G => n1118, D => n1156, Q => 
                           bht_0_13_port);
   bht_reg_2_13_inst : DLH_X1 port map( G => n1202, D => n1156, Q => 
                           bht_2_13_port);
   bht_reg_4_13_inst : DLH_X1 port map( G => n1208, D => n1156, Q => 
                           bht_4_13_port);
   bht_reg_6_13_inst : DLH_X1 port map( G => n1214, D => n1156, Q => 
                           bht_6_13_port);
   bht_reg_8_13_inst : DLH_X1 port map( G => n1220, D => n1156, Q => 
                           bht_8_13_port);
   bht_reg_10_13_inst : DLH_X1 port map( G => n1226, D => n1156, Q => 
                           bht_10_13_port);
   bht_reg_12_13_inst : DLH_X1 port map( G => n1232, D => n1156, Q => 
                           bht_12_13_port);
   bht_reg_14_13_inst : DLH_X1 port map( G => n1238, D => n1156, Q => 
                           bht_14_13_port);
   bht_reg_16_13_inst : DLH_X1 port map( G => n1244, D => n1156, Q => 
                           bht_16_13_port);
   bht_reg_18_13_inst : DLH_X1 port map( G => n1250, D => n1156, Q => 
                           bht_18_13_port);
   bht_reg_20_13_inst : DLH_X1 port map( G => n1256, D => n1156, Q => 
                           bht_20_13_port);
   bht_reg_22_13_inst : DLH_X1 port map( G => n1262, D => n1157, Q => 
                           bht_22_13_port);
   bht_reg_24_13_inst : DLH_X1 port map( G => n1268, D => n1157, Q => 
                           bht_24_13_port);
   bht_reg_26_13_inst : DLH_X1 port map( G => n1274, D => n1157, Q => 
                           bht_26_13_port);
   bht_reg_28_13_inst : DLH_X1 port map( G => n1280, D => n1157, Q => 
                           bht_28_13_port);
   bht_reg_30_13_inst : DLH_X1 port map( G => n1286, D => n1157, Q => 
                           bht_30_13_port);
   bht_reg_31_13_inst : DLH_X1 port map( G => n1289, D => n1157, Q => 
                           bht_31_13_port);
   bht_reg_29_13_inst : DLH_X1 port map( G => n1283, D => n1157, Q => 
                           bht_29_13_port);
   bht_reg_27_13_inst : DLH_X1 port map( G => n1277, D => n1157, Q => 
                           bht_27_13_port);
   bht_reg_25_13_inst : DLH_X1 port map( G => n1271, D => n1157, Q => 
                           bht_25_13_port);
   bht_reg_23_13_inst : DLH_X1 port map( G => n1265, D => n1157, Q => 
                           bht_23_13_port);
   bht_reg_21_13_inst : DLH_X1 port map( G => n1259, D => n1157, Q => 
                           bht_21_13_port);
   bht_reg_19_13_inst : DLH_X1 port map( G => n1253, D => n1158, Q => 
                           bht_19_13_port);
   bht_reg_17_13_inst : DLH_X1 port map( G => n1247, D => n1158, Q => 
                           bht_17_13_port);
   bht_reg_15_13_inst : DLH_X1 port map( G => n1241, D => n1158, Q => 
                           bht_15_13_port);
   bht_reg_13_13_inst : DLH_X1 port map( G => n1235, D => n1158, Q => 
                           bht_13_13_port);
   bht_reg_11_13_inst : DLH_X1 port map( G => n1229, D => n1158, Q => 
                           bht_11_13_port);
   bht_reg_9_13_inst : DLH_X1 port map( G => n1223, D => n1158, Q => 
                           bht_9_13_port);
   bht_reg_7_13_inst : DLH_X1 port map( G => n1217, D => n1158, Q => 
                           bht_7_13_port);
   bht_reg_5_13_inst : DLH_X1 port map( G => n1211, D => n1158, Q => 
                           bht_5_13_port);
   bht_reg_3_13_inst : DLH_X1 port map( G => n1205, D => n1158, Q => 
                           bht_3_13_port);
   bht_reg_1_13_inst : DLH_X1 port map( G => n1199, D => n1158, Q => 
                           bht_1_13_port);
   entry_r_reg_12_inst : DLH_X1 port map( G => n961, D => N137, Q => 
                           entry_r_12_port);
   entry_r_delay_reg_12_inst : DFFR_X1 port map( D => entry_r_12_port, CK => 
                           clk, RN => rst, Q => net108077, QN => n20);
   bht_reg_0_12_inst : DLH_X1 port map( G => n1118, D => n1159, Q => 
                           bht_0_12_port);
   bht_reg_2_12_inst : DLH_X1 port map( G => n1202, D => n1159, Q => 
                           bht_2_12_port);
   bht_reg_4_12_inst : DLH_X1 port map( G => n1208, D => n1159, Q => 
                           bht_4_12_port);
   bht_reg_6_12_inst : DLH_X1 port map( G => n1214, D => n1159, Q => 
                           bht_6_12_port);
   bht_reg_8_12_inst : DLH_X1 port map( G => n1220, D => n1159, Q => 
                           bht_8_12_port);
   bht_reg_10_12_inst : DLH_X1 port map( G => n1226, D => n1159, Q => 
                           bht_10_12_port);
   bht_reg_12_12_inst : DLH_X1 port map( G => n1232, D => n1159, Q => 
                           bht_12_12_port);
   bht_reg_14_12_inst : DLH_X1 port map( G => n1238, D => n1159, Q => 
                           bht_14_12_port);
   bht_reg_16_12_inst : DLH_X1 port map( G => n1244, D => n1159, Q => 
                           bht_16_12_port);
   bht_reg_18_12_inst : DLH_X1 port map( G => n1250, D => n1159, Q => 
                           bht_18_12_port);
   bht_reg_20_12_inst : DLH_X1 port map( G => n1256, D => n1159, Q => 
                           bht_20_12_port);
   bht_reg_22_12_inst : DLH_X1 port map( G => n1262, D => n1160, Q => 
                           bht_22_12_port);
   bht_reg_24_12_inst : DLH_X1 port map( G => n1268, D => n1160, Q => 
                           bht_24_12_port);
   bht_reg_26_12_inst : DLH_X1 port map( G => n1274, D => n1160, Q => 
                           bht_26_12_port);
   bht_reg_28_12_inst : DLH_X1 port map( G => n1280, D => n1160, Q => 
                           bht_28_12_port);
   bht_reg_30_12_inst : DLH_X1 port map( G => n1286, D => n1160, Q => 
                           bht_30_12_port);
   bht_reg_31_12_inst : DLH_X1 port map( G => n1289, D => n1160, Q => 
                           bht_31_12_port);
   bht_reg_29_12_inst : DLH_X1 port map( G => n1283, D => n1160, Q => 
                           bht_29_12_port);
   bht_reg_27_12_inst : DLH_X1 port map( G => n1277, D => n1160, Q => 
                           bht_27_12_port);
   bht_reg_25_12_inst : DLH_X1 port map( G => n1271, D => n1160, Q => 
                           bht_25_12_port);
   bht_reg_23_12_inst : DLH_X1 port map( G => n1265, D => n1160, Q => 
                           bht_23_12_port);
   bht_reg_21_12_inst : DLH_X1 port map( G => n1259, D => n1160, Q => 
                           bht_21_12_port);
   bht_reg_19_12_inst : DLH_X1 port map( G => n1253, D => n1161, Q => 
                           bht_19_12_port);
   bht_reg_17_12_inst : DLH_X1 port map( G => n1247, D => n1161, Q => 
                           bht_17_12_port);
   bht_reg_15_12_inst : DLH_X1 port map( G => n1241, D => n1161, Q => 
                           bht_15_12_port);
   bht_reg_13_12_inst : DLH_X1 port map( G => n1235, D => n1161, Q => 
                           bht_13_12_port);
   bht_reg_11_12_inst : DLH_X1 port map( G => n1229, D => n1161, Q => 
                           bht_11_12_port);
   bht_reg_9_12_inst : DLH_X1 port map( G => n1223, D => n1161, Q => 
                           bht_9_12_port);
   bht_reg_7_12_inst : DLH_X1 port map( G => n1217, D => n1161, Q => 
                           bht_7_12_port);
   bht_reg_5_12_inst : DLH_X1 port map( G => n1211, D => n1161, Q => 
                           bht_5_12_port);
   bht_reg_3_12_inst : DLH_X1 port map( G => n1205, D => n1161, Q => 
                           bht_3_12_port);
   bht_reg_1_12_inst : DLH_X1 port map( G => n1199, D => n1161, Q => 
                           bht_1_12_port);
   entry_r_reg_11_inst : DLH_X1 port map( G => n961, D => N136, Q => 
                           entry_r_11_port);
   entry_r_delay_reg_11_inst : DFFR_X1 port map( D => entry_r_11_port, CK => 
                           clk, RN => rst, Q => net108076, QN => n19);
   bht_reg_0_11_inst : DLH_X1 port map( G => n1118, D => n1162, Q => 
                           bht_0_11_port);
   bht_reg_2_11_inst : DLH_X1 port map( G => n1202, D => n1162, Q => 
                           bht_2_11_port);
   bht_reg_4_11_inst : DLH_X1 port map( G => n1208, D => n1162, Q => 
                           bht_4_11_port);
   bht_reg_6_11_inst : DLH_X1 port map( G => n1214, D => n1162, Q => 
                           bht_6_11_port);
   bht_reg_8_11_inst : DLH_X1 port map( G => n1220, D => n1162, Q => 
                           bht_8_11_port);
   bht_reg_10_11_inst : DLH_X1 port map( G => n1226, D => n1162, Q => 
                           bht_10_11_port);
   bht_reg_12_11_inst : DLH_X1 port map( G => n1232, D => n1162, Q => 
                           bht_12_11_port);
   bht_reg_14_11_inst : DLH_X1 port map( G => n1238, D => n1162, Q => 
                           bht_14_11_port);
   bht_reg_16_11_inst : DLH_X1 port map( G => n1244, D => n1162, Q => 
                           bht_16_11_port);
   bht_reg_18_11_inst : DLH_X1 port map( G => n1250, D => n1162, Q => 
                           bht_18_11_port);
   bht_reg_20_11_inst : DLH_X1 port map( G => n1256, D => n1162, Q => 
                           bht_20_11_port);
   bht_reg_22_11_inst : DLH_X1 port map( G => n1262, D => n1163, Q => 
                           bht_22_11_port);
   bht_reg_24_11_inst : DLH_X1 port map( G => n1268, D => n1163, Q => 
                           bht_24_11_port);
   bht_reg_26_11_inst : DLH_X1 port map( G => n1274, D => n1163, Q => 
                           bht_26_11_port);
   bht_reg_28_11_inst : DLH_X1 port map( G => n1280, D => n1163, Q => 
                           bht_28_11_port);
   bht_reg_30_11_inst : DLH_X1 port map( G => n1286, D => n1163, Q => 
                           bht_30_11_port);
   bht_reg_31_11_inst : DLH_X1 port map( G => n1289, D => n1163, Q => 
                           bht_31_11_port);
   bht_reg_29_11_inst : DLH_X1 port map( G => n1283, D => n1163, Q => 
                           bht_29_11_port);
   bht_reg_27_11_inst : DLH_X1 port map( G => n1277, D => n1163, Q => 
                           bht_27_11_port);
   bht_reg_25_11_inst : DLH_X1 port map( G => n1271, D => n1163, Q => 
                           bht_25_11_port);
   bht_reg_23_11_inst : DLH_X1 port map( G => n1265, D => n1163, Q => 
                           bht_23_11_port);
   bht_reg_21_11_inst : DLH_X1 port map( G => n1259, D => n1163, Q => 
                           bht_21_11_port);
   bht_reg_19_11_inst : DLH_X1 port map( G => n1253, D => n1164, Q => 
                           bht_19_11_port);
   bht_reg_17_11_inst : DLH_X1 port map( G => n1247, D => n1164, Q => 
                           bht_17_11_port);
   bht_reg_15_11_inst : DLH_X1 port map( G => n1241, D => n1164, Q => 
                           bht_15_11_port);
   bht_reg_13_11_inst : DLH_X1 port map( G => n1235, D => n1164, Q => 
                           bht_13_11_port);
   bht_reg_11_11_inst : DLH_X1 port map( G => n1229, D => n1164, Q => 
                           bht_11_11_port);
   bht_reg_9_11_inst : DLH_X1 port map( G => n1223, D => n1164, Q => 
                           bht_9_11_port);
   bht_reg_7_11_inst : DLH_X1 port map( G => n1217, D => n1164, Q => 
                           bht_7_11_port);
   bht_reg_5_11_inst : DLH_X1 port map( G => n1211, D => n1164, Q => 
                           bht_5_11_port);
   bht_reg_3_11_inst : DLH_X1 port map( G => n1205, D => n1164, Q => 
                           bht_3_11_port);
   bht_reg_1_11_inst : DLH_X1 port map( G => n1199, D => n1164, Q => 
                           bht_1_11_port);
   entry_r_reg_10_inst : DLH_X1 port map( G => n961, D => N135, Q => 
                           entry_r_10_port);
   entry_r_delay_reg_10_inst : DFFR_X1 port map( D => entry_r_10_port, CK => 
                           clk, RN => rst, Q => net108075, QN => n18);
   bht_reg_0_10_inst : DLH_X1 port map( G => n1117, D => n1165, Q => 
                           bht_0_10_port);
   bht_reg_2_10_inst : DLH_X1 port map( G => n1201, D => n1165, Q => 
                           bht_2_10_port);
   bht_reg_4_10_inst : DLH_X1 port map( G => n1207, D => n1165, Q => 
                           bht_4_10_port);
   bht_reg_6_10_inst : DLH_X1 port map( G => n1213, D => n1165, Q => 
                           bht_6_10_port);
   bht_reg_8_10_inst : DLH_X1 port map( G => n1219, D => n1165, Q => 
                           bht_8_10_port);
   bht_reg_10_10_inst : DLH_X1 port map( G => n1225, D => n1165, Q => 
                           bht_10_10_port);
   bht_reg_12_10_inst : DLH_X1 port map( G => n1231, D => n1165, Q => 
                           bht_12_10_port);
   bht_reg_14_10_inst : DLH_X1 port map( G => n1237, D => n1165, Q => 
                           bht_14_10_port);
   bht_reg_16_10_inst : DLH_X1 port map( G => n1243, D => n1165, Q => 
                           bht_16_10_port);
   bht_reg_18_10_inst : DLH_X1 port map( G => n1249, D => n1165, Q => 
                           bht_18_10_port);
   bht_reg_20_10_inst : DLH_X1 port map( G => n1255, D => n1165, Q => 
                           bht_20_10_port);
   bht_reg_22_10_inst : DLH_X1 port map( G => n1261, D => n1166, Q => 
                           bht_22_10_port);
   bht_reg_24_10_inst : DLH_X1 port map( G => n1267, D => n1166, Q => 
                           bht_24_10_port);
   bht_reg_26_10_inst : DLH_X1 port map( G => n1273, D => n1166, Q => 
                           bht_26_10_port);
   bht_reg_28_10_inst : DLH_X1 port map( G => n1279, D => n1166, Q => 
                           bht_28_10_port);
   bht_reg_30_10_inst : DLH_X1 port map( G => n1285, D => n1166, Q => 
                           bht_30_10_port);
   bht_reg_31_10_inst : DLH_X1 port map( G => n1288, D => n1166, Q => 
                           bht_31_10_port);
   bht_reg_29_10_inst : DLH_X1 port map( G => n1282, D => n1166, Q => 
                           bht_29_10_port);
   bht_reg_27_10_inst : DLH_X1 port map( G => n1276, D => n1166, Q => 
                           bht_27_10_port);
   bht_reg_25_10_inst : DLH_X1 port map( G => n1270, D => n1166, Q => 
                           bht_25_10_port);
   bht_reg_23_10_inst : DLH_X1 port map( G => n1264, D => n1166, Q => 
                           bht_23_10_port);
   bht_reg_21_10_inst : DLH_X1 port map( G => n1258, D => n1166, Q => 
                           bht_21_10_port);
   bht_reg_19_10_inst : DLH_X1 port map( G => n1252, D => n1167, Q => 
                           bht_19_10_port);
   bht_reg_17_10_inst : DLH_X1 port map( G => n1246, D => n1167, Q => 
                           bht_17_10_port);
   bht_reg_15_10_inst : DLH_X1 port map( G => n1240, D => n1167, Q => 
                           bht_15_10_port);
   bht_reg_13_10_inst : DLH_X1 port map( G => n1234, D => n1167, Q => 
                           bht_13_10_port);
   bht_reg_11_10_inst : DLH_X1 port map( G => n1228, D => n1167, Q => 
                           bht_11_10_port);
   bht_reg_9_10_inst : DLH_X1 port map( G => n1222, D => n1167, Q => 
                           bht_9_10_port);
   bht_reg_7_10_inst : DLH_X1 port map( G => n1216, D => n1167, Q => 
                           bht_7_10_port);
   bht_reg_5_10_inst : DLH_X1 port map( G => n1210, D => n1167, Q => 
                           bht_5_10_port);
   bht_reg_3_10_inst : DLH_X1 port map( G => n1204, D => n1167, Q => 
                           bht_3_10_port);
   bht_reg_1_10_inst : DLH_X1 port map( G => n1198, D => n1167, Q => 
                           bht_1_10_port);
   entry_r_reg_9_inst : DLH_X1 port map( G => n961, D => N134, Q => 
                           entry_r_9_port);
   entry_r_delay_reg_9_inst : DFFR_X1 port map( D => entry_r_9_port, CK => clk,
                           RN => rst, Q => net108074, QN => n17);
   bht_reg_0_9_inst : DLH_X1 port map( G => n1117, D => n1168, Q => 
                           bht_0_9_port);
   bht_reg_2_9_inst : DLH_X1 port map( G => n1201, D => n1168, Q => 
                           bht_2_9_port);
   bht_reg_4_9_inst : DLH_X1 port map( G => n1207, D => n1168, Q => 
                           bht_4_9_port);
   bht_reg_6_9_inst : DLH_X1 port map( G => n1213, D => n1168, Q => 
                           bht_6_9_port);
   bht_reg_8_9_inst : DLH_X1 port map( G => n1219, D => n1168, Q => 
                           bht_8_9_port);
   bht_reg_10_9_inst : DLH_X1 port map( G => n1225, D => n1168, Q => 
                           bht_10_9_port);
   bht_reg_12_9_inst : DLH_X1 port map( G => n1231, D => n1168, Q => 
                           bht_12_9_port);
   bht_reg_14_9_inst : DLH_X1 port map( G => n1237, D => n1168, Q => 
                           bht_14_9_port);
   bht_reg_16_9_inst : DLH_X1 port map( G => n1243, D => n1168, Q => 
                           bht_16_9_port);
   bht_reg_18_9_inst : DLH_X1 port map( G => n1249, D => n1168, Q => 
                           bht_18_9_port);
   bht_reg_20_9_inst : DLH_X1 port map( G => n1255, D => n1168, Q => 
                           bht_20_9_port);
   bht_reg_22_9_inst : DLH_X1 port map( G => n1261, D => n1169, Q => 
                           bht_22_9_port);
   bht_reg_24_9_inst : DLH_X1 port map( G => n1267, D => n1169, Q => 
                           bht_24_9_port);
   bht_reg_26_9_inst : DLH_X1 port map( G => n1273, D => n1169, Q => 
                           bht_26_9_port);
   bht_reg_28_9_inst : DLH_X1 port map( G => n1279, D => n1169, Q => 
                           bht_28_9_port);
   bht_reg_30_9_inst : DLH_X1 port map( G => n1285, D => n1169, Q => 
                           bht_30_9_port);
   bht_reg_31_9_inst : DLH_X1 port map( G => n1288, D => n1169, Q => 
                           bht_31_9_port);
   bht_reg_29_9_inst : DLH_X1 port map( G => n1282, D => n1169, Q => 
                           bht_29_9_port);
   bht_reg_27_9_inst : DLH_X1 port map( G => n1276, D => n1169, Q => 
                           bht_27_9_port);
   bht_reg_25_9_inst : DLH_X1 port map( G => n1270, D => n1169, Q => 
                           bht_25_9_port);
   bht_reg_23_9_inst : DLH_X1 port map( G => n1264, D => n1169, Q => 
                           bht_23_9_port);
   bht_reg_21_9_inst : DLH_X1 port map( G => n1258, D => n1169, Q => 
                           bht_21_9_port);
   bht_reg_19_9_inst : DLH_X1 port map( G => n1252, D => n1170, Q => 
                           bht_19_9_port);
   bht_reg_17_9_inst : DLH_X1 port map( G => n1246, D => n1170, Q => 
                           bht_17_9_port);
   bht_reg_15_9_inst : DLH_X1 port map( G => n1240, D => n1170, Q => 
                           bht_15_9_port);
   bht_reg_13_9_inst : DLH_X1 port map( G => n1234, D => n1170, Q => 
                           bht_13_9_port);
   bht_reg_11_9_inst : DLH_X1 port map( G => n1228, D => n1170, Q => 
                           bht_11_9_port);
   bht_reg_9_9_inst : DLH_X1 port map( G => n1222, D => n1170, Q => 
                           bht_9_9_port);
   bht_reg_7_9_inst : DLH_X1 port map( G => n1216, D => n1170, Q => 
                           bht_7_9_port);
   bht_reg_5_9_inst : DLH_X1 port map( G => n1210, D => n1170, Q => 
                           bht_5_9_port);
   bht_reg_3_9_inst : DLH_X1 port map( G => n1204, D => n1170, Q => 
                           bht_3_9_port);
   bht_reg_1_9_inst : DLH_X1 port map( G => n1198, D => n1170, Q => 
                           bht_1_9_port);
   entry_r_reg_8_inst : DLH_X1 port map( G => n961, D => N133, Q => 
                           entry_r_8_port);
   entry_r_delay_reg_8_inst : DFFR_X1 port map( D => entry_r_8_port, CK => clk,
                           RN => rst, Q => net108073, QN => n16);
   bht_reg_0_8_inst : DLH_X1 port map( G => n1117, D => n1171, Q => 
                           bht_0_8_port);
   bht_reg_2_8_inst : DLH_X1 port map( G => n1201, D => n1171, Q => 
                           bht_2_8_port);
   bht_reg_4_8_inst : DLH_X1 port map( G => n1207, D => n1171, Q => 
                           bht_4_8_port);
   bht_reg_6_8_inst : DLH_X1 port map( G => n1213, D => n1171, Q => 
                           bht_6_8_port);
   bht_reg_8_8_inst : DLH_X1 port map( G => n1219, D => n1171, Q => 
                           bht_8_8_port);
   bht_reg_10_8_inst : DLH_X1 port map( G => n1225, D => n1171, Q => 
                           bht_10_8_port);
   bht_reg_12_8_inst : DLH_X1 port map( G => n1231, D => n1171, Q => 
                           bht_12_8_port);
   bht_reg_14_8_inst : DLH_X1 port map( G => n1237, D => n1171, Q => 
                           bht_14_8_port);
   bht_reg_16_8_inst : DLH_X1 port map( G => n1243, D => n1171, Q => 
                           bht_16_8_port);
   bht_reg_18_8_inst : DLH_X1 port map( G => n1249, D => n1171, Q => 
                           bht_18_8_port);
   bht_reg_20_8_inst : DLH_X1 port map( G => n1255, D => n1171, Q => 
                           bht_20_8_port);
   bht_reg_22_8_inst : DLH_X1 port map( G => n1261, D => n1172, Q => 
                           bht_22_8_port);
   bht_reg_24_8_inst : DLH_X1 port map( G => n1267, D => n1172, Q => 
                           bht_24_8_port);
   bht_reg_26_8_inst : DLH_X1 port map( G => n1273, D => n1172, Q => 
                           bht_26_8_port);
   bht_reg_28_8_inst : DLH_X1 port map( G => n1279, D => n1172, Q => 
                           bht_28_8_port);
   bht_reg_30_8_inst : DLH_X1 port map( G => n1285, D => n1172, Q => 
                           bht_30_8_port);
   bht_reg_31_8_inst : DLH_X1 port map( G => n1288, D => n1172, Q => 
                           bht_31_8_port);
   bht_reg_29_8_inst : DLH_X1 port map( G => n1282, D => n1172, Q => 
                           bht_29_8_port);
   bht_reg_27_8_inst : DLH_X1 port map( G => n1276, D => n1172, Q => 
                           bht_27_8_port);
   bht_reg_25_8_inst : DLH_X1 port map( G => n1270, D => n1172, Q => 
                           bht_25_8_port);
   bht_reg_23_8_inst : DLH_X1 port map( G => n1264, D => n1172, Q => 
                           bht_23_8_port);
   bht_reg_21_8_inst : DLH_X1 port map( G => n1258, D => n1172, Q => 
                           bht_21_8_port);
   bht_reg_19_8_inst : DLH_X1 port map( G => n1252, D => n1173, Q => 
                           bht_19_8_port);
   bht_reg_17_8_inst : DLH_X1 port map( G => n1246, D => n1173, Q => 
                           bht_17_8_port);
   bht_reg_15_8_inst : DLH_X1 port map( G => n1240, D => n1173, Q => 
                           bht_15_8_port);
   bht_reg_13_8_inst : DLH_X1 port map( G => n1234, D => n1173, Q => 
                           bht_13_8_port);
   bht_reg_11_8_inst : DLH_X1 port map( G => n1228, D => n1173, Q => 
                           bht_11_8_port);
   bht_reg_9_8_inst : DLH_X1 port map( G => n1222, D => n1173, Q => 
                           bht_9_8_port);
   bht_reg_7_8_inst : DLH_X1 port map( G => n1216, D => n1173, Q => 
                           bht_7_8_port);
   bht_reg_5_8_inst : DLH_X1 port map( G => n1210, D => n1173, Q => 
                           bht_5_8_port);
   bht_reg_3_8_inst : DLH_X1 port map( G => n1204, D => n1173, Q => 
                           bht_3_8_port);
   bht_reg_1_8_inst : DLH_X1 port map( G => n1198, D => n1173, Q => 
                           bht_1_8_port);
   entry_r_reg_7_inst : DLH_X1 port map( G => n961, D => N132, Q => 
                           entry_r_7_port);
   entry_r_delay_reg_7_inst : DFFR_X1 port map( D => entry_r_7_port, CK => clk,
                           RN => rst, Q => net108072, QN => n15);
   bht_reg_0_7_inst : DLH_X1 port map( G => n1117, D => n1174, Q => 
                           bht_0_7_port);
   bht_reg_2_7_inst : DLH_X1 port map( G => n1201, D => n1174, Q => 
                           bht_2_7_port);
   bht_reg_4_7_inst : DLH_X1 port map( G => n1207, D => n1174, Q => 
                           bht_4_7_port);
   bht_reg_6_7_inst : DLH_X1 port map( G => n1213, D => n1174, Q => 
                           bht_6_7_port);
   bht_reg_8_7_inst : DLH_X1 port map( G => n1219, D => n1174, Q => 
                           bht_8_7_port);
   bht_reg_10_7_inst : DLH_X1 port map( G => n1225, D => n1174, Q => 
                           bht_10_7_port);
   bht_reg_12_7_inst : DLH_X1 port map( G => n1231, D => n1174, Q => 
                           bht_12_7_port);
   bht_reg_14_7_inst : DLH_X1 port map( G => n1237, D => n1174, Q => 
                           bht_14_7_port);
   bht_reg_16_7_inst : DLH_X1 port map( G => n1243, D => n1174, Q => 
                           bht_16_7_port);
   bht_reg_18_7_inst : DLH_X1 port map( G => n1249, D => n1174, Q => 
                           bht_18_7_port);
   bht_reg_20_7_inst : DLH_X1 port map( G => n1255, D => n1174, Q => 
                           bht_20_7_port);
   bht_reg_22_7_inst : DLH_X1 port map( G => n1261, D => n1175, Q => 
                           bht_22_7_port);
   bht_reg_24_7_inst : DLH_X1 port map( G => n1267, D => n1175, Q => 
                           bht_24_7_port);
   bht_reg_26_7_inst : DLH_X1 port map( G => n1273, D => n1175, Q => 
                           bht_26_7_port);
   bht_reg_28_7_inst : DLH_X1 port map( G => n1279, D => n1175, Q => 
                           bht_28_7_port);
   bht_reg_30_7_inst : DLH_X1 port map( G => n1285, D => n1175, Q => 
                           bht_30_7_port);
   bht_reg_31_7_inst : DLH_X1 port map( G => n1288, D => n1175, Q => 
                           bht_31_7_port);
   bht_reg_29_7_inst : DLH_X1 port map( G => n1282, D => n1175, Q => 
                           bht_29_7_port);
   bht_reg_27_7_inst : DLH_X1 port map( G => n1276, D => n1175, Q => 
                           bht_27_7_port);
   bht_reg_25_7_inst : DLH_X1 port map( G => n1270, D => n1175, Q => 
                           bht_25_7_port);
   bht_reg_23_7_inst : DLH_X1 port map( G => n1264, D => n1175, Q => 
                           bht_23_7_port);
   bht_reg_21_7_inst : DLH_X1 port map( G => n1258, D => n1175, Q => 
                           bht_21_7_port);
   bht_reg_19_7_inst : DLH_X1 port map( G => n1252, D => n1176, Q => 
                           bht_19_7_port);
   bht_reg_17_7_inst : DLH_X1 port map( G => n1246, D => n1176, Q => 
                           bht_17_7_port);
   bht_reg_15_7_inst : DLH_X1 port map( G => n1240, D => n1176, Q => 
                           bht_15_7_port);
   bht_reg_13_7_inst : DLH_X1 port map( G => n1234, D => n1176, Q => 
                           bht_13_7_port);
   bht_reg_11_7_inst : DLH_X1 port map( G => n1228, D => n1176, Q => 
                           bht_11_7_port);
   bht_reg_9_7_inst : DLH_X1 port map( G => n1222, D => n1176, Q => 
                           bht_9_7_port);
   bht_reg_7_7_inst : DLH_X1 port map( G => n1216, D => n1176, Q => 
                           bht_7_7_port);
   bht_reg_5_7_inst : DLH_X1 port map( G => n1210, D => n1176, Q => 
                           bht_5_7_port);
   bht_reg_3_7_inst : DLH_X1 port map( G => n1204, D => n1176, Q => 
                           bht_3_7_port);
   bht_reg_1_7_inst : DLH_X1 port map( G => n1198, D => n1176, Q => 
                           bht_1_7_port);
   entry_r_reg_6_inst : DLH_X1 port map( G => n961, D => N131, Q => 
                           entry_r_6_port);
   entry_r_delay_reg_6_inst : DFFR_X1 port map( D => entry_r_6_port, CK => clk,
                           RN => rst, Q => net108071, QN => n14);
   bht_reg_0_6_inst : DLH_X1 port map( G => n1117, D => n1177, Q => 
                           bht_0_6_port);
   bht_reg_2_6_inst : DLH_X1 port map( G => n1201, D => n1177, Q => 
                           bht_2_6_port);
   bht_reg_4_6_inst : DLH_X1 port map( G => n1207, D => n1177, Q => 
                           bht_4_6_port);
   bht_reg_6_6_inst : DLH_X1 port map( G => n1213, D => n1177, Q => 
                           bht_6_6_port);
   bht_reg_8_6_inst : DLH_X1 port map( G => n1219, D => n1177, Q => 
                           bht_8_6_port);
   bht_reg_10_6_inst : DLH_X1 port map( G => n1225, D => n1177, Q => 
                           bht_10_6_port);
   bht_reg_12_6_inst : DLH_X1 port map( G => n1231, D => n1177, Q => 
                           bht_12_6_port);
   bht_reg_14_6_inst : DLH_X1 port map( G => n1237, D => n1177, Q => 
                           bht_14_6_port);
   bht_reg_16_6_inst : DLH_X1 port map( G => n1243, D => n1177, Q => 
                           bht_16_6_port);
   bht_reg_18_6_inst : DLH_X1 port map( G => n1249, D => n1177, Q => 
                           bht_18_6_port);
   bht_reg_20_6_inst : DLH_X1 port map( G => n1255, D => n1177, Q => 
                           bht_20_6_port);
   bht_reg_22_6_inst : DLH_X1 port map( G => n1261, D => n1178, Q => 
                           bht_22_6_port);
   bht_reg_24_6_inst : DLH_X1 port map( G => n1267, D => n1178, Q => 
                           bht_24_6_port);
   bht_reg_26_6_inst : DLH_X1 port map( G => n1273, D => n1178, Q => 
                           bht_26_6_port);
   bht_reg_28_6_inst : DLH_X1 port map( G => n1279, D => n1178, Q => 
                           bht_28_6_port);
   bht_reg_30_6_inst : DLH_X1 port map( G => n1285, D => n1178, Q => 
                           bht_30_6_port);
   bht_reg_31_6_inst : DLH_X1 port map( G => n1288, D => n1178, Q => 
                           bht_31_6_port);
   bht_reg_29_6_inst : DLH_X1 port map( G => n1282, D => n1178, Q => 
                           bht_29_6_port);
   bht_reg_27_6_inst : DLH_X1 port map( G => n1276, D => n1178, Q => 
                           bht_27_6_port);
   bht_reg_25_6_inst : DLH_X1 port map( G => n1270, D => n1178, Q => 
                           bht_25_6_port);
   bht_reg_23_6_inst : DLH_X1 port map( G => n1264, D => n1178, Q => 
                           bht_23_6_port);
   bht_reg_21_6_inst : DLH_X1 port map( G => n1258, D => n1178, Q => 
                           bht_21_6_port);
   bht_reg_19_6_inst : DLH_X1 port map( G => n1252, D => n1179, Q => 
                           bht_19_6_port);
   bht_reg_17_6_inst : DLH_X1 port map( G => n1246, D => n1179, Q => 
                           bht_17_6_port);
   bht_reg_15_6_inst : DLH_X1 port map( G => n1240, D => n1179, Q => 
                           bht_15_6_port);
   bht_reg_13_6_inst : DLH_X1 port map( G => n1234, D => n1179, Q => 
                           bht_13_6_port);
   bht_reg_11_6_inst : DLH_X1 port map( G => n1228, D => n1179, Q => 
                           bht_11_6_port);
   bht_reg_9_6_inst : DLH_X1 port map( G => n1222, D => n1179, Q => 
                           bht_9_6_port);
   bht_reg_7_6_inst : DLH_X1 port map( G => n1216, D => n1179, Q => 
                           bht_7_6_port);
   bht_reg_5_6_inst : DLH_X1 port map( G => n1210, D => n1179, Q => 
                           bht_5_6_port);
   bht_reg_3_6_inst : DLH_X1 port map( G => n1204, D => n1179, Q => 
                           bht_3_6_port);
   bht_reg_1_6_inst : DLH_X1 port map( G => n1198, D => n1179, Q => 
                           bht_1_6_port);
   entry_r_reg_5_inst : DLH_X1 port map( G => n961, D => N130, Q => 
                           entry_r_5_port);
   entry_r_delay_reg_5_inst : DFFR_X1 port map( D => entry_r_5_port, CK => clk,
                           RN => rst, Q => net108070, QN => n13);
   bht_reg_0_5_inst : DLH_X1 port map( G => n1117, D => n1180, Q => 
                           bht_0_5_port);
   bht_reg_2_5_inst : DLH_X1 port map( G => n1201, D => n1180, Q => 
                           bht_2_5_port);
   bht_reg_4_5_inst : DLH_X1 port map( G => n1207, D => n1180, Q => 
                           bht_4_5_port);
   bht_reg_6_5_inst : DLH_X1 port map( G => n1213, D => n1180, Q => 
                           bht_6_5_port);
   bht_reg_8_5_inst : DLH_X1 port map( G => n1219, D => n1180, Q => 
                           bht_8_5_port);
   bht_reg_10_5_inst : DLH_X1 port map( G => n1225, D => n1180, Q => 
                           bht_10_5_port);
   bht_reg_12_5_inst : DLH_X1 port map( G => n1231, D => n1180, Q => 
                           bht_12_5_port);
   bht_reg_14_5_inst : DLH_X1 port map( G => n1237, D => n1180, Q => 
                           bht_14_5_port);
   bht_reg_16_5_inst : DLH_X1 port map( G => n1243, D => n1180, Q => 
                           bht_16_5_port);
   bht_reg_18_5_inst : DLH_X1 port map( G => n1249, D => n1180, Q => 
                           bht_18_5_port);
   bht_reg_20_5_inst : DLH_X1 port map( G => n1255, D => n1180, Q => 
                           bht_20_5_port);
   bht_reg_22_5_inst : DLH_X1 port map( G => n1261, D => n1181, Q => 
                           bht_22_5_port);
   bht_reg_24_5_inst : DLH_X1 port map( G => n1267, D => n1181, Q => 
                           bht_24_5_port);
   bht_reg_26_5_inst : DLH_X1 port map( G => n1273, D => n1181, Q => 
                           bht_26_5_port);
   bht_reg_28_5_inst : DLH_X1 port map( G => n1279, D => n1181, Q => 
                           bht_28_5_port);
   bht_reg_30_5_inst : DLH_X1 port map( G => n1285, D => n1181, Q => 
                           bht_30_5_port);
   bht_reg_31_5_inst : DLH_X1 port map( G => n1288, D => n1181, Q => 
                           bht_31_5_port);
   bht_reg_29_5_inst : DLH_X1 port map( G => n1282, D => n1181, Q => 
                           bht_29_5_port);
   bht_reg_27_5_inst : DLH_X1 port map( G => n1276, D => n1181, Q => 
                           bht_27_5_port);
   bht_reg_25_5_inst : DLH_X1 port map( G => n1270, D => n1181, Q => 
                           bht_25_5_port);
   bht_reg_23_5_inst : DLH_X1 port map( G => n1264, D => n1181, Q => 
                           bht_23_5_port);
   bht_reg_21_5_inst : DLH_X1 port map( G => n1258, D => n1181, Q => 
                           bht_21_5_port);
   bht_reg_19_5_inst : DLH_X1 port map( G => n1252, D => n1182, Q => 
                           bht_19_5_port);
   bht_reg_17_5_inst : DLH_X1 port map( G => n1246, D => n1182, Q => 
                           bht_17_5_port);
   bht_reg_15_5_inst : DLH_X1 port map( G => n1240, D => n1182, Q => 
                           bht_15_5_port);
   bht_reg_13_5_inst : DLH_X1 port map( G => n1234, D => n1182, Q => 
                           bht_13_5_port);
   bht_reg_11_5_inst : DLH_X1 port map( G => n1228, D => n1182, Q => 
                           bht_11_5_port);
   bht_reg_9_5_inst : DLH_X1 port map( G => n1222, D => n1182, Q => 
                           bht_9_5_port);
   bht_reg_7_5_inst : DLH_X1 port map( G => n1216, D => n1182, Q => 
                           bht_7_5_port);
   bht_reg_5_5_inst : DLH_X1 port map( G => n1210, D => n1182, Q => 
                           bht_5_5_port);
   bht_reg_3_5_inst : DLH_X1 port map( G => n1204, D => n1182, Q => 
                           bht_3_5_port);
   bht_reg_1_5_inst : DLH_X1 port map( G => n1198, D => n1182, Q => 
                           bht_1_5_port);
   entry_r_reg_4_inst : DLH_X1 port map( G => n961, D => N129, Q => 
                           entry_r_4_port);
   entry_r_delay_reg_4_inst : DFFR_X1 port map( D => entry_r_4_port, CK => clk,
                           RN => rst, Q => net108069, QN => n12);
   bht_reg_0_4_inst : DLH_X1 port map( G => n1117, D => n1183, Q => 
                           bht_0_4_port);
   bht_reg_2_4_inst : DLH_X1 port map( G => n1201, D => n1183, Q => 
                           bht_2_4_port);
   bht_reg_4_4_inst : DLH_X1 port map( G => n1207, D => n1183, Q => 
                           bht_4_4_port);
   bht_reg_6_4_inst : DLH_X1 port map( G => n1213, D => n1183, Q => 
                           bht_6_4_port);
   bht_reg_8_4_inst : DLH_X1 port map( G => n1219, D => n1183, Q => 
                           bht_8_4_port);
   bht_reg_10_4_inst : DLH_X1 port map( G => n1225, D => n1183, Q => 
                           bht_10_4_port);
   bht_reg_12_4_inst : DLH_X1 port map( G => n1231, D => n1183, Q => 
                           bht_12_4_port);
   bht_reg_14_4_inst : DLH_X1 port map( G => n1237, D => n1183, Q => 
                           bht_14_4_port);
   bht_reg_16_4_inst : DLH_X1 port map( G => n1243, D => n1183, Q => 
                           bht_16_4_port);
   bht_reg_18_4_inst : DLH_X1 port map( G => n1249, D => n1183, Q => 
                           bht_18_4_port);
   bht_reg_20_4_inst : DLH_X1 port map( G => n1255, D => n1183, Q => 
                           bht_20_4_port);
   bht_reg_22_4_inst : DLH_X1 port map( G => n1261, D => n1184, Q => 
                           bht_22_4_port);
   bht_reg_24_4_inst : DLH_X1 port map( G => n1267, D => n1184, Q => 
                           bht_24_4_port);
   bht_reg_26_4_inst : DLH_X1 port map( G => n1273, D => n1184, Q => 
                           bht_26_4_port);
   bht_reg_28_4_inst : DLH_X1 port map( G => n1279, D => n1184, Q => 
                           bht_28_4_port);
   bht_reg_30_4_inst : DLH_X1 port map( G => n1285, D => n1184, Q => 
                           bht_30_4_port);
   bht_reg_31_4_inst : DLH_X1 port map( G => n1288, D => n1184, Q => 
                           bht_31_4_port);
   bht_reg_29_4_inst : DLH_X1 port map( G => n1282, D => n1184, Q => 
                           bht_29_4_port);
   bht_reg_27_4_inst : DLH_X1 port map( G => n1276, D => n1184, Q => 
                           bht_27_4_port);
   bht_reg_25_4_inst : DLH_X1 port map( G => n1270, D => n1184, Q => 
                           bht_25_4_port);
   bht_reg_23_4_inst : DLH_X1 port map( G => n1264, D => n1184, Q => 
                           bht_23_4_port);
   bht_reg_21_4_inst : DLH_X1 port map( G => n1258, D => n1184, Q => 
                           bht_21_4_port);
   bht_reg_19_4_inst : DLH_X1 port map( G => n1252, D => n1185, Q => 
                           bht_19_4_port);
   bht_reg_17_4_inst : DLH_X1 port map( G => n1246, D => n1185, Q => 
                           bht_17_4_port);
   bht_reg_15_4_inst : DLH_X1 port map( G => n1240, D => n1185, Q => 
                           bht_15_4_port);
   bht_reg_13_4_inst : DLH_X1 port map( G => n1234, D => n1185, Q => 
                           bht_13_4_port);
   bht_reg_11_4_inst : DLH_X1 port map( G => n1228, D => n1185, Q => 
                           bht_11_4_port);
   bht_reg_9_4_inst : DLH_X1 port map( G => n1222, D => n1185, Q => 
                           bht_9_4_port);
   bht_reg_7_4_inst : DLH_X1 port map( G => n1216, D => n1185, Q => 
                           bht_7_4_port);
   bht_reg_5_4_inst : DLH_X1 port map( G => n1210, D => n1185, Q => 
                           bht_5_4_port);
   bht_reg_3_4_inst : DLH_X1 port map( G => n1204, D => n1185, Q => 
                           bht_3_4_port);
   bht_reg_1_4_inst : DLH_X1 port map( G => n1198, D => n1185, Q => 
                           bht_1_4_port);
   entry_r_reg_3_inst : DLH_X1 port map( G => n961, D => N128, Q => 
                           entry_r_3_port);
   entry_r_delay_reg_3_inst : DFFR_X1 port map( D => entry_r_3_port, CK => clk,
                           RN => rst, Q => net108068, QN => n11);
   bht_reg_0_3_inst : DLH_X1 port map( G => n1117, D => n1186, Q => 
                           bht_0_3_port);
   bht_reg_2_3_inst : DLH_X1 port map( G => n1201, D => n1186, Q => 
                           bht_2_3_port);
   bht_reg_4_3_inst : DLH_X1 port map( G => n1207, D => n1186, Q => 
                           bht_4_3_port);
   bht_reg_6_3_inst : DLH_X1 port map( G => n1213, D => n1186, Q => 
                           bht_6_3_port);
   bht_reg_8_3_inst : DLH_X1 port map( G => n1219, D => n1186, Q => 
                           bht_8_3_port);
   bht_reg_10_3_inst : DLH_X1 port map( G => n1225, D => n1186, Q => 
                           bht_10_3_port);
   bht_reg_12_3_inst : DLH_X1 port map( G => n1231, D => n1186, Q => 
                           bht_12_3_port);
   bht_reg_14_3_inst : DLH_X1 port map( G => n1237, D => n1186, Q => 
                           bht_14_3_port);
   bht_reg_16_3_inst : DLH_X1 port map( G => n1243, D => n1186, Q => 
                           bht_16_3_port);
   bht_reg_18_3_inst : DLH_X1 port map( G => n1249, D => n1186, Q => 
                           bht_18_3_port);
   bht_reg_20_3_inst : DLH_X1 port map( G => n1255, D => n1186, Q => 
                           bht_20_3_port);
   bht_reg_22_3_inst : DLH_X1 port map( G => n1261, D => n1187, Q => 
                           bht_22_3_port);
   bht_reg_24_3_inst : DLH_X1 port map( G => n1267, D => n1187, Q => 
                           bht_24_3_port);
   bht_reg_26_3_inst : DLH_X1 port map( G => n1273, D => n1187, Q => 
                           bht_26_3_port);
   bht_reg_28_3_inst : DLH_X1 port map( G => n1279, D => n1187, Q => 
                           bht_28_3_port);
   bht_reg_30_3_inst : DLH_X1 port map( G => n1285, D => n1187, Q => 
                           bht_30_3_port);
   bht_reg_31_3_inst : DLH_X1 port map( G => n1288, D => n1187, Q => 
                           bht_31_3_port);
   bht_reg_29_3_inst : DLH_X1 port map( G => n1282, D => n1187, Q => 
                           bht_29_3_port);
   bht_reg_27_3_inst : DLH_X1 port map( G => n1276, D => n1187, Q => 
                           bht_27_3_port);
   bht_reg_25_3_inst : DLH_X1 port map( G => n1270, D => n1187, Q => 
                           bht_25_3_port);
   bht_reg_23_3_inst : DLH_X1 port map( G => n1264, D => n1187, Q => 
                           bht_23_3_port);
   bht_reg_21_3_inst : DLH_X1 port map( G => n1258, D => n1187, Q => 
                           bht_21_3_port);
   bht_reg_19_3_inst : DLH_X1 port map( G => n1252, D => n1188, Q => 
                           bht_19_3_port);
   bht_reg_17_3_inst : DLH_X1 port map( G => n1246, D => n1188, Q => 
                           bht_17_3_port);
   bht_reg_15_3_inst : DLH_X1 port map( G => n1240, D => n1188, Q => 
                           bht_15_3_port);
   bht_reg_13_3_inst : DLH_X1 port map( G => n1234, D => n1188, Q => 
                           bht_13_3_port);
   bht_reg_11_3_inst : DLH_X1 port map( G => n1228, D => n1188, Q => 
                           bht_11_3_port);
   bht_reg_9_3_inst : DLH_X1 port map( G => n1222, D => n1188, Q => 
                           bht_9_3_port);
   bht_reg_7_3_inst : DLH_X1 port map( G => n1216, D => n1188, Q => 
                           bht_7_3_port);
   bht_reg_5_3_inst : DLH_X1 port map( G => n1210, D => n1188, Q => 
                           bht_5_3_port);
   bht_reg_3_3_inst : DLH_X1 port map( G => n1204, D => n1188, Q => 
                           bht_3_3_port);
   bht_reg_1_3_inst : DLH_X1 port map( G => n1198, D => n1188, Q => 
                           bht_1_3_port);
   entry_r_reg_2_inst : DLH_X1 port map( G => n961, D => N127, Q => 
                           entry_r_2_port);
   entry_r_delay_reg_2_inst : DFFR_X1 port map( D => entry_r_2_port, CK => clk,
                           RN => rst, Q => net108067, QN => n10);
   bht_reg_0_2_inst : DLH_X1 port map( G => n1117, D => n1189, Q => 
                           bht_0_2_port);
   bht_reg_2_2_inst : DLH_X1 port map( G => n1201, D => n1189, Q => 
                           bht_2_2_port);
   bht_reg_4_2_inst : DLH_X1 port map( G => n1207, D => n1189, Q => 
                           bht_4_2_port);
   bht_reg_6_2_inst : DLH_X1 port map( G => n1213, D => n1189, Q => 
                           bht_6_2_port);
   bht_reg_8_2_inst : DLH_X1 port map( G => n1219, D => n1189, Q => 
                           bht_8_2_port);
   bht_reg_10_2_inst : DLH_X1 port map( G => n1225, D => n1189, Q => 
                           bht_10_2_port);
   bht_reg_12_2_inst : DLH_X1 port map( G => n1231, D => n1189, Q => 
                           bht_12_2_port);
   bht_reg_14_2_inst : DLH_X1 port map( G => n1237, D => n1189, Q => 
                           bht_14_2_port);
   bht_reg_16_2_inst : DLH_X1 port map( G => n1243, D => n1189, Q => 
                           bht_16_2_port);
   bht_reg_18_2_inst : DLH_X1 port map( G => n1249, D => n1189, Q => 
                           bht_18_2_port);
   bht_reg_20_2_inst : DLH_X1 port map( G => n1255, D => n1189, Q => 
                           bht_20_2_port);
   bht_reg_22_2_inst : DLH_X1 port map( G => n1261, D => n1190, Q => 
                           bht_22_2_port);
   bht_reg_24_2_inst : DLH_X1 port map( G => n1267, D => n1190, Q => 
                           bht_24_2_port);
   bht_reg_26_2_inst : DLH_X1 port map( G => n1273, D => n1190, Q => 
                           bht_26_2_port);
   bht_reg_28_2_inst : DLH_X1 port map( G => n1279, D => n1190, Q => 
                           bht_28_2_port);
   bht_reg_30_2_inst : DLH_X1 port map( G => n1285, D => n1190, Q => 
                           bht_30_2_port);
   bht_reg_31_2_inst : DLH_X1 port map( G => n1288, D => n1190, Q => 
                           bht_31_2_port);
   bht_reg_29_2_inst : DLH_X1 port map( G => n1282, D => n1190, Q => 
                           bht_29_2_port);
   bht_reg_27_2_inst : DLH_X1 port map( G => n1276, D => n1190, Q => 
                           bht_27_2_port);
   bht_reg_25_2_inst : DLH_X1 port map( G => n1270, D => n1190, Q => 
                           bht_25_2_port);
   bht_reg_23_2_inst : DLH_X1 port map( G => n1264, D => n1190, Q => 
                           bht_23_2_port);
   bht_reg_21_2_inst : DLH_X1 port map( G => n1258, D => n1190, Q => 
                           bht_21_2_port);
   bht_reg_19_2_inst : DLH_X1 port map( G => n1252, D => n1191, Q => 
                           bht_19_2_port);
   bht_reg_17_2_inst : DLH_X1 port map( G => n1246, D => n1191, Q => 
                           bht_17_2_port);
   bht_reg_15_2_inst : DLH_X1 port map( G => n1240, D => n1191, Q => 
                           bht_15_2_port);
   bht_reg_13_2_inst : DLH_X1 port map( G => n1234, D => n1191, Q => 
                           bht_13_2_port);
   bht_reg_11_2_inst : DLH_X1 port map( G => n1228, D => n1191, Q => 
                           bht_11_2_port);
   bht_reg_9_2_inst : DLH_X1 port map( G => n1222, D => n1191, Q => 
                           bht_9_2_port);
   bht_reg_7_2_inst : DLH_X1 port map( G => n1216, D => n1191, Q => 
                           bht_7_2_port);
   bht_reg_5_2_inst : DLH_X1 port map( G => n1210, D => n1191, Q => 
                           bht_5_2_port);
   bht_reg_3_2_inst : DLH_X1 port map( G => n1204, D => n1191, Q => 
                           bht_3_2_port);
   bht_reg_1_2_inst : DLH_X1 port map( G => n1198, D => n1191, Q => 
                           bht_1_2_port);
   sig_brt_delay_reg : DFFR_X1 port map( D => n797, CK => clk, RN => rst, Q => 
                           sig_brt_delay, QN => n799);
   bht_reg_0_0_inst : DLH_X1 port map( G => n1117, D => n1197, Q => 
                           bht_0_0_port);
   bht_reg_2_0_inst : DLH_X1 port map( G => n1201, D => n1197, Q => 
                           bht_2_0_port);
   bht_reg_4_0_inst : DLH_X1 port map( G => n1207, D => n1197, Q => 
                           bht_4_0_port);
   bht_reg_6_0_inst : DLH_X1 port map( G => n1213, D => n1197, Q => 
                           bht_6_0_port);
   bht_reg_8_0_inst : DLH_X1 port map( G => n1219, D => n1197, Q => 
                           bht_8_0_port);
   bht_reg_10_0_inst : DLH_X1 port map( G => n1225, D => n1197, Q => 
                           bht_10_0_port);
   bht_reg_12_0_inst : DLH_X1 port map( G => n1231, D => n1197, Q => 
                           bht_12_0_port);
   bht_reg_14_0_inst : DLH_X1 port map( G => n1237, D => n1197, Q => 
                           bht_14_0_port);
   bht_reg_16_0_inst : DLH_X1 port map( G => n1243, D => n1197, Q => 
                           bht_16_0_port);
   bht_reg_18_0_inst : DLH_X1 port map( G => n1249, D => n1197, Q => 
                           bht_18_0_port);
   bht_reg_20_0_inst : DLH_X1 port map( G => n1255, D => n1196, Q => 
                           bht_20_0_port);
   bht_reg_22_0_inst : DLH_X1 port map( G => n1261, D => n1196, Q => 
                           bht_22_0_port);
   bht_reg_24_0_inst : DLH_X1 port map( G => n1267, D => n1196, Q => 
                           bht_24_0_port);
   bht_reg_26_0_inst : DLH_X1 port map( G => n1273, D => n1196, Q => 
                           bht_26_0_port);
   bht_reg_28_0_inst : DLH_X1 port map( G => n1279, D => n1196, Q => 
                           bht_28_0_port);
   bht_reg_30_0_inst : DLH_X1 port map( G => n1285, D => n1196, Q => 
                           bht_30_0_port);
   bht_reg_31_0_inst : DLH_X1 port map( G => n1288, D => n1196, Q => 
                           bht_31_0_port);
   bht_reg_29_0_inst : DLH_X1 port map( G => n1282, D => n1196, Q => 
                           bht_29_0_port);
   bht_reg_27_0_inst : DLH_X1 port map( G => n1276, D => n1196, Q => 
                           bht_27_0_port);
   bht_reg_25_0_inst : DLH_X1 port map( G => n1270, D => n1196, Q => 
                           bht_25_0_port);
   bht_reg_23_0_inst : DLH_X1 port map( G => n1264, D => n1196, Q => 
                           bht_23_0_port);
   bht_reg_21_0_inst : DLH_X1 port map( G => n1258, D => n1195, Q => 
                           bht_21_0_port);
   bht_reg_19_0_inst : DLH_X1 port map( G => n1252, D => n1195, Q => 
                           bht_19_0_port);
   bht_reg_17_0_inst : DLH_X1 port map( G => n1246, D => n1195, Q => 
                           bht_17_0_port);
   bht_reg_15_0_inst : DLH_X1 port map( G => n1240, D => n1195, Q => 
                           bht_15_0_port);
   bht_reg_13_0_inst : DLH_X1 port map( G => n1234, D => n1195, Q => 
                           bht_13_0_port);
   bht_reg_11_0_inst : DLH_X1 port map( G => n1228, D => n1195, Q => 
                           bht_11_0_port);
   bht_reg_9_0_inst : DLH_X1 port map( G => n1222, D => n1195, Q => 
                           bht_9_0_port);
   bht_reg_7_0_inst : DLH_X1 port map( G => n1216, D => n1195, Q => 
                           bht_7_0_port);
   bht_reg_5_0_inst : DLH_X1 port map( G => n1210, D => n1195, Q => 
                           bht_5_0_port);
   bht_reg_3_0_inst : DLH_X1 port map( G => n1204, D => n1195, Q => 
                           bht_3_0_port);
   bht_reg_1_0_inst : DLH_X1 port map( G => n1198, D => n1195, Q => 
                           bht_1_0_port);
   entry_r_reg_0_inst : DLH_X1 port map( G => n1292, D => N125, Q => 
                           entry_r_0_port);
   entry_r_delay_reg_0_inst : DFFR_X1 port map( D => entry_r_0_port, CK => clk,
                           RN => rst, Q => net108066, QN => n860);
   bht_reg_0_1_inst : DLH_X1 port map( G => n1117, D => n1194, Q => 
                           bht_0_1_port);
   bht_reg_2_1_inst : DLH_X1 port map( G => n1201, D => n1194, Q => 
                           bht_2_1_port);
   bht_reg_4_1_inst : DLH_X1 port map( G => n1207, D => n1194, Q => 
                           bht_4_1_port);
   bht_reg_6_1_inst : DLH_X1 port map( G => n1213, D => n1194, Q => 
                           bht_6_1_port);
   bht_reg_8_1_inst : DLH_X1 port map( G => n1219, D => n1194, Q => 
                           bht_8_1_port);
   bht_reg_10_1_inst : DLH_X1 port map( G => n1225, D => n1194, Q => 
                           bht_10_1_port);
   bht_reg_12_1_inst : DLH_X1 port map( G => n1231, D => n1194, Q => 
                           bht_12_1_port);
   bht_reg_14_1_inst : DLH_X1 port map( G => n1237, D => n1194, Q => 
                           bht_14_1_port);
   bht_reg_16_1_inst : DLH_X1 port map( G => n1243, D => n1194, Q => 
                           bht_16_1_port);
   bht_reg_18_1_inst : DLH_X1 port map( G => n1249, D => n1194, Q => 
                           bht_18_1_port);
   bht_reg_20_1_inst : DLH_X1 port map( G => n1255, D => n1193, Q => 
                           bht_20_1_port);
   bht_reg_22_1_inst : DLH_X1 port map( G => n1261, D => n1193, Q => 
                           bht_22_1_port);
   bht_reg_24_1_inst : DLH_X1 port map( G => n1267, D => n1193, Q => 
                           bht_24_1_port);
   bht_reg_26_1_inst : DLH_X1 port map( G => n1273, D => n1193, Q => 
                           bht_26_1_port);
   bht_reg_28_1_inst : DLH_X1 port map( G => n1279, D => n1193, Q => 
                           bht_28_1_port);
   bht_reg_30_1_inst : DLH_X1 port map( G => n1285, D => n1193, Q => 
                           bht_30_1_port);
   bht_reg_31_1_inst : DLH_X1 port map( G => n1288, D => n1193, Q => 
                           bht_31_1_port);
   bht_reg_29_1_inst : DLH_X1 port map( G => n1282, D => n1193, Q => 
                           bht_29_1_port);
   bht_reg_27_1_inst : DLH_X1 port map( G => n1276, D => n1193, Q => 
                           bht_27_1_port);
   bht_reg_25_1_inst : DLH_X1 port map( G => n1270, D => n1193, Q => 
                           bht_25_1_port);
   bht_reg_23_1_inst : DLH_X1 port map( G => n1264, D => n1193, Q => 
                           bht_23_1_port);
   bht_reg_21_1_inst : DLH_X1 port map( G => n1258, D => n1192, Q => 
                           bht_21_1_port);
   bht_reg_19_1_inst : DLH_X1 port map( G => n1252, D => n1192, Q => 
                           bht_19_1_port);
   bht_reg_17_1_inst : DLH_X1 port map( G => n1246, D => n1192, Q => 
                           bht_17_1_port);
   bht_reg_15_1_inst : DLH_X1 port map( G => n1240, D => n1192, Q => 
                           bht_15_1_port);
   bht_reg_13_1_inst : DLH_X1 port map( G => n1234, D => n1192, Q => 
                           bht_13_1_port);
   bht_reg_11_1_inst : DLH_X1 port map( G => n1228, D => n1192, Q => 
                           bht_11_1_port);
   bht_reg_9_1_inst : DLH_X1 port map( G => n1222, D => n1192, Q => 
                           bht_9_1_port);
   bht_reg_7_1_inst : DLH_X1 port map( G => n1216, D => n1192, Q => 
                           bht_7_1_port);
   bht_reg_5_1_inst : DLH_X1 port map( G => n1210, D => n1192, Q => 
                           bht_5_1_port);
   bht_reg_3_1_inst : DLH_X1 port map( G => n1204, D => n1192, Q => 
                           bht_3_1_port);
   bht_reg_1_1_inst : DLH_X1 port map( G => n1198, D => n1192, Q => 
                           bht_1_1_port);
   entry_r_reg_1_inst : DLH_X1 port map( G => n1292, D => N126, Q => 
                           entry_r_1_port);
   entry_r_delay_reg_1_inst : DFFR_X1 port map( D => entry_r_1_port, CK => clk,
                           RN => rst, Q => n854, QN => net108065);
   entry_r_reg_25_inst : DLH_X1 port map( G => n962, D => N150, Q => 
                           entry_r_25_port);
   entry_r_delay_reg_25_inst : DFFR_X1 port map( D => entry_r_25_port, CK => 
                           clk, RN => rst, Q => net108064, QN => n9);
   bht_reg_0_25_inst : DLH_X1 port map( G => n1119, D => n1120, Q => 
                           bht_0_25_port);
   bht_reg_2_25_inst : DLH_X1 port map( G => n1203, D => n1120, Q => 
                           bht_2_25_port);
   bht_reg_4_25_inst : DLH_X1 port map( G => n1209, D => n1120, Q => 
                           bht_4_25_port);
   bht_reg_6_25_inst : DLH_X1 port map( G => n1215, D => n1120, Q => 
                           bht_6_25_port);
   bht_reg_8_25_inst : DLH_X1 port map( G => n1221, D => n1120, Q => 
                           bht_8_25_port);
   bht_reg_10_25_inst : DLH_X1 port map( G => n1227, D => n1120, Q => 
                           bht_10_25_port);
   bht_reg_12_25_inst : DLH_X1 port map( G => n1233, D => n1120, Q => 
                           bht_12_25_port);
   bht_reg_14_25_inst : DLH_X1 port map( G => n1239, D => n1120, Q => 
                           bht_14_25_port);
   bht_reg_16_25_inst : DLH_X1 port map( G => n1245, D => n1120, Q => 
                           bht_16_25_port);
   bht_reg_18_25_inst : DLH_X1 port map( G => n1251, D => n1120, Q => 
                           bht_18_25_port);
   bht_reg_20_25_inst : DLH_X1 port map( G => n1257, D => n1121, Q => 
                           bht_20_25_port);
   bht_reg_22_25_inst : DLH_X1 port map( G => n1263, D => n1121, Q => 
                           bht_22_25_port);
   bht_reg_24_25_inst : DLH_X1 port map( G => n1269, D => n1121, Q => 
                           bht_24_25_port);
   bht_reg_26_25_inst : DLH_X1 port map( G => n1275, D => n1121, Q => 
                           bht_26_25_port);
   bht_reg_28_25_inst : DLH_X1 port map( G => n1281, D => n1121, Q => 
                           bht_28_25_port);
   bht_reg_30_25_inst : DLH_X1 port map( G => n1287, D => n1121, Q => 
                           bht_30_25_port);
   bht_reg_29_25_inst : DLH_X1 port map( G => n1284, D => n1121, Q => 
                           bht_29_25_port);
   bht_reg_27_25_inst : DLH_X1 port map( G => n1278, D => n1121, Q => 
                           bht_27_25_port);
   bht_reg_25_25_inst : DLH_X1 port map( G => n1272, D => n1121, Q => 
                           bht_25_25_port);
   bht_reg_23_25_inst : DLH_X1 port map( G => n1266, D => n1121, Q => 
                           bht_23_25_port);
   bht_reg_21_25_inst : DLH_X1 port map( G => n1260, D => n1121, Q => 
                           bht_21_25_port);
   bht_reg_19_25_inst : DLH_X1 port map( G => n1254, D => n1122, Q => 
                           bht_19_25_port);
   bht_reg_17_25_inst : DLH_X1 port map( G => n1248, D => n1122, Q => 
                           bht_17_25_port);
   bht_reg_15_25_inst : DLH_X1 port map( G => n1242, D => n1122, Q => 
                           bht_15_25_port);
   bht_reg_13_25_inst : DLH_X1 port map( G => n1236, D => n1122, Q => 
                           bht_13_25_port);
   bht_reg_11_25_inst : DLH_X1 port map( G => n1230, D => n1122, Q => 
                           bht_11_25_port);
   bht_reg_9_25_inst : DLH_X1 port map( G => n1224, D => n1122, Q => 
                           bht_9_25_port);
   bht_reg_7_25_inst : DLH_X1 port map( G => n1218, D => n1122, Q => 
                           bht_7_25_port);
   bht_reg_5_25_inst : DLH_X1 port map( G => n1212, D => n1122, Q => 
                           bht_5_25_port);
   bht_reg_3_25_inst : DLH_X1 port map( G => n1206, D => n1122, Q => 
                           bht_3_25_port);
   bht_reg_1_25_inst : DLH_X1 port map( G => n1200, D => n1122, Q => 
                           bht_1_25_port);
   U823 : AND2_X2 port map( A1 => n851, A2 => addr(4), ZN => n828);
   U837 : XOR2_X1 port map( A => n107, B => n108, Z => n105);
   U838 : NAND3_X1 port map( A1 => n859, A2 => n855, A3 => sig_bal_delay, ZN =>
                           n97);
   U839 : NAND3_X1 port map( A1 => sig_bal_delay, A2 => n859, A3 => n8, ZN => 
                           n130_port);
   U840 : NAND3_X1 port map( A1 => sig_bal_delay, A2 => n855, A3 => n4, ZN => 
                           n131_port);
   U841 : NAND3_X1 port map( A1 => n200, A2 => n858, A3 => n34, ZN => n98);
   U842 : NAND3_X1 port map( A1 => n800, A2 => n858, A3 => n34, ZN => n121);
   U843 : NAND3_X1 port map( A1 => n34, A2 => n200, A3 => n5, ZN => n122);
   U844 : NAND3_X1 port map( A1 => n34, A2 => n800, A3 => n5, ZN => n123);
   U845 : NAND3_X1 port map( A1 => n853, A2 => n858, A3 => n200, ZN => n124);
   U846 : NAND3_X1 port map( A1 => n853, A2 => n858, A3 => n800, ZN => 
                           n125_port);
   U847 : NAND3_X1 port map( A1 => n200, A2 => n853, A3 => n5, ZN => n126_port)
                           ;
   U848 : NAND3_X1 port map( A1 => n8, A2 => sig_bal_delay, A3 => n4, ZN => 
                           n132_port);
   U849 : NAND3_X1 port map( A1 => n800, A2 => n853, A3 => n5, ZN => n127_port)
                           ;
   U3 : AND4_X1 port map( A1 => n680, A2 => n681, A3 => n682, A4 => n683, ZN =>
                           n918);
   U4 : BUF_X2 port map( A => n245, Z => n1028);
   U5 : BUF_X2 port map( A => n230, Z => n1060);
   U6 : BUF_X2 port map( A => n241, Z => n1039);
   U7 : BUF_X1 port map( A => n246, Z => n1024);
   U8 : BUF_X1 port map( A => n241, Z => n1040);
   U9 : BUF_X2 port map( A => n239, Z => n1045);
   U10 : BUF_X2 port map( A => n245, Z => n1027);
   U11 : AND4_X1 port map( A1 => n692, A2 => n693, A3 => n694, A4 => n695, ZN 
                           => n919);
   U12 : AND4_X1 port map( A1 => n684, A2 => n685, A3 => n686, A4 => n687, ZN 
                           => n916);
   U13 : AND4_X1 port map( A1 => n771, A2 => n770, A3 => n769, A4 => n772, ZN 
                           => n1005);
   U14 : NOR2_X1 port map( A1 => n94, A2 => n856, ZN => sig_bpw);
   U15 : AND4_X1 port map( A1 => n562, A2 => n563, A3 => n564, A4 => n565, ZN 
                           => n901);
   U16 : AND4_X1 port map( A1 => n582, A2 => n583, A3 => n584, A4 => n585, ZN 
                           => n914);
   U17 : INV_X1 port map( A => n898, ZN => n147_port);
   U18 : AND4_X1 port map( A1 => n805, A2 => n806, A3 => n807, A4 => n808, ZN 
                           => n896);
   U19 : AND4_X1 port map( A1 => n801, A2 => n802, A3 => n803, A4 => n804, ZN 
                           => n897);
   U20 : BUF_X1 port map( A => n1291, Z => n961);
   U21 : CLKBUF_X1 port map( A => sig_brt_port, Z => n797);
   U22 : CLKBUF_X1 port map( A => n208, Z => n798);
   U23 : BUF_X1 port map( A => n1308, Z => n1306);
   U24 : AND4_X1 port map( A1 => n248, A2 => n1002, A3 => n250, A4 => n251, ZN 
                           => n852);
   U25 : AND3_X1 port map( A1 => n250, A2 => n251, A3 => n248, ZN => n857);
   U26 : BUF_X1 port map( A => n204, Z => n1103);
   U27 : BUF_X1 port map( A => n203, Z => n861);
   U28 : AND4_X1 port map( A1 => n558, A2 => n559, A3 => n560, A4 => n561, ZN 
                           => n902);
   U29 : BUF_X2 port map( A => n243, Z => n1034);
   U30 : BUF_X1 port map( A => n220, Z => n1019);
   U31 : BUF_X2 port map( A => n230, Z => n1061);
   U32 : BUF_X1 port map( A => n230, Z => n1062);
   U33 : BUF_X1 port map( A => n203, Z => n1015);
   U34 : BUF_X2 port map( A => n201, Z => n1109);
   U35 : CLKBUF_X1 port map( A => n208, Z => n862);
   U36 : CLKBUF_X1 port map( A => n208, Z => n863);
   U37 : BUF_X1 port map( A => n203, Z => n1014);
   U38 : BUF_X1 port map( A => n203, Z => n1105);
   U39 : NOR2_X1 port map( A1 => n864, A2 => addr(4), ZN => n829);
   U40 : INV_X1 port map( A => addr(3), ZN => n864);
   U41 : BUF_X1 port map( A => n203, Z => n865);
   U42 : CLKBUF_X1 port map( A => n470, Z => n866);
   U43 : BUF_X1 port map( A => n216, Z => n868);
   U44 : BUF_X1 port map( A => n216, Z => n867);
   U45 : BUF_X1 port map( A => n205, Z => n1100);
   U46 : BUF_X1 port map( A => n208, Z => n869);
   U47 : BUF_X1 port map( A => n234, Z => n1048);
   U48 : CLKBUF_X1 port map( A => n208, Z => n870);
   U49 : OR4_X2 port map( A1 => n636, A2 => n637, A3 => n638, A4 => n639, ZN =>
                           n165);
   U50 : AND2_X1 port map( A1 => n825, A2 => n829, ZN => n205);
   U51 : BUF_X1 port map( A => n242, Z => n1037);
   U52 : CLKBUF_X1 port map( A => n208, Z => n871);
   U53 : CLKBUF_X1 port map( A => n1099, Z => n872);
   U54 : AND2_X1 port map( A1 => n828, A2 => n849, ZN => n242);
   U55 : BUF_X2 port map( A => n220, Z => n1080);
   U56 : BUF_X2 port map( A => n218, Z => n1081);
   U57 : BUF_X2 port map( A => n234, Z => n1049);
   U58 : AND3_X1 port map( A1 => n888, A2 => n966, A3 => addr(6), ZN => n827);
   U59 : AND2_X1 port map( A1 => n827, A2 => n828, ZN => n201);
   U60 : AND2_X1 port map( A1 => n827, A2 => n826, ZN => n198);
   U61 : AND2_X1 port map( A1 => n827, A2 => n829, ZN => n204);
   U62 : BUF_X2 port map( A => n220, Z => n1079);
   U63 : AND4_X2 port map( A1 => n762, A2 => n763, A3 => n761, A4 => n764, ZN 
                           => n1007);
   U64 : BUF_X2 port map( A => n241, Z => n1041);
   U65 : AND2_X2 port map( A1 => n825, A2 => n828, ZN => n203);
   U66 : CLKBUF_X1 port map( A => n145_port, Z => n873);
   U67 : BUF_X2 port map( A => n204, Z => n875);
   U68 : BUF_X1 port map( A => n204, Z => n874);
   U69 : BUF_X1 port map( A => n204, Z => n1102);
   U70 : BUF_X2 port map( A => n205, Z => n1101);
   U71 : BUF_X2 port map( A => n217, Z => n1084);
   U72 : BUF_X2 port map( A => n242, Z => n876);
   U73 : CLKBUF_X1 port map( A => n471, Z => n877);
   U74 : BUF_X2 port map( A => n198, Z => n1111);
   U75 : BUF_X2 port map( A => n227, Z => n1069);
   U76 : BUF_X2 port map( A => n215, Z => n1090);
   U77 : BUF_X2 port map( A => n246, Z => n1026);
   U78 : BUF_X2 port map( A => n246, Z => n1025);
   U79 : BUF_X2 port map( A => n243, Z => n1033);
   U80 : BUF_X2 port map( A => n206, Z => n1096);
   U81 : AND2_X4 port map( A1 => n825, A2 => n830, ZN => n208);
   U82 : AND3_X2 port map( A1 => n966, A2 => n831, A3 => addr(6), ZN => n825);
   U83 : NAND4_X1 port map( A1 => n1004, A2 => n1005, A3 => n1006, A4 => n1007,
                           ZN => n878);
   U84 : BUF_X2 port map( A => n244, Z => n1031);
   U85 : AND4_X1 port map( A1 => n879, A2 => n880, A3 => n881, A4 => n882, ZN 
                           => n185);
   U86 : AND4_X1 port map( A1 => n529, A2 => n530, A3 => n531, A4 => n532, ZN 
                           => n879);
   U87 : AND4_X1 port map( A1 => n525, A2 => n526, A3 => n527, A4 => n528, ZN 
                           => n880);
   U88 : AND4_X1 port map( A1 => n521, A2 => n522, A3 => n523, A4 => n524, ZN 
                           => n881);
   U89 : AND4_X1 port map( A1 => n517, A2 => n518, A3 => n519, A4 => n520, ZN 
                           => n882);
   U90 : BUF_X2 port map( A => n228, Z => n1067);
   U91 : AND4_X1 port map( A1 => n883, A2 => n884, A3 => n885, A4 => n886, ZN 
                           => n188_port);
   U92 : AND4_X1 port map( A1 => n549, A2 => n550, A3 => n551, A4 => n552, ZN 
                           => n883);
   U93 : AND4_X1 port map( A1 => n545, A2 => n546, A3 => n547, A4 => n548, ZN 
                           => n884);
   U94 : AND4_X1 port map( A1 => n541, A2 => n542, A3 => n543, A4 => n544, ZN 
                           => n885);
   U95 : AND4_X1 port map( A1 => n537, A2 => n538, A3 => n539, A4 => n540, ZN 
                           => n886);
   U96 : NAND4_X1 port map( A1 => n971, A2 => n972, A3 => n973, A4 => n974, ZN 
                           => n887);
   U97 : CLKBUF_X1 port map( A => addr(2), Z => n888);
   U98 : AOI211_X2 port map( C1 => n147_port, C2 => n268, A => n269, B => n270,
                           ZN => n250);
   U99 : OR4_X1 port map( A1 => n877, A2 => n866, A3 => n468, A4 => n469, ZN =>
                           n889);
   U100 : OR4_X2 port map( A1 => n656, A2 => n657, A3 => n658, A4 => n659, ZN 
                           => n167);
   U101 : BUF_X2 port map( A => n240, Z => n1043);
   U102 : BUF_X2 port map( A => n239, Z => n1046);
   U103 : NAND4_X1 port map( A1 => n890, A2 => n891, A3 => n892, A4 => n893, ZN
                           => n181);
   U104 : AND4_X1 port map( A1 => n732, A2 => n733, A3 => n734, A4 => n735, ZN 
                           => n890);
   U105 : AND4_X1 port map( A1 => n728, A2 => n729, A3 => n730, A4 => n731, ZN 
                           => n891);
   U106 : AND4_X1 port map( A1 => n724, A2 => n725, A3 => n726, A4 => n727, ZN 
                           => n892);
   U107 : AND4_X1 port map( A1 => n720, A2 => n721, A3 => n722, A4 => n723, ZN 
                           => n893);
   U108 : OR4_X2 port map( A1 => n616, A2 => n619, A3 => n618, A4 => n617, ZN 
                           => n175);
   U109 : OR4_X2 port map( A1 => n736, A2 => n737, A3 => n738, A4 => n739, ZN 
                           => n946);
   U110 : BUF_X2 port map( A => n233, Z => n1052);
   U111 : NAND4_X1 port map( A1 => n894, A2 => n895, A3 => n896, A4 => n897, ZN
                           => n139_port);
   U112 : AND4_X1 port map( A1 => n813, A2 => n814, A3 => n815, A4 => n816, ZN 
                           => n894);
   U113 : AND4_X1 port map( A1 => n809, A2 => n810, A3 => n811, A4 => n812, ZN 
                           => n895);
   U114 : BUF_X2 port map( A => n217, Z => n1085);
   U115 : BUF_X2 port map( A => n198, Z => n1110);
   U116 : NAND4_X1 port map( A1 => n979, A2 => n980, A3 => n981, A4 => n982, ZN
                           => n898);
   U117 : NAND4_X1 port map( A1 => n899, A2 => n900, A3 => n901, A4 => n902, ZN
                           => n183);
   U118 : AND4_X1 port map( A1 => n570, A2 => n571, A3 => n572, A4 => n573, ZN 
                           => n899);
   U119 : AND4_X1 port map( A1 => n566, A2 => n567, A3 => n568, A4 => n569, ZN 
                           => n900);
   U120 : NAND4_X1 port map( A1 => n903, A2 => n904, A3 => n905, A4 => n906, ZN
                           => n157);
   U121 : AND4_X1 port map( A1 => n363, A2 => n364, A3 => n365, A4 => n366, ZN 
                           => n903);
   U122 : AND4_X1 port map( A1 => n359, A2 => n360, A3 => n361, A4 => n362, ZN 
                           => n904);
   U123 : AND4_X1 port map( A1 => n351, A2 => n352, A3 => n354, A4 => n353, ZN 
                           => n905);
   U124 : AND4_X1 port map( A1 => n355, A2 => n356, A3 => n357, A4 => n358, ZN 
                           => n906);
   U125 : OAI222_X1 port map( A1 => n265, A2 => n155, B1 => n266, B2 => n159, 
                           C1 => n267, C2 => n157, ZN => n252);
   U126 : BUF_X2 port map( A => n244, Z => n1030);
   U127 : INV_X1 port map( A => n1001, ZN => n907);
   U128 : NAND4_X1 port map( A1 => n908, A2 => n909, A3 => n910, A4 => n911, ZN
                           => n159);
   U129 : AND4_X1 port map( A1 => n384, A2 => n385, A3 => n386, A4 => n387, ZN 
                           => n908);
   U130 : AND4_X1 port map( A1 => n380, A2 => n381, A3 => n382, A4 => n383, ZN 
                           => n909);
   U131 : AND4_X1 port map( A1 => n376, A2 => n377, A3 => n378, A4 => n379, ZN 
                           => n910);
   U132 : AND4_X1 port map( A1 => n372, A2 => n373, A3 => n374, A4 => n375, ZN 
                           => n911);
   U133 : BUF_X2 port map( A => n232, Z => n1055);
   U134 : BUF_X2 port map( A => n231, Z => n1058);
   U135 : BUF_X2 port map( A => n240, Z => n1042);
   U136 : NAND4_X1 port map( A1 => n912, A2 => n913, A3 => n914, A4 => n915, ZN
                           => n179);
   U137 : AND4_X1 port map( A1 => n590, A2 => n591, A3 => n592, A4 => n593, ZN 
                           => n912);
   U138 : AND4_X1 port map( A1 => n578, A2 => n579, A3 => n580, A4 => n581, ZN 
                           => n913);
   U139 : AND4_X1 port map( A1 => n586, A2 => n587, A3 => n588, A4 => n589, ZN 
                           => n915);
   U140 : AND4_X2 port map( A1 => n916, A2 => n917, A3 => n918, A4 => n919, ZN 
                           => n281);
   U141 : AND4_X1 port map( A1 => n688, A2 => n689, A3 => n690, A4 => n691, ZN 
                           => n917);
   U142 : OAI222_X1 port map( A1 => n262, A2 => n181, B1 => n263, B2 => n179, 
                           C1 => n264, C2 => n183, ZN => n253);
   U143 : BUF_X2 port map( A => n227, Z => n1070);
   U144 : BUF_X2 port map( A => n231, Z => n1057);
   U145 : BUF_X2 port map( A => n232, Z => n1054);
   U146 : AND2_X1 port map( A1 => n1002, A2 => n920, ZN => N126);
   U147 : NOR2_X1 port map( A1 => n936, A2 => n189, ZN => n920);
   U148 : BUF_X2 port map( A => n201, Z => n1108);
   U149 : NAND4_X1 port map( A1 => n921, A2 => n922, A3 => n923, A4 => n924, ZN
                           => n155);
   U150 : AND4_X1 port map( A1 => n343, A2 => n344, A3 => n345, A4 => n346, ZN 
                           => n921);
   U151 : AND4_X1 port map( A1 => n339, A2 => n341, A3 => n340, A4 => n342, ZN 
                           => n922);
   U152 : AND4_X1 port map( A1 => n335, A2 => n336, A3 => n337, A4 => n338, ZN 
                           => n923);
   U153 : AND4_X1 port map( A1 => n333, A2 => n332, A3 => n331, A4 => n334, ZN 
                           => n924);
   U154 : BUF_X2 port map( A => n228, Z => n1066);
   U155 : BUF_X2 port map( A => n233, Z => n1051);
   U156 : NAND4_X1 port map( A1 => n925, A2 => n926, A3 => n927, A4 => n928, ZN
                           => n161);
   U157 : AND4_X1 port map( A1 => n404, A2 => n405, A3 => n406, A4 => n407, ZN 
                           => n925);
   U158 : AND4_X1 port map( A1 => n400, A2 => n401, A3 => n402, A4 => n403, ZN 
                           => n926);
   U159 : AND4_X1 port map( A1 => n396, A2 => n397, A3 => n398, A4 => n399, ZN 
                           => n927);
   U160 : AND4_X1 port map( A1 => n392, A2 => n393, A3 => n394, A4 => n395, ZN 
                           => n928);
   U161 : INV_X1 port map( A => addr(2), ZN => n929);
   U162 : AND2_X1 port map( A1 => bht_17_6_port, A2 => n1096, ZN => n930);
   U163 : AND2_X1 port map( A1 => n208, A2 => bht_16_6_port, ZN => n931);
   U164 : NOR2_X1 port map( A1 => n930, A2 => n931, ZN => n578);
   U165 : BUF_X2 port map( A => n206, Z => n1097);
   U166 : OR4_X2 port map( A1 => n468, A2 => n469, A3 => n470, A4 => n471, ZN 
                           => n153);
   U167 : OAI222_X1 port map( A1 => n273, A2 => n887, B1 => n274, B2 => 
                           n141_port, C1 => n275, C2 => n889, ZN => n269);
   U168 : BUF_X2 port map( A => n220, Z => n1018);
   U169 : BUF_X2 port map( A => n218, Z => n1082);
   U170 : NAND4_X1 port map( A1 => n932, A2 => n933, A3 => n934, A4 => n935, ZN
                           => n141_port);
   U171 : AND4_X1 port map( A1 => n506, A2 => n507, A3 => n508, A4 => n509, ZN 
                           => n932);
   U172 : AND4_X1 port map( A1 => n502, A2 => n503, A3 => n504, A4 => n505, ZN 
                           => n933);
   U173 : AND4_X1 port map( A1 => n498, A2 => n499, A3 => n500, A4 => n501, ZN 
                           => n934);
   U174 : AND4_X1 port map( A1 => n496, A2 => n494, A3 => n495, A4 => n497, ZN 
                           => n935);
   U175 : BUF_X2 port map( A => n215, Z => n1091);
   U176 : NAND3_X1 port map( A1 => n251, A2 => n250, A3 => n248, ZN => n936);
   U177 : NOR4_X2 port map( A1 => n252, A2 => n253, A3 => n255, A4 => n254, ZN 
                           => n251);
   U178 : AND2_X1 port map( A1 => n262, A2 => n181, ZN => n937);
   U179 : AND2_X1 port map( A1 => n256, A2 => n163, ZN => n938);
   U180 : AND2_X1 port map( A1 => n283, A2 => n171, ZN => n939);
   U181 : NOR3_X1 port map( A1 => n937, A2 => n938, A3 => n939, ZN => n299);
   U182 : OR4_X2 port map( A1 => n696, A2 => n697, A3 => n698, A4 => n699, ZN 
                           => n163);
   U183 : CLKBUF_X1 port map( A => n1062, Z => n965);
   U184 : BUF_X2 port map( A => n229, Z => n1064);
   U185 : AND3_X1 port map( A1 => n940, A2 => n941, A3 => n942, ZN => n304);
   U186 : NAND2_X1 port map( A1 => n153, A2 => n275, ZN => n940);
   U187 : NAND2_X1 port map( A1 => n151_port, A2 => n273, ZN => n941);
   U188 : NAND2_X1 port map( A1 => n149_port, A2 => n272, ZN => n942);
   U189 : BUF_X2 port map( A => n201, Z => n1107);
   U190 : NAND2_X1 port map( A1 => n157, A2 => n267, ZN => n943);
   U191 : NAND2_X1 port map( A1 => n155, A2 => n265, ZN => n944);
   U192 : NAND2_X1 port map( A1 => n169, A2 => n259, ZN => n945);
   U193 : AND3_X1 port map( A1 => n943, A2 => n944, A3 => n945, ZN => n306);
   U194 : BUF_X2 port map( A => n229, Z => n1063);
   U195 : BUF_X2 port map( A => n217, Z => n1086);
   U196 : BUF_X2 port map( A => n205, Z => n1099);
   U197 : BUF_X2 port map( A => n242, Z => n1036);
   U198 : CLKBUF_X1 port map( A => n1291, Z => n962);
   U199 : BUF_X1 port map( A => n852, Z => n955);
   U200 : BUF_X1 port map( A => n852, Z => n956);
   U201 : BUF_X1 port map( A => n852, Z => n957);
   U202 : BUF_X1 port map( A => n852, Z => n959);
   U203 : BUF_X1 port map( A => n852, Z => n958);
   U204 : BUF_X1 port map( A => n955, Z => n960);
   U205 : BUF_X1 port map( A => N188, Z => n1291);
   U206 : CLKBUF_X1 port map( A => N188, Z => n1292);
   U207 : BUF_X1 port map( A => n221, Z => n1076);
   U208 : BUF_X1 port map( A => n216, Z => n1088);
   U209 : NOR2_X1 port map( A1 => n1306, A2 => n1293, ZN => N188);
   U210 : BUF_X1 port map( A => n221, Z => n1075);
   U211 : BUF_X1 port map( A => n222, Z => n1072);
   U212 : BUF_X1 port map( A => n216, Z => n1087);
   U213 : BUF_X1 port map( A => n213, Z => n1094);
   U214 : BUF_X1 port map( A => n213, Z => n1093);
   U215 : BUF_X1 port map( A => n222, Z => n1074);
   U216 : BUF_X1 port map( A => n222, Z => n1008);
   U217 : CLKBUF_X1 port map( A => n244, Z => n1032);
   U218 : BUF_X1 port map( A => n222, Z => n1009);
   U219 : CLKBUF_X1 port map( A => n233, Z => n1053);
   U220 : CLKBUF_X1 port map( A => n245, Z => n1029);
   U221 : CLKBUF_X1 port map( A => n243, Z => n1035);
   U222 : CLKBUF_X1 port map( A => n227, Z => n1071);
   U223 : CLKBUF_X1 port map( A => n239, Z => n1047);
   U224 : CLKBUF_X1 port map( A => n228, Z => n1068);
   U225 : CLKBUF_X1 port map( A => n231, Z => n1059);
   U226 : CLKBUF_X1 port map( A => n234, Z => n1050);
   U227 : CLKBUF_X1 port map( A => n240, Z => n1044);
   U228 : CLKBUF_X1 port map( A => n232, Z => n1056);
   U229 : CLKBUF_X1 port map( A => n229, Z => n1065);
   U230 : CLKBUF_X1 port map( A => n242, Z => n1038);
   U231 : CLKBUF_X1 port map( A => n198, Z => n1112);
   U232 : CLKBUF_X1 port map( A => n218, Z => n1083);
   U233 : CLKBUF_X1 port map( A => n221, Z => n1077);
   U234 : CLKBUF_X1 port map( A => n206, Z => n1098);
   U235 : CLKBUF_X1 port map( A => n216, Z => n1089);
   U236 : CLKBUF_X1 port map( A => n213, Z => n1095);
   U237 : BUF_X1 port map( A => N3730, Z => n1198);
   U238 : BUF_X1 port map( A => N3622, Z => n1204);
   U239 : BUF_X1 port map( A => N3514, Z => n1210);
   U240 : BUF_X1 port map( A => N3406, Z => n1216);
   U241 : BUF_X1 port map( A => N3460, Z => n1213);
   U242 : BUF_X1 port map( A => N3568, Z => n1207);
   U243 : BUF_X1 port map( A => N3676, Z => n1201);
   U244 : BUF_X1 port map( A => N3784, Z => n1117);
   U245 : BUF_X1 port map( A => N3730, Z => n1199);
   U246 : BUF_X1 port map( A => N3622, Z => n1205);
   U247 : BUF_X1 port map( A => N3514, Z => n1211);
   U248 : BUF_X1 port map( A => N3406, Z => n1217);
   U249 : BUF_X1 port map( A => N3460, Z => n1214);
   U250 : BUF_X1 port map( A => N3568, Z => n1208);
   U251 : BUF_X1 port map( A => N3676, Z => n1202);
   U252 : BUF_X1 port map( A => N3784, Z => n1118);
   U253 : BUF_X1 port map( A => N3298, Z => n1222);
   U254 : BUF_X1 port map( A => N3190, Z => n1228);
   U255 : BUF_X1 port map( A => N3082, Z => n1234);
   U256 : BUF_X1 port map( A => N2974, Z => n1240);
   U257 : BUF_X1 port map( A => N2866, Z => n1246);
   U258 : BUF_X1 port map( A => N2758, Z => n1252);
   U259 : BUF_X1 port map( A => N2650, Z => n1258);
   U260 : BUF_X1 port map( A => N2542, Z => n1264);
   U261 : BUF_X1 port map( A => N2434, Z => n1270);
   U262 : BUF_X1 port map( A => N2326, Z => n1276);
   U263 : BUF_X1 port map( A => N2218, Z => n1282);
   U264 : BUF_X1 port map( A => N2110, Z => n1288);
   U265 : BUF_X1 port map( A => N2164, Z => n1285);
   U266 : BUF_X1 port map( A => N2272, Z => n1279);
   U267 : BUF_X1 port map( A => N2380, Z => n1273);
   U268 : BUF_X1 port map( A => N2488, Z => n1267);
   U269 : BUF_X1 port map( A => N2596, Z => n1261);
   U270 : BUF_X1 port map( A => N2704, Z => n1255);
   U271 : BUF_X1 port map( A => N2812, Z => n1249);
   U272 : BUF_X1 port map( A => N2920, Z => n1243);
   U273 : BUF_X1 port map( A => N3028, Z => n1237);
   U274 : BUF_X1 port map( A => N3136, Z => n1231);
   U275 : BUF_X1 port map( A => N3244, Z => n1225);
   U276 : BUF_X1 port map( A => N3352, Z => n1219);
   U277 : BUF_X1 port map( A => N3298, Z => n1223);
   U278 : BUF_X1 port map( A => N3190, Z => n1229);
   U279 : BUF_X1 port map( A => N3082, Z => n1235);
   U280 : BUF_X1 port map( A => N2974, Z => n1241);
   U281 : BUF_X1 port map( A => N2866, Z => n1247);
   U282 : BUF_X1 port map( A => N2758, Z => n1253);
   U283 : BUF_X1 port map( A => N2650, Z => n1259);
   U284 : BUF_X1 port map( A => N2542, Z => n1265);
   U285 : BUF_X1 port map( A => N2434, Z => n1271);
   U286 : BUF_X1 port map( A => N2326, Z => n1277);
   U287 : BUF_X1 port map( A => N2218, Z => n1283);
   U288 : BUF_X1 port map( A => N2110, Z => n1289);
   U289 : BUF_X1 port map( A => N2164, Z => n1286);
   U290 : BUF_X1 port map( A => N2272, Z => n1280);
   U291 : BUF_X1 port map( A => N2380, Z => n1274);
   U292 : BUF_X1 port map( A => N2488, Z => n1268);
   U293 : BUF_X1 port map( A => N2596, Z => n1262);
   U294 : BUF_X1 port map( A => N2704, Z => n1256);
   U295 : BUF_X1 port map( A => N2812, Z => n1250);
   U296 : BUF_X1 port map( A => N2920, Z => n1244);
   U297 : BUF_X1 port map( A => N3028, Z => n1238);
   U298 : BUF_X1 port map( A => N3136, Z => n1232);
   U299 : BUF_X1 port map( A => N3244, Z => n1226);
   U300 : BUF_X1 port map( A => N3352, Z => n1220);
   U301 : BUF_X1 port map( A => N3735, Z => n1192);
   U302 : BUF_X1 port map( A => N3735, Z => n1193);
   U303 : BUF_X1 port map( A => N3735, Z => n1194);
   U304 : BUF_X1 port map( A => N3730, Z => n1200);
   U305 : BUF_X1 port map( A => N3622, Z => n1206);
   U306 : BUF_X1 port map( A => N3514, Z => n1212);
   U307 : BUF_X1 port map( A => N3406, Z => n1218);
   U308 : BUF_X1 port map( A => N3460, Z => n1215);
   U309 : BUF_X1 port map( A => N3568, Z => n1209);
   U310 : BUF_X1 port map( A => N3676, Z => n1203);
   U311 : BUF_X1 port map( A => N3784, Z => n1119);
   U312 : BUF_X1 port map( A => N3298, Z => n1224);
   U313 : BUF_X1 port map( A => N3190, Z => n1230);
   U314 : BUF_X1 port map( A => N3082, Z => n1236);
   U315 : BUF_X1 port map( A => N2974, Z => n1242);
   U316 : BUF_X1 port map( A => N2866, Z => n1248);
   U317 : BUF_X1 port map( A => N2758, Z => n1254);
   U318 : BUF_X1 port map( A => N2650, Z => n1260);
   U319 : BUF_X1 port map( A => N2542, Z => n1266);
   U320 : BUF_X1 port map( A => N2434, Z => n1272);
   U321 : BUF_X1 port map( A => N2326, Z => n1278);
   U322 : BUF_X1 port map( A => N2218, Z => n1284);
   U323 : BUF_X1 port map( A => N2164, Z => n1287);
   U324 : BUF_X1 port map( A => N2272, Z => n1281);
   U325 : BUF_X1 port map( A => N2380, Z => n1275);
   U326 : BUF_X1 port map( A => N2488, Z => n1269);
   U327 : BUF_X1 port map( A => N2596, Z => n1263);
   U328 : BUF_X1 port map( A => N2704, Z => n1257);
   U329 : BUF_X1 port map( A => N2812, Z => n1251);
   U330 : BUF_X1 port map( A => N2920, Z => n1245);
   U331 : BUF_X1 port map( A => N3028, Z => n1239);
   U332 : BUF_X1 port map( A => N3136, Z => n1233);
   U333 : BUF_X1 port map( A => N3244, Z => n1227);
   U334 : BUF_X1 port map( A => N3352, Z => n1221);
   U335 : BUF_X1 port map( A => N2110, Z => n1290);
   U336 : NOR4_X1 port map( A1 => n288, A2 => n289, A3 => n290, A4 => n291, ZN 
                           => n287);
   U337 : NAND4_X1 port map( A1 => n272, A2 => n274, A3 => n293, A4 => n294, ZN
                           => n288);
   U338 : NAND4_X1 port map( A1 => n263, A2 => n292, A3 => n275, A4 => n271, ZN
                           => n289);
   U339 : NAND4_X1 port map( A1 => n259, A2 => n260, A3 => n264, A4 => n262, ZN
                           => n290);
   U340 : AND4_X1 port map( A1 => n793, A2 => n794, A3 => n795, A4 => n796, ZN 
                           => n994);
   U341 : AND4_X1 port map( A1 => n781, A2 => n782, A3 => n783, A4 => n784, ZN 
                           => n997);
   U342 : AND4_X1 port map( A1 => n604, A2 => n605, A3 => n606, A4 => n607, ZN 
                           => n969);
   U343 : AND4_X1 port map( A1 => n436, A2 => n437, A3 => n438, A4 => n439, ZN 
                           => n977);
   U344 : AND4_X1 port map( A1 => n432, A2 => n433, A3 => n434, A4 => n435, ZN 
                           => n978);
   U345 : AND4_X1 port map( A1 => n464, A2 => n465, A3 => n466, A4 => n467, ZN 
                           => n971);
   U346 : NOR4_X1 port map( A1 => n190, A2 => n191, A3 => n192, A4 => n193, ZN 
                           => n189);
   U347 : NAND4_X1 port map( A1 => n235, A2 => n236, A3 => n237, A4 => n238, ZN
                           => n190);
   U348 : NAND2_X1 port map( A1 => rst, A2 => n100, ZN => n94);
   U349 : NAND4_X1 port map( A1 => n258, A2 => n256, A3 => n257, A4 => n261, ZN
                           => n291);
   U350 : NAND4_X1 port map( A1 => n632, A2 => n633, A3 => n634, A4 => n635, ZN
                           => n616);
   U351 : NAND4_X1 port map( A1 => n712, A2 => n713, A3 => n714, A4 => n715, ZN
                           => n696);
   U352 : NAND4_X1 port map( A1 => n708, A2 => n709, A3 => n710, A4 => n711, ZN
                           => n697);
   U353 : NAND4_X1 port map( A1 => n672, A2 => n673, A3 => n674, A4 => n675, ZN
                           => n656);
   U354 : NAND4_X1 port map( A1 => n664, A2 => n665, A3 => n666, A4 => n667, ZN
                           => n658);
   U355 : NAND4_X1 port map( A1 => n668, A2 => n669, A3 => n670, A4 => n671, ZN
                           => n657);
   U356 : NAND4_X1 port map( A1 => n652, A2 => n653, A3 => n654, A4 => n655, ZN
                           => n636);
   U357 : NAND4_X1 port map( A1 => n640, A2 => n641, A3 => n642, A4 => n643, ZN
                           => n639);
   U358 : AND2_X1 port map( A1 => n837, A2 => n829, ZN => n220);
   U359 : AND2_X1 port map( A1 => n837, A2 => n830, ZN => n222);
   U360 : AND2_X1 port map( A1 => n849, A2 => n829, ZN => n244);
   U361 : AND2_X1 port map( A1 => n826, A2 => n838, ZN => n213);
   U362 : AND2_X1 port map( A1 => n830, A2 => n838, ZN => n221);
   U363 : AND2_X1 port map( A1 => n829, A2 => n838, ZN => n218);
   U364 : AND3_X1 port map( A1 => n489, A2 => n948, A3 => n947, ZN => n303);
   U365 : NAND2_X1 port map( A1 => n139_port, A2 => n292, ZN => n947);
   U366 : NAND2_X1 port map( A1 => n141_port, A2 => n274, ZN => n948);
   U367 : AND3_X1 port map( A1 => n949, A2 => n950, A3 => n595, ZN => n300);
   U368 : NAND2_X1 port map( A1 => n260, A2 => n167, ZN => n949);
   U369 : NAND2_X1 port map( A1 => n261, A2 => n165, ZN => n950);
   U370 : AND4_X1 port map( A1 => n276, A2 => n298, A3 => n283, A4 => n273, ZN 
                           => n284);
   U371 : INV_X1 port map( A => n276, ZN => n268);
   U372 : INV_X1 port map( A => n1295, ZN => n1293);
   U373 : OAI22_X1 port map( A1 => n94, A2 => n860, B1 => n100, B2 => n101, ZN 
                           => N3735);
   U374 : NAND2_X1 port map( A1 => rst, A2 => n854, ZN => n101);
   U375 : OAI21_X1 port map( B1 => n97, B2 => n121, A => rst, ZN => N3730);
   U376 : OAI21_X1 port map( B1 => n97, B2 => n123, A => rst, ZN => N3622);
   U377 : OAI21_X1 port map( B1 => n97, B2 => n125_port, A => rst, ZN => N3514)
                           ;
   U378 : OAI21_X1 port map( B1 => n97, B2 => n127_port, A => rst, ZN => N3406)
                           ;
   U379 : OAI21_X1 port map( B1 => n97, B2 => n126_port, A => rst, ZN => N3460)
                           ;
   U380 : OAI21_X1 port map( B1 => n97, B2 => n124, A => rst, ZN => N3568);
   U381 : OAI21_X1 port map( B1 => n97, B2 => n122, A => rst, ZN => N3676);
   U382 : OAI21_X1 port map( B1 => n97, B2 => n98, A => rst, ZN => N3784);
   U383 : OAI21_X1 port map( B1 => n121, B2 => n130_port, A => rst, ZN => N3298
                           );
   U384 : OAI21_X1 port map( B1 => n123, B2 => n130_port, A => rst, ZN => N3190
                           );
   U385 : OAI21_X1 port map( B1 => n125_port, B2 => n130_port, A => rst, ZN => 
                           N3082);
   U386 : OAI21_X1 port map( B1 => n127_port, B2 => n130_port, A => rst, ZN => 
                           N2974);
   U387 : OAI21_X1 port map( B1 => n121, B2 => n131_port, A => rst, ZN => N2866
                           );
   U388 : OAI21_X1 port map( B1 => n123, B2 => n131_port, A => rst, ZN => N2758
                           );
   U389 : OAI21_X1 port map( B1 => n125_port, B2 => n131_port, A => rst, ZN => 
                           N2650);
   U390 : OAI21_X1 port map( B1 => n127_port, B2 => n131_port, A => rst, ZN => 
                           N2542);
   U391 : OAI21_X1 port map( B1 => n121, B2 => n132_port, A => rst, ZN => N2434
                           );
   U392 : OAI21_X1 port map( B1 => n123, B2 => n132_port, A => rst, ZN => N2326
                           );
   U393 : OAI21_X1 port map( B1 => n125_port, B2 => n132_port, A => rst, ZN => 
                           N2218);
   U394 : OAI21_X1 port map( B1 => n126_port, B2 => n132_port, A => rst, ZN => 
                           N2164);
   U395 : OAI21_X1 port map( B1 => n124, B2 => n132_port, A => rst, ZN => N2272
                           );
   U396 : OAI21_X1 port map( B1 => n122, B2 => n132_port, A => rst, ZN => N2380
                           );
   U397 : OAI21_X1 port map( B1 => n98, B2 => n132_port, A => rst, ZN => N2488)
                           ;
   U398 : OAI21_X1 port map( B1 => n126_port, B2 => n131_port, A => rst, ZN => 
                           N2596);
   U399 : OAI21_X1 port map( B1 => n124, B2 => n131_port, A => rst, ZN => N2704
                           );
   U400 : OAI21_X1 port map( B1 => n122, B2 => n131_port, A => rst, ZN => N2812
                           );
   U401 : OAI21_X1 port map( B1 => n98, B2 => n131_port, A => rst, ZN => N2920)
                           ;
   U402 : OAI21_X1 port map( B1 => n126_port, B2 => n130_port, A => rst, ZN => 
                           N3028);
   U403 : OAI21_X1 port map( B1 => n124, B2 => n130_port, A => rst, ZN => N3136
                           );
   U404 : OAI21_X1 port map( B1 => n122, B2 => n130_port, A => rst, ZN => N3244
                           );
   U405 : OAI21_X1 port map( B1 => n98, B2 => n130_port, A => rst, ZN => N3352)
                           ;
   U406 : OAI21_X1 port map( B1 => n127_port, B2 => n132_port, A => rst, ZN => 
                           N2110);
   U407 : NOR2_X1 port map( A1 => n247, A2 => n953, ZN => N125);
   U408 : NOR4_X1 port map( A1 => n817, A2 => n818, A3 => n819, A4 => n820, ZN 
                           => n247);
   U409 : NAND4_X1 port map( A1 => n845, A2 => n846, A3 => n847, A4 => n848, ZN
                           => n817);
   U410 : NAND4_X1 port map( A1 => n839, A2 => n840, A3 => n841, A4 => n842, ZN
                           => n818);
   U411 : BUF_X1 port map( A => N3733, Z => n1195);
   U412 : BUF_X1 port map( A => N3733, Z => n1196);
   U413 : BUF_X1 port map( A => N3737, Z => n1190);
   U414 : BUF_X1 port map( A => N3737, Z => n1189);
   U415 : BUF_X1 port map( A => N3783, Z => n1121);
   U416 : BUF_X1 port map( A => N3739, Z => n1187);
   U417 : BUF_X1 port map( A => N3739, Z => n1186);
   U418 : BUF_X1 port map( A => N3741, Z => n1184);
   U419 : BUF_X1 port map( A => N3741, Z => n1183);
   U420 : BUF_X1 port map( A => N3743, Z => n1181);
   U421 : BUF_X1 port map( A => N3743, Z => n1180);
   U422 : BUF_X1 port map( A => N3745, Z => n1178);
   U423 : BUF_X1 port map( A => N3745, Z => n1177);
   U424 : BUF_X1 port map( A => N3747, Z => n1175);
   U425 : BUF_X1 port map( A => N3747, Z => n1174);
   U426 : BUF_X1 port map( A => N3749, Z => n1172);
   U427 : BUF_X1 port map( A => N3749, Z => n1171);
   U428 : BUF_X1 port map( A => N3751, Z => n1169);
   U429 : BUF_X1 port map( A => N3751, Z => n1168);
   U430 : BUF_X1 port map( A => N3753, Z => n1166);
   U431 : BUF_X1 port map( A => N3753, Z => n1165);
   U432 : BUF_X1 port map( A => N3755, Z => n1163);
   U433 : BUF_X1 port map( A => N3755, Z => n1162);
   U434 : BUF_X1 port map( A => N3757, Z => n1160);
   U435 : BUF_X1 port map( A => N3757, Z => n1159);
   U436 : BUF_X1 port map( A => N3759, Z => n1157);
   U437 : BUF_X1 port map( A => N3759, Z => n1156);
   U438 : BUF_X1 port map( A => N3761, Z => n1154);
   U439 : BUF_X1 port map( A => N3761, Z => n1153);
   U440 : BUF_X1 port map( A => N3763, Z => n1151);
   U441 : BUF_X1 port map( A => N3763, Z => n1150);
   U442 : BUF_X1 port map( A => N3765, Z => n1148);
   U443 : BUF_X1 port map( A => N3765, Z => n1147);
   U444 : BUF_X1 port map( A => N3767, Z => n1145);
   U445 : BUF_X1 port map( A => N3767, Z => n1144);
   U446 : BUF_X1 port map( A => N3769, Z => n1142);
   U447 : BUF_X1 port map( A => N3769, Z => n1141);
   U448 : BUF_X1 port map( A => N3771, Z => n1139);
   U449 : BUF_X1 port map( A => N3771, Z => n1138);
   U450 : BUF_X1 port map( A => N3773, Z => n1136);
   U451 : BUF_X1 port map( A => N3773, Z => n1135);
   U452 : BUF_X1 port map( A => N3775, Z => n1133);
   U453 : BUF_X1 port map( A => N3775, Z => n1132);
   U454 : BUF_X1 port map( A => N3777, Z => n1130);
   U455 : BUF_X1 port map( A => N3777, Z => n1129);
   U456 : BUF_X1 port map( A => N3779, Z => n1127);
   U457 : BUF_X1 port map( A => N3779, Z => n1126);
   U458 : BUF_X1 port map( A => N3781, Z => n1124);
   U459 : BUF_X1 port map( A => N3781, Z => n1123);
   U460 : BUF_X1 port map( A => N3785, Z => n1115);
   U461 : BUF_X1 port map( A => N3785, Z => n1114);
   U462 : BUF_X1 port map( A => N3783, Z => n1120);
   U463 : BUF_X1 port map( A => n1307, Z => n1305);
   U464 : BUF_X1 port map( A => n1303, Z => n1304);
   U465 : BUF_X1 port map( A => n1307, Z => n1303);
   U466 : BUF_X1 port map( A => n1307, Z => n1302);
   U467 : BUF_X1 port map( A => n1307, Z => n1301);
   U468 : BUF_X1 port map( A => n1302, Z => n1300);
   U469 : BUF_X1 port map( A => N3733, Z => n1197);
   U470 : BUF_X1 port map( A => N3737, Z => n1191);
   U471 : BUF_X1 port map( A => N3783, Z => n1122);
   U472 : BUF_X1 port map( A => N3739, Z => n1188);
   U473 : BUF_X1 port map( A => N3741, Z => n1185);
   U474 : BUF_X1 port map( A => N3743, Z => n1182);
   U475 : BUF_X1 port map( A => N3745, Z => n1179);
   U476 : BUF_X1 port map( A => N3747, Z => n1176);
   U477 : BUF_X1 port map( A => N3749, Z => n1173);
   U478 : BUF_X1 port map( A => N3751, Z => n1170);
   U479 : BUF_X1 port map( A => N3753, Z => n1167);
   U480 : BUF_X1 port map( A => N3755, Z => n1164);
   U481 : BUF_X1 port map( A => N3757, Z => n1161);
   U482 : BUF_X1 port map( A => N3759, Z => n1158);
   U483 : BUF_X1 port map( A => N3761, Z => n1155);
   U484 : BUF_X1 port map( A => N3763, Z => n1152);
   U485 : BUF_X1 port map( A => N3765, Z => n1149);
   U486 : BUF_X1 port map( A => N3767, Z => n1146);
   U487 : BUF_X1 port map( A => N3769, Z => n1143);
   U488 : BUF_X1 port map( A => N3771, Z => n1140);
   U489 : BUF_X1 port map( A => N3773, Z => n1137);
   U490 : BUF_X1 port map( A => N3775, Z => n1134);
   U491 : BUF_X1 port map( A => N3777, Z => n1131);
   U492 : BUF_X1 port map( A => N3779, Z => n1128);
   U493 : BUF_X1 port map( A => N3781, Z => n1125);
   U494 : BUF_X1 port map( A => N3785, Z => n1116);
   U495 : CLKBUF_X1 port map( A => n1308, Z => n1307);
   U496 : NOR4_X1 port map( A1 => ld_a(23), A2 => ld_a(22), A3 => ld_a(21), A4 
                           => ld_a(20), ZN => n114);
   U497 : NOR4_X1 port map( A1 => ld_a(9), A2 => ld_a(8), A3 => ld_a(7), A4 => 
                           ld_a(6), ZN => n118);
   U498 : AOI22_X1 port map( A1 => n1293, A2 => reg_a(20), B1 => n1295, B2 => 
                           addr(27), ZN => n276);
   U499 : AOI22_X1 port map( A1 => n1293, A2 => reg_a(13), B1 => n1295, B2 => 
                           addr(20), ZN => n271);
   U500 : AOI22_X1 port map( A1 => n1293, A2 => reg_a(3), B1 => n1299, B2 => 
                           addr(10), ZN => n262);
   U501 : AOI22_X1 port map( A1 => n1293, A2 => reg_a(22), B1 => n1299, B2 => 
                           addr(29), ZN => n294);
   U502 : AOI22_X1 port map( A1 => n1293, A2 => reg_a(16), B1 => n1295, B2 => 
                           addr(23), ZN => n265);
   U503 : AOI22_X1 port map( A1 => n1293, A2 => reg_a(21), B1 => n1298, B2 => 
                           addr(28), ZN => n293);
   U504 : AOI22_X1 port map( A1 => n1293, A2 => reg_a(14), B1 => n1297, B2 => 
                           addr(21), ZN => n266);
   U505 : AOI22_X1 port map( A1 => n1293, A2 => reg_a(2), B1 => n1297, B2 => 
                           addr(9), ZN => n264);
   U506 : AOI22_X1 port map( A1 => n1293, A2 => reg_a(8), B1 => n1298, B2 => 
                           addr(15), ZN => n283);
   U507 : AOI22_X1 port map( A1 => n1293, A2 => reg_a(5), B1 => n1297, B2 => 
                           addr(12), ZN => n257);
   U508 : AOI22_X1 port map( A1 => n1293, A2 => reg_a(7), B1 => n1299, B2 => 
                           addr(14), ZN => n298);
   U509 : AOI22_X1 port map( A1 => n1293, A2 => reg_a(15), B1 => n1295, B2 => 
                           addr(22), ZN => n267);
   U510 : AOI22_X1 port map( A1 => n1293, A2 => reg_a(12), B1 => n1298, B2 => 
                           addr(19), ZN => n256);
   U511 : AOI22_X1 port map( A1 => n1293, A2 => reg_a(11), B1 => n1298, B2 => 
                           addr(18), ZN => n261);
   U512 : AOI22_X1 port map( A1 => n1293, A2 => reg_a(18), B1 => n1296, B2 => 
                           addr(25), ZN => n273);
   U513 : AOI22_X1 port map( A1 => n1293, A2 => reg_a(6), B1 => addr(13), B2 =>
                           n1294, ZN => n258);
   U514 : AOI22_X1 port map( A1 => n1293, A2 => reg_a(4), B1 => n1297, B2 => 
                           addr(11), ZN => n263);
   U515 : AOI22_X1 port map( A1 => n1293, A2 => reg_a(17), B1 => n1296, B2 => 
                           addr(24), ZN => n275);
   U516 : AOI22_X1 port map( A1 => n1293, A2 => reg_a(9), B1 => n1294, B2 => 
                           addr(16), ZN => n259);
   U517 : AOI22_X1 port map( A1 => n1293, A2 => reg_a(23), B1 => n1296, B2 => 
                           addr(30), ZN => n274);
   U518 : AOI22_X1 port map( A1 => n1293, A2 => reg_a(24), B1 => n1299, B2 => 
                           addr(31), ZN => n292);
   U519 : AOI22_X1 port map( A1 => n1293, A2 => reg_a(10), B1 => n1298, B2 => 
                           addr(17), ZN => n260);
   U520 : AOI22_X1 port map( A1 => n1293, A2 => reg_a(19), B1 => n1296, B2 => 
                           addr(26), ZN => n272);
   U521 : NAND4_X1 port map( A1 => opcd_delay_2_port, A2 => n214, A3 => n105, 
                           A4 => n106, ZN => n100);
   U522 : NOR3_X1 port map( A1 => opcd_delay_3_port, A2 => opcd_delay_5_port, 
                           A3 => opcd_delay_4_port, ZN => n106);
   U523 : NOR2_X1 port map( A1 => n109, A2 => n110, ZN => n108);
   U524 : AOI22_X1 port map( A1 => bht_7_2_port, A2 => n1070, B1 => 
                           bht_6_2_port, B2 => n1067, ZN => n540);
   U525 : AOI22_X1 port map( A1 => bht_15_26_port, A2 => n1047, B1 => 
                           bht_14_26_port, B2 => n1044, ZN => n808);
   U526 : AOI22_X1 port map( A1 => bht_7_14_port, A2 => n1070, B1 => 
                           bht_6_14_port, B2 => n1067, ZN => n711);
   U527 : AOI22_X1 port map( A1 => bht_7_12_port, A2 => n1070, B1 => 
                           bht_6_12_port, B2 => n1068, ZN => n671);
   U528 : AOI22_X1 port map( A1 => bht_7_5_port, A2 => n1070, B1 => 
                           bht_6_5_port, B2 => n1067, ZN => n731);
   U529 : AOI22_X1 port map( A1 => bht_5_26_port, A2 => n1064, B1 => 
                           bht_4_26_port, B2 => n1060, ZN => n803);
   U530 : AOI22_X1 port map( A1 => bht_13_26_port, A2 => n1039, B1 => 
                           bht_12_26_port, B2 => n1036, ZN => n807);
   U531 : AOI22_X1 port map( A1 => bht_11_26_port, A2 => n1035, B1 => 
                           bht_10_26_port, B2 => n1032, ZN => n806);
   U532 : AOI22_X1 port map( A1 => bht_1_14_port, A2 => n1052, B1 => 
                           bht_0_14_port, B2 => n1050, ZN => n708);
   U533 : AOI22_X1 port map( A1 => bht_1_12_port, A2 => n1052, B1 => 
                           bht_0_12_port, B2 => n1049, ZN => n668);
   U534 : AOI22_X1 port map( A1 => bht_1_5_port, A2 => n1052, B1 => 
                           bht_0_5_port, B2 => n1049, ZN => n728);
   U535 : AOI22_X1 port map( A1 => bht_1_17_port, A2 => n1051, B1 => 
                           bht_0_17_port, B2 => n1049, ZN => n351);
   U536 : AOI22_X1 port map( A1 => bht_1_3_port, A2 => n1051, B1 => 
                           bht_0_3_port, B2 => n1050, ZN => n517);
   U537 : AOI22_X1 port map( A1 => bht_9_2_port, A2 => n1028, B1 => 
                           bht_8_2_port, B2 => n1024, ZN => n541);
   U538 : AOI22_X1 port map( A1 => bht_9_26_port, A2 => n1029, B1 => 
                           bht_8_26_port, B2 => n1026, ZN => n805);
   U539 : AOI22_X1 port map( A1 => bht_9_8_port, A2 => n1028, B1 => 
                           bht_8_8_port, B2 => n1024, ZN => n632);
   U540 : AOI22_X1 port map( A1 => bht_9_6_port, A2 => n1028, B1 => 
                           bht_8_6_port, B2 => n1026, ZN => n590);
   U541 : AOI22_X1 port map( A1 => bht_9_4_port, A2 => n1028, B1 => 
                           bht_8_4_port, B2 => n1026, ZN => n570);
   U542 : AOI22_X1 port map( A1 => bht_9_13_port, A2 => n1028, B1 => 
                           bht_8_13_port, B2 => n1026, ZN => n652);
   U543 : AOI22_X1 port map( A1 => bht_9_14_port, A2 => n1028, B1 => 
                           bht_8_14_port, B2 => n1024, ZN => n712);
   U544 : AOI22_X1 port map( A1 => bht_9_12_port, A2 => n1028, B1 => 
                           bht_8_12_port, B2 => n1026, ZN => n672);
   U545 : AOI22_X1 port map( A1 => bht_9_5_port, A2 => n1028, B1 => 
                           bht_8_5_port, B2 => n1024, ZN => n732);
   U546 : AOI22_X1 port map( A1 => bht_23_26_port, A2 => n1112, B1 => 
                           bht_22_26_port, B2 => n990, ZN => n812);
   U547 : NAND4_X1 port map( A1 => n111, A2 => n112, A3 => n113, A4 => n114, ZN
                           => n110);
   U548 : NOR4_X1 port map( A1 => ld_a(12), A2 => ld_a(11), A3 => ld_a(10), A4 
                           => ld_a(0), ZN => n111);
   U549 : NOR4_X1 port map( A1 => ld_a(16), A2 => ld_a(15), A3 => ld_a(14), A4 
                           => ld_a(13), ZN => n112);
   U550 : NOR4_X1 port map( A1 => ld_a(1), A2 => ld_a(19), A3 => ld_a(18), A4 
                           => ld_a(17), ZN => n113);
   U551 : NAND4_X1 port map( A1 => n115, A2 => n116, A3 => n117, A4 => n118, ZN
                           => n109);
   U552 : NOR4_X1 port map( A1 => ld_a(27), A2 => ld_a(26), A3 => ld_a(25), A4 
                           => ld_a(24), ZN => n115);
   U553 : NOR4_X1 port map( A1 => ld_a(30), A2 => ld_a(2), A3 => ld_a(29), A4 
                           => ld_a(28), ZN => n116);
   U554 : NOR4_X1 port map( A1 => ld_a(5), A2 => ld_a(4), A3 => ld_a(3), A4 => 
                           ld_a(31), ZN => n117);
   U555 : AOI22_X1 port map( A1 => bht_15_23_port, A2 => n1047, B1 => 
                           bht_14_23_port, B2 => n1044, ZN => n796);
   U556 : AOI22_X1 port map( A1 => bht_7_9_port, A2 => n1070, B1 => 
                           bht_6_9_port, B2 => n1066, ZN => n743);
   U557 : AOI22_X1 port map( A1 => bht_7_8_port, A2 => n1070, B1 => 
                           bht_6_8_port, B2 => n1067, ZN => n631);
   U558 : AOI22_X1 port map( A1 => bht_7_10_port, A2 => n1070, B1 => 
                           bht_6_10_port, B2 => n1068, ZN => n691);
   U559 : AOI22_X1 port map( A1 => bht_7_6_port, A2 => n1070, B1 => 
                           bht_6_6_port, B2 => n1067, ZN => n589);
   U560 : AOI22_X1 port map( A1 => bht_7_4_port, A2 => n1070, B1 => 
                           bht_6_4_port, B2 => n1068, ZN => n569);
   U561 : AOI22_X1 port map( A1 => bht_7_13_port, A2 => n1070, B1 => 
                           bht_6_13_port, B2 => n1067, ZN => n651);
   U562 : AOI22_X1 port map( A1 => bht_13_23_port, A2 => n1039, B1 => 
                           bht_12_23_port, B2 => n876, ZN => n795);
   U563 : AOI22_X1 port map( A1 => bht_11_23_port, A2 => n1035, B1 => 
                           bht_10_23_port, B2 => n1030, ZN => n794);
   U564 : AOI22_X1 port map( A1 => bht_27_26_port, A2 => n1083, B1 => 
                           bht_26_26_port, B2 => n1078, ZN => n814);
   U565 : AOI22_X1 port map( A1 => bht_1_8_port, A2 => n1052, B1 => 
                           bht_0_8_port, B2 => n1049, ZN => n628);
   U566 : AOI22_X1 port map( A1 => bht_1_4_port, A2 => n1052, B1 => 
                           bht_0_4_port, B2 => n1049, ZN => n566);
   U567 : AOI22_X1 port map( A1 => bht_1_13_port, A2 => n1052, B1 => 
                           bht_0_13_port, B2 => n1050, ZN => n648);
   U568 : AOI22_X1 port map( A1 => bht_25_21_port, A2 => n1075, B1 => 
                           bht_24_21_port, B2 => n1074, ZN => n444);
   U569 : AOI22_X1 port map( A1 => bht_25_20_port, A2 => n1075, B1 => 
                           bht_24_20_port, B2 => n1074, ZN => n464);
   U570 : AOI22_X1 port map( A1 => bht_1_21_port, A2 => n1051, B1 => 
                           bht_0_21_port, B2 => n1049, ZN => n432);
   U571 : AOI22_X1 port map( A1 => bht_9_23_port, A2 => n1029, B1 => 
                           bht_8_23_port, B2 => n1025, ZN => n793);
   U572 : AOI22_X1 port map( A1 => bht_25_19_port, A2 => n1075, B1 => 
                           bht_24_19_port, B2 => n1074, ZN => n484);
   U573 : AOI22_X1 port map( A1 => bht_1_19_port, A2 => n1051, B1 => 
                           bht_0_19_port, B2 => n1048, ZN => n472);
   U574 : AOI22_X1 port map( A1 => bht_1_16_port, A2 => n1051, B1 => 
                           bht_0_16_port, B2 => n1050, ZN => n372);
   U575 : AOI22_X1 port map( A1 => bht_1_15_port, A2 => n1051, B1 => 
                           bht_0_15_port, B2 => n1049, ZN => n392);
   U576 : AOI22_X1 port map( A1 => bht_9_10_port, A2 => n1028, B1 => 
                           bht_8_10_port, B2 => n1024, ZN => n692);
   U577 : AOI22_X1 port map( A1 => bht_1_25_port, A2 => n1051, B1 => 
                           bht_0_25_port, B2 => n1049, ZN => n502);
   U578 : AOI22_X1 port map( A1 => bht_9_9_port, A2 => n1028, B1 => 
                           bht_8_9_port, B2 => n1025, ZN => n744);
   U579 : NAND4_X1 port map( A1 => n194, A2 => n195, A3 => n196, A4 => n197, ZN
                           => n193);
   U580 : NAND4_X1 port map( A1 => n209, A2 => n210, A3 => n211, A4 => n212, ZN
                           => n192);
   U581 : AOI22_X1 port map( A1 => bht_7_23_port, A2 => n1071, B1 => 
                           bht_6_23_port, B2 => n1066, ZN => n792);
   U582 : AOI22_X1 port map( A1 => bht_5_23_port, A2 => n1063, B1 => 
                           bht_4_23_port, B2 => n1061, ZN => n791);
   U583 : AOI22_X1 port map( A1 => bht_3_23_port, A2 => n1059, B1 => 
                           bht_2_23_port, B2 => n1054, ZN => n790);
   U584 : AOI22_X1 port map( A1 => bht_1_22_port, A2 => n1051, B1 => 
                           bht_0_22_port, B2 => n1048, ZN => n412);
   U585 : AOI22_X1 port map( A1 => bht_9_7_port, A2 => n1028, B1 => 
                           bht_8_7_port, B2 => n1024, ZN => n612);
   U586 : AOI22_X1 port map( A1 => bht_1_11_port, A2 => n1051, B1 => 
                           bht_0_11_port, B2 => n1049, ZN => n319);
   U587 : AOI22_X1 port map( A1 => bht_1_23_port, A2 => n1053, B1 => 
                           bht_0_23_port, B2 => n1049, ZN => n789);
   U588 : NAND4_X1 port map( A1 => n223, A2 => n224, A3 => n225, A4 => n226, ZN
                           => n191);
   U589 : AOI22_X1 port map( A1 => bht_1_1_port, A2 => n1051, B1 => 
                           bht_0_1_port, B2 => n1050, ZN => n223);
   U590 : NAND4_X1 port map( A1 => n644, A2 => n645, A3 => n646, A4 => n647, ZN
                           => n638);
   U591 : NAND4_X1 port map( A1 => n700, A2 => n701, A3 => n702, A4 => n703, ZN
                           => n699);
   U592 : NAND4_X1 port map( A1 => n660, A2 => n661, A3 => n662, A4 => n663, ZN
                           => n659);
   U593 : XNOR2_X1 port map( A => n219, B => n799, ZN => n107);
   U594 : AND2_X1 port map( A1 => n951, A2 => n952, ZN => n686);
   U595 : NAND2_X1 port map( A1 => bht_29_10_port, A2 => n868, ZN => n951);
   U596 : NAND2_X1 port map( A1 => bht_28_10_port, A2 => n1086, ZN => n952);
   U597 : AOI22_X1 port map( A1 => bht_1_26_port, A2 => n1053, B1 => 
                           bht_0_26_port, B2 => n1049, ZN => n801);
   U598 : AOI22_X1 port map( A1 => bht_3_26_port, A2 => n1059, B1 => 
                           bht_2_26_port, B2 => n1055, ZN => n802);
   U599 : AOI22_X1 port map( A1 => bht_7_26_port, A2 => n1071, B1 => 
                           bht_6_26_port, B2 => n1067, ZN => n804);
   U600 : NOR4_X1 port map( A1 => n295, A2 => n296, A3 => reg_a(29), A4 => 
                           reg_a(28), ZN => n286);
   U601 : AND4_X1 port map( A1 => n600, A2 => n601, A3 => n602, A4 => n603, ZN 
                           => n970);
   U602 : AND4_X1 port map( A1 => n452, A2 => n453, A3 => n454, A4 => n455, ZN 
                           => n974);
   U603 : AOI22_X1 port map( A1 => bht_1_20_port, A2 => n1051, B1 => 
                           bht_0_20_port, B2 => n1049, ZN => n452);
   U604 : AND4_X1 port map( A1 => n315, A2 => n316, A3 => n317, A4 => n318, ZN 
                           => n985);
   U605 : AND4_X1 port map( A1 => n444, A2 => n445, A3 => n446, A4 => n447, ZN 
                           => n975);
   U606 : AND4_X1 port map( A1 => n297, A2 => n267, A3 => n266, A4 => n265, ZN 
                           => n285);
   U607 : INV_X1 port map( A => reg_a(0), ZN => n297);
   U608 : INV_X1 port map( A => rst, ZN => n1308);
   U609 : OAI22_X1 port map( A1 => n103, A2 => n94, B1 => n100, B2 => n104, ZN 
                           => N3733);
   U610 : NAND2_X1 port map( A1 => sig_brt_delay, A2 => rst, ZN => n104);
   U611 : AOI22_X1 port map( A1 => n120, A2 => n799, B1 => n854, B2 => n860, ZN
                           => n103);
   U612 : NAND2_X1 port map( A1 => net108065, A2 => net108066, ZN => n120);
   U613 : INV_X1 port map( A => addr(27), ZN => n146_port);
   U614 : OAI22_X1 port map( A1 => n955, A2 => n186, B1 => n188_port, B2 => 
                           n953, ZN => N127);
   U615 : INV_X1 port map( A => addr(7), ZN => n186);
   U616 : OAI22_X1 port map( A1 => n955, A2 => n184, B1 => n185, B2 => n953, ZN
                           => N128);
   U617 : INV_X1 port map( A => addr(8), ZN => n184);
   U618 : AOI22_X1 port map( A1 => bht_7_0_port, A2 => n1071, B1 => 
                           bht_6_0_port, B2 => n1067, ZN => n842);
   U619 : AOI22_X1 port map( A1 => bht_15_0_port, A2 => n1047, B1 => 
                           bht_14_0_port, B2 => n1044, ZN => n848);
   U620 : AOI22_X1 port map( A1 => bht_5_0_port, A2 => n1064, B1 => 
                           bht_4_0_port, B2 => n1061, ZN => n841);
   U621 : AOI22_X1 port map( A1 => bht_13_0_port, A2 => n1039, B1 => 
                           bht_12_0_port, B2 => n1038, ZN => n847);
   U622 : AOI22_X1 port map( A1 => bht_3_0_port, A2 => n1059, B1 => 
                           bht_2_0_port, B2 => n1055, ZN => n840);
   U623 : AOI22_X1 port map( A1 => bht_11_0_port, A2 => n1035, B1 => 
                           bht_10_0_port, B2 => n1031, ZN => n846);
   U624 : AOI22_X1 port map( A1 => bht_1_0_port, A2 => n1053, B1 => 
                           bht_0_0_port, B2 => n1049, ZN => n839);
   U625 : AOI22_X1 port map( A1 => bht_9_0_port, A2 => n1029, B1 => 
                           bht_8_0_port, B2 => n1024, ZN => n845);
   U626 : NOR2_X1 port map( A1 => n1306, A2 => n10, ZN => N3737);
   U627 : NOR2_X1 port map( A1 => n1305, A2 => n11, ZN => N3739);
   U628 : NOR2_X1 port map( A1 => n1305, A2 => n12, ZN => N3741);
   U629 : NOR2_X1 port map( A1 => n1305, A2 => n13, ZN => N3743);
   U630 : NOR2_X1 port map( A1 => n1305, A2 => n14, ZN => N3745);
   U631 : NOR2_X1 port map( A1 => n1304, A2 => n15, ZN => N3747);
   U632 : NOR2_X1 port map( A1 => n1304, A2 => n16, ZN => N3749);
   U633 : NOR2_X1 port map( A1 => n1304, A2 => n17, ZN => N3751);
   U634 : NOR2_X1 port map( A1 => n1304, A2 => n18, ZN => N3753);
   U635 : NOR2_X1 port map( A1 => n1303, A2 => n19, ZN => N3755);
   U636 : NOR2_X1 port map( A1 => n1303, A2 => n20, ZN => N3757);
   U637 : NOR2_X1 port map( A1 => n1303, A2 => n21, ZN => N3759);
   U638 : NOR2_X1 port map( A1 => n1303, A2 => n22, ZN => N3761);
   U639 : NOR2_X1 port map( A1 => n1302, A2 => n23, ZN => N3763);
   U640 : NOR2_X1 port map( A1 => n1302, A2 => n24, ZN => N3765);
   U641 : NOR2_X1 port map( A1 => n1302, A2 => n25, ZN => N3767);
   U642 : NOR2_X1 port map( A1 => n1302, A2 => n26, ZN => N3769);
   U643 : NOR2_X1 port map( A1 => n1301, A2 => n27, ZN => N3771);
   U644 : NOR2_X1 port map( A1 => n1301, A2 => n28, ZN => N3773);
   U645 : NOR2_X1 port map( A1 => n1301, A2 => n29, ZN => N3775);
   U646 : NOR2_X1 port map( A1 => n1301, A2 => n30, ZN => N3777);
   U647 : NOR2_X1 port map( A1 => n1300, A2 => n31, ZN => N3779);
   U648 : NOR2_X1 port map( A1 => n1300, A2 => n32, ZN => N3781);
   U649 : NOR2_X1 port map( A1 => n1300, A2 => n33, ZN => N3785);
   U650 : NOR2_X1 port map( A1 => n1300, A2 => n9, ZN => N3783);
   U651 : NAND4_X1 port map( A1 => n821, A2 => n822, A3 => n823, A4 => n824, ZN
                           => n820);
   U652 : AOI22_X1 port map( A1 => bht_21_0_port, A2 => n1107, B1 => 
                           bht_20_0_port, B2 => n865, ZN => n823);
   U653 : AOI22_X1 port map( A1 => bht_23_0_port, A2 => n1111, B1 => 
                           bht_22_0_port, B2 => n990, ZN => n824);
   U654 : NAND4_X1 port map( A1 => n833, A2 => n834, A3 => n835, A4 => n836, ZN
                           => n819);
   U655 : AOI22_X1 port map( A1 => bht_25_0_port, A2 => n1077, B1 => 
                           bht_24_0_port, B2 => n1072, ZN => n833);
   U656 : AOI22_X1 port map( A1 => bht_27_0_port, A2 => n1083, B1 => 
                           bht_26_0_port, B2 => n1080, ZN => n834);
   U657 : BUF_X1 port map( A => sig_bal, Z => n1295);
   U658 : BUF_X1 port map( A => sig_bal, Z => n1296);
   U659 : OR4_X1 port map( A1 => reg_a(25), A2 => reg_a(1), A3 => reg_a(27), A4
                           => reg_a(26), ZN => n295);
   U660 : BUF_X1 port map( A => sig_bal, Z => n1294);
   U661 : BUF_X1 port map( A => sig_bal, Z => n1297);
   U662 : BUF_X1 port map( A => sig_bal, Z => n1299);
   U663 : BUF_X1 port map( A => sig_bal, Z => n1298);
   U664 : OR3_X1 port map( A1 => n1294, A2 => reg_a(31), A3 => reg_a(30), ZN =>
                           n296);
   U665 : INV_X1 port map( A => n182, ZN => N129);
   U666 : INV_X1 port map( A => n180, ZN => N130);
   U667 : INV_X1 port map( A => n178, ZN => N131);
   U668 : INV_X1 port map( A => n176, ZN => N132);
   U669 : INV_X1 port map( A => n174, ZN => N133);
   U670 : INV_X1 port map( A => n172, ZN => N134);
   U671 : INV_X1 port map( A => n170, ZN => N135);
   U672 : INV_X1 port map( A => n168, ZN => N136);
   U673 : INV_X1 port map( A => n166, ZN => N137);
   U674 : INV_X1 port map( A => n164, ZN => N138);
   U675 : INV_X1 port map( A => n162, ZN => N139);
   U676 : INV_X1 port map( A => n158, ZN => N141);
   U677 : INV_X1 port map( A => n137_port, ZN => N151);
   U678 : INV_X1 port map( A => n156, ZN => N142);
   U679 : AOI22_X1 port map( A1 => n953, A2 => addr(22), B1 => n157, B2 => n955
                           , ZN => n156);
   U680 : INV_X1 port map( A => n140_port, ZN => N150);
   U681 : INV_X1 port map( A => n160, ZN => N140);
   U682 : INV_X1 port map( A => n154, ZN => N143);
   U683 : INV_X1 port map( A => n152, ZN => N144);
   U684 : INV_X1 port map( A => n150_port, ZN => N145);
   U685 : INV_X1 port map( A => n148_port, ZN => N146);
   U686 : INV_X1 port map( A => n144_port, ZN => N148);
   U687 : INV_X1 port map( A => n142_port, ZN => N149);
   U688 : AOI22_X1 port map( A1 => bht_19_0_port, A2 => n1102, B1 => 
                           bht_18_0_port, B2 => n872, ZN => n822);
   U689 : AND4_X1 port map( A1 => n789, A2 => n790, A3 => n791, A4 => n792, ZN 
                           => n995);
   U690 : AND4_X1 port map( A1 => n785, A2 => n786, A3 => n787, A4 => n788, ZN 
                           => n996);
   U691 : AND2_X1 port map( A1 => n825, A2 => n826, ZN => n990);
   U692 : CLKBUF_X1 port map( A => n208, Z => n963);
   U693 : INV_X1 port map( A => n956, ZN => n953);
   U694 : INV_X1 port map( A => n956, ZN => n954);
   U695 : NAND2_X1 port map( A1 => n1020, A2 => n964, ZN => n1013);
   U696 : NOR2_X1 port map( A1 => opcd(1), A2 => n1010, ZN => n964);
   U697 : AOI22_X1 port map( A1 => bht_11_1_port, A2 => n1033, B1 => 
                           bht_10_1_port, B2 => n1032, ZN => n236);
   U698 : AOI22_X1 port map( A1 => bht_11_11_port, A2 => n1033, B1 => 
                           bht_10_11_port, B2 => n1032, ZN => n324);
   U699 : AOI22_X1 port map( A1 => bht_11_22_port, A2 => n1033, B1 => 
                           bht_10_22_port, B2 => n1031, ZN => n417);
   U700 : AOI22_X1 port map( A1 => bht_11_25_port, A2 => n1033, B1 => 
                           bht_10_25_port, B2 => n1031, ZN => n507);
   U701 : AOI22_X1 port map( A1 => bht_11_3_port, A2 => n1033, B1 => 
                           bht_10_3_port, B2 => n1031, ZN => n522);
   U702 : AOI22_X1 port map( A1 => bht_11_16_port, A2 => n1033, B1 => 
                           bht_10_16_port, B2 => n1030, ZN => n377);
   U703 : AOI22_X1 port map( A1 => bht_11_19_port, A2 => n1033, B1 => 
                           bht_10_19_port, B2 => n1030, ZN => n477);
   U704 : AOI22_X1 port map( A1 => bht_11_17_port, A2 => n1033, B1 => 
                           bht_10_17_port, B2 => n1032, ZN => n356);
   U705 : AOI22_X1 port map( A1 => bht_11_18_port, A2 => n1033, B1 => 
                           bht_10_18_port, B2 => n1030, ZN => n336);
   U706 : NAND4_X1 port map( A1 => n704, A2 => n705, A3 => n706, A4 => n707, ZN
                           => n698);
   U707 : AND2_X1 port map( A1 => n828, A2 => n838, ZN => n216);
   U708 : AOI22_X1 port map( A1 => bht_17_26_port, A2 => n1097, B1 => n863, B2 
                           => bht_16_26_port, ZN => n809);
   U709 : AOI22_X1 port map( A1 => bht_17_0_port, A2 => n1098, B1 => 
                           bht_16_0_port, B2 => n869, ZN => n821);
   U710 : INV_X1 port map( A => addr(5), ZN => n966);
   U711 : NAND4_X1 port map( A1 => n967, A2 => n968, A3 => n969, A4 => n970, ZN
                           => n177);
   U712 : AND4_X1 port map( A1 => n612, A2 => n613, A3 => n614, A4 => n615, ZN 
                           => n967);
   U713 : AND4_X1 port map( A1 => n608, A2 => n609, A3 => n610, A4 => n611, ZN 
                           => n968);
   U714 : AND2_X1 port map( A1 => n837, A2 => n826, ZN => n215);
   U715 : NAND4_X1 port map( A1 => n971, A2 => n972, A3 => n973, A4 => n974, ZN
                           => n151_port);
   U716 : AND4_X1 port map( A1 => n460, A2 => n461, A3 => n462, A4 => n463, ZN 
                           => n972);
   U717 : AND4_X1 port map( A1 => n456, A2 => n457, A3 => n458, A4 => n459, ZN 
                           => n973);
   U718 : AOI22_X1 port map( A1 => bht_11_5_port, A2 => n1034, B1 => 
                           bht_10_5_port, B2 => n1031, ZN => n733);
   U719 : AOI22_X1 port map( A1 => bht_11_12_port, A2 => n1034, B1 => 
                           bht_10_12_port, B2 => n1031, ZN => n673);
   U720 : AOI22_X1 port map( A1 => bht_11_13_port, A2 => n1034, B1 => 
                           bht_10_13_port, B2 => n1031, ZN => n653);
   U721 : AOI22_X1 port map( A1 => bht_11_14_port, A2 => n1034, B1 => 
                           bht_10_14_port, B2 => n1031, ZN => n713);
   U722 : AOI22_X1 port map( A1 => bht_11_4_port, A2 => n1034, B1 => 
                           bht_10_4_port, B2 => n1031, ZN => n571);
   U723 : AOI22_X1 port map( A1 => bht_11_6_port, A2 => n1034, B1 => 
                           bht_10_6_port, B2 => n1032, ZN => n591);
   U724 : AOI22_X1 port map( A1 => bht_11_7_port, A2 => n1034, B1 => 
                           bht_10_7_port, B2 => n1032, ZN => n613);
   U725 : AOI22_X1 port map( A1 => bht_11_8_port, A2 => n1034, B1 => 
                           bht_10_8_port, B2 => n1031, ZN => n633);
   U726 : AOI22_X1 port map( A1 => bht_11_9_port, A2 => n1034, B1 => 
                           bht_10_9_port, B2 => n1030, ZN => n745);
   U727 : AOI22_X1 port map( A1 => bht_11_2_port, A2 => n1034, B1 => 
                           bht_10_2_port, B2 => n1031, ZN => n542);
   U728 : AOI22_X1 port map( A1 => bht_11_10_port, A2 => n1034, B1 => 
                           bht_10_10_port, B2 => n1031, ZN => n693);
   U729 : AOI22_X1 port map( A1 => bht_11_24_port, A2 => n1034, B1 => 
                           bht_10_24_port, B2 => n1030, ZN => n774);
   U730 : BUF_X1 port map( A => n215, Z => n1092);
   U731 : AOI22_X1 port map( A1 => bht_9_1_port, A2 => n1027, B1 => 
                           bht_8_1_port, B2 => n1026, ZN => n235);
   U732 : AOI22_X1 port map( A1 => bht_9_11_port, A2 => n1027, B1 => 
                           bht_8_11_port, B2 => n1024, ZN => n323);
   U733 : AOI22_X1 port map( A1 => bht_9_21_port, A2 => n1027, B1 => 
                           bht_8_21_port, B2 => n1024, ZN => n436);
   U734 : AOI22_X1 port map( A1 => bht_9_22_port, A2 => n1027, B1 => 
                           bht_8_22_port, B2 => n1025, ZN => n416);
   U735 : AOI22_X1 port map( A1 => bht_9_25_port, A2 => n1027, B1 => 
                           bht_8_25_port, B2 => n1024, ZN => n506);
   U736 : AOI22_X1 port map( A1 => bht_9_3_port, A2 => n1027, B1 => 
                           bht_8_3_port, B2 => n1026, ZN => n521);
   U737 : AOI22_X1 port map( A1 => bht_9_16_port, A2 => n1027, B1 => 
                           bht_8_16_port, B2 => n1026, ZN => n376);
   U738 : AOI22_X1 port map( A1 => bht_9_17_port, A2 => n1027, B1 => 
                           bht_8_17_port, B2 => n1026, ZN => n355);
   U739 : AOI22_X1 port map( A1 => bht_9_19_port, A2 => n1027, B1 => 
                           bht_8_19_port, B2 => n1026, ZN => n476);
   U740 : AOI22_X1 port map( A1 => bht_9_18_port, A2 => n1027, B1 => 
                           bht_8_18_port, B2 => n1025, ZN => n335);
   U741 : AOI22_X1 port map( A1 => bht_9_20_port, A2 => n1027, B1 => 
                           bht_8_20_port, B2 => n1026, ZN => n456);
   U742 : AOI22_X1 port map( A1 => bht_9_24_port, A2 => n1028, B1 => 
                           bht_8_24_port, B2 => n1025, ZN => n773);
   U743 : BUF_X1 port map( A => n222, Z => n1073);
   U744 : AOI22_X1 port map( A1 => bht_7_7_port, A2 => n1070, B1 => 
                           bht_6_7_port, B2 => n1067, ZN => n611);
   U745 : AOI22_X1 port map( A1 => bht_29_1_port, A2 => n867, B1 => 
                           bht_28_1_port, B2 => n1086, ZN => n211);
   U746 : NAND4_X1 port map( A1 => n484, A2 => n485, A3 => n486, A4 => n487, ZN
                           => n468);
   U747 : AND2_X1 port map( A1 => addr(3), A2 => addr(4), ZN => n826);
   U748 : AOI22_X1 port map( A1 => bht_11_15_port, A2 => n1033, B1 => 
                           bht_10_15_port, B2 => n1031, ZN => n397);
   U749 : AOI22_X1 port map( A1 => bht_9_15_port, A2 => n1027, B1 => 
                           bht_8_15_port, B2 => n1024, ZN => n396);
   U750 : AOI22_X1 port map( A1 => bht_15_5_port, A2 => n1046, B1 => 
                           bht_14_5_port, B2 => n1043, ZN => n735);
   U751 : AOI22_X1 port map( A1 => bht_15_12_port, A2 => n1046, B1 => 
                           bht_14_12_port, B2 => n1043, ZN => n675);
   U752 : AOI22_X1 port map( A1 => bht_15_13_port, A2 => n1046, B1 => 
                           bht_14_13_port, B2 => n1043, ZN => n655);
   U753 : AND4_X1 port map( A1 => n773, A2 => n774, A3 => n775, A4 => n776, ZN 
                           => n1004);
   U754 : AOI22_X1 port map( A1 => bht_15_14_port, A2 => n1046, B1 => 
                           bht_14_14_port, B2 => n1043, ZN => n715);
   U755 : AOI22_X1 port map( A1 => bht_15_4_port, A2 => n1046, B1 => 
                           bht_14_4_port, B2 => n1043, ZN => n573);
   U756 : AOI22_X1 port map( A1 => bht_15_6_port, A2 => n1046, B1 => 
                           bht_14_6_port, B2 => n1043, ZN => n593);
   U757 : AOI22_X1 port map( A1 => bht_15_8_port, A2 => n1046, B1 => 
                           bht_14_8_port, B2 => n1043, ZN => n635);
   U758 : AOI22_X1 port map( A1 => bht_15_7_port, A2 => n1046, B1 => 
                           bht_14_7_port, B2 => n1043, ZN => n615);
   U759 : AOI22_X1 port map( A1 => bht_15_9_port, A2 => n1046, B1 => 
                           bht_14_9_port, B2 => n1043, ZN => n747);
   U760 : AOI22_X1 port map( A1 => bht_15_2_port, A2 => n1046, B1 => 
                           bht_14_2_port, B2 => n1043, ZN => n544);
   U761 : AOI22_X1 port map( A1 => bht_15_10_port, A2 => n1046, B1 => 
                           bht_14_10_port, B2 => n1043, ZN => n695);
   U762 : AOI22_X1 port map( A1 => bht_15_24_port, A2 => n1046, B1 => 
                           bht_14_24_port, B2 => n1043, ZN => n776);
   U763 : AND2_X1 port map( A1 => n827, A2 => n830, ZN => n206);
   U764 : BUF_X1 port map( A => n204, Z => n1104);
   U765 : AOI22_X1 port map( A1 => bht_21_26_port, A2 => n1107, B1 => 
                           bht_20_26_port, B2 => n1015, ZN => n811);
   U766 : AOI22_X1 port map( A1 => bht_1_24_port, A2 => n1052, B1 => 
                           bht_0_24_port, B2 => n1048, ZN => n769);
   U767 : AOI22_X1 port map( A1 => bht_1_7_port, A2 => n1052, B1 => 
                           bht_0_7_port, B2 => n1050, ZN => n608);
   U768 : AOI22_X1 port map( A1 => bht_1_2_port, A2 => n1052, B1 => 
                           bht_0_2_port, B2 => n1050, ZN => n537);
   U769 : AOI22_X1 port map( A1 => bht_1_9_port, A2 => n1052, B1 => 
                           bht_0_9_port, B2 => n1048, ZN => n740);
   U770 : AOI22_X1 port map( A1 => bht_1_10_port, A2 => n1052, B1 => 
                           bht_0_10_port, B2 => n1049, ZN => n688);
   U771 : AOI22_X1 port map( A1 => bht_1_6_port, A2 => n1052, B1 => 
                           bht_0_6_port, B2 => n1049, ZN => n586);
   U772 : OAI222_X1 port map( A1 => n256, A2 => n163, B1 => n257, B2 => n177, 
                           C1 => n258, C2 => n175, ZN => n255);
   U773 : AOI22_X1 port map( A1 => bht_11_20_port, A2 => n1033, B1 => 
                           bht_10_20_port, B2 => n1032, ZN => n457);
   U774 : BUF_X1 port map( A => n220, Z => n1078);
   U775 : AOI22_X1 port map( A1 => n953, A2 => addr(21), B1 => n159, B2 => n956
                           , ZN => n158);
   U776 : AOI22_X1 port map( A1 => bht_19_26_port, A2 => n874, B1 => 
                           bht_18_26_port, B2 => n1099, ZN => n810);
   U777 : BUF_X1 port map( A => n203, Z => n1106);
   U778 : NAND4_X1 port map( A1 => n482, A2 => n480, A3 => n483, A4 => n481, ZN
                           => n469);
   U779 : AOI22_X1 port map( A1 => n954, A2 => addr(20), B1 => n161, B2 => n960
                           , ZN => n160);
   U780 : AOI22_X1 port map( A1 => bht_15_1_port, A2 => n1045, B1 => 
                           bht_14_1_port, B2 => n1042, ZN => n238);
   U781 : AOI22_X1 port map( A1 => bht_15_11_port, A2 => n1045, B1 => 
                           bht_14_11_port, B2 => n1042, ZN => n326);
   U782 : AOI22_X1 port map( A1 => bht_15_25_port, A2 => n1045, B1 => 
                           bht_14_25_port, B2 => n1042, ZN => n509);
   U783 : AOI22_X1 port map( A1 => bht_15_3_port, A2 => n1045, B1 => 
                           bht_14_3_port, B2 => n1042, ZN => n524);
   U784 : AOI22_X1 port map( A1 => bht_15_17_port, A2 => n1045, B1 => 
                           bht_14_17_port, B2 => n1042, ZN => n358);
   U785 : AOI22_X1 port map( A1 => bht_15_15_port, A2 => n1045, B1 => 
                           bht_14_15_port, B2 => n1042, ZN => n399);
   U786 : NAND4_X1 port map( A1 => n975, A2 => n976, A3 => n977, A4 => n978, ZN
                           => n149_port);
   U787 : AND4_X1 port map( A1 => n440, A2 => n441, A3 => n442, A4 => n443, ZN 
                           => n976);
   U788 : AOI22_X1 port map( A1 => bht_3_1_port, A2 => n1057, B1 => 
                           bht_2_1_port, B2 => n1056, ZN => n224);
   U789 : OAI222_X1 port map( A1 => n259, A2 => n169, B1 => n260, B2 => n167, 
                           C1 => n261, C2 => n165, ZN => n254);
   U790 : AOI22_X1 port map( A1 => bht_3_11_port, A2 => n1057, B1 => 
                           bht_2_11_port, B2 => n1056, ZN => n320);
   U791 : AOI22_X1 port map( A1 => bht_3_22_port, A2 => n1057, B1 => 
                           bht_2_22_port, B2 => n1054, ZN => n413);
   U792 : AOI22_X1 port map( A1 => bht_3_25_port, A2 => n1057, B1 => 
                           bht_2_25_port, B2 => n1055, ZN => n503);
   U793 : AOI22_X1 port map( A1 => bht_3_3_port, A2 => n1057, B1 => 
                           bht_2_3_port, B2 => n1055, ZN => n518);
   U794 : AOI22_X1 port map( A1 => bht_3_16_port, A2 => n1057, B1 => 
                           bht_2_16_port, B2 => n1055, ZN => n373);
   U795 : AOI22_X1 port map( A1 => bht_3_17_port, A2 => n1057, B1 => 
                           bht_2_17_port, B2 => n1055, ZN => n352);
   U796 : AOI22_X1 port map( A1 => bht_3_20_port, A2 => n1057, B1 => 
                           bht_2_20_port, B2 => n1056, ZN => n453);
   U797 : AOI22_X1 port map( A1 => n954, A2 => addr(30), B1 => n141_port, B2 =>
                           n960, ZN => n140_port);
   U798 : NAND4_X1 port map( A1 => n628, A2 => n629, A3 => n630, A4 => n631, ZN
                           => n617);
   U799 : NAND4_X1 port map( A1 => n624, A2 => n625, A3 => n626, A4 => n627, ZN
                           => n618);
   U800 : AOI22_X1 port map( A1 => bht_7_24_port, A2 => n1070, B1 => 
                           bht_6_24_port, B2 => n1066, ZN => n772);
   U801 : NAND4_X1 port map( A1 => n474, A2 => n472, A3 => n473, A4 => n475, ZN
                           => n471);
   U802 : AOI22_X1 port map( A1 => bht_3_19_port, A2 => n1057, B1 => 
                           bht_2_19_port, B2 => n1054, ZN => n473);
   U803 : NAND4_X1 port map( A1 => n476, A2 => n479, A3 => n477, A4 => n478, ZN
                           => n470);
   U804 : NAND4_X1 port map( A1 => n648, A2 => n649, A3 => n650, A4 => n651, ZN
                           => n637);
   U805 : AOI22_X1 port map( A1 => bht_3_12_port, A2 => n1058, B1 => 
                           bht_2_12_port, B2 => n1056, ZN => n669);
   U806 : AOI22_X1 port map( A1 => bht_3_5_port, A2 => n1058, B1 => 
                           bht_2_5_port, B2 => n1055, ZN => n729);
   U807 : AOI22_X1 port map( A1 => bht_3_13_port, A2 => n1058, B1 => 
                           bht_2_13_port, B2 => n1055, ZN => n649);
   U808 : AOI22_X1 port map( A1 => bht_3_14_port, A2 => n1058, B1 => 
                           bht_2_14_port, B2 => n1055, ZN => n709);
   U809 : AOI22_X1 port map( A1 => bht_3_6_port, A2 => n1058, B1 => 
                           bht_2_6_port, B2 => n1055, ZN => n587);
   U810 : AOI22_X1 port map( A1 => bht_3_4_port, A2 => n1058, B1 => 
                           bht_2_4_port, B2 => n1056, ZN => n567);
   U811 : AOI22_X1 port map( A1 => bht_3_9_port, A2 => n1058, B1 => 
                           bht_2_9_port, B2 => n1054, ZN => n741);
   U812 : AOI22_X1 port map( A1 => bht_3_10_port, A2 => n1058, B1 => 
                           bht_2_10_port, B2 => n1056, ZN => n689);
   U813 : AOI22_X1 port map( A1 => bht_3_8_port, A2 => n1058, B1 => 
                           bht_2_8_port, B2 => n1055, ZN => n629);
   U814 : AOI22_X1 port map( A1 => bht_3_2_port, A2 => n1058, B1 => 
                           bht_2_2_port, B2 => n1056, ZN => n538);
   U815 : AOI22_X1 port map( A1 => bht_3_7_port, A2 => n1058, B1 => 
                           bht_2_7_port, B2 => n1055, ZN => n609);
   U816 : AOI22_X1 port map( A1 => bht_3_24_port, A2 => n1058, B1 => 
                           bht_2_24_port, B2 => n1054, ZN => n770);
   U817 : AOI22_X1 port map( A1 => n954, A2 => addr(26), B1 => n149_port, B2 =>
                           n960, ZN => n148_port);
   U818 : OAI22_X1 port map( A1 => n271, A2 => n161, B1 => n272, B2 => 
                           n149_port, ZN => n270);
   U819 : AOI22_X1 port map( A1 => bht_3_15_port, A2 => n1057, B1 => 
                           bht_2_15_port, B2 => n1056, ZN => n393);
   U820 : AND4_X1 port map( A1 => n767, A2 => n768, A3 => n766, A4 => n765, ZN 
                           => n1006);
   U821 : NAND4_X1 port map( A1 => n620, A2 => n621, A3 => n622, A4 => n623, ZN
                           => n619);
   U822 : AOI22_X1 port map( A1 => n954, A2 => addr(24), B1 => n889, B2 => n960
                           , ZN => n152);
   U824 : AND4_X1 port map( A1 => n424, A2 => n425, A3 => n426, A4 => n427, ZN 
                           => n979);
   U825 : AND4_X1 port map( A1 => n420, A2 => n421, A3 => n422, A4 => n423, ZN 
                           => n980);
   U826 : AND4_X1 port map( A1 => n416, A2 => n417, A3 => n418, A4 => n419, ZN 
                           => n981);
   U827 : AND4_X1 port map( A1 => n412, A2 => n413, A3 => n414, A4 => n415, ZN 
                           => n982);
   U828 : AND2_X1 port map( A1 => n843, A2 => n826, ZN => n228);
   U829 : AND2_X1 port map( A1 => n829, A2 => n843, ZN => n232);
   U830 : AOI22_X1 port map( A1 => n954, A2 => addr(23), B1 => n155, B2 => n959
                           , ZN => n154);
   U831 : NAND4_X1 port map( A1 => n983, A2 => n984, A3 => n985, A4 => n986, ZN
                           => n169);
   U832 : AND4_X1 port map( A1 => n323, A2 => n324, A3 => n325, A4 => n326, ZN 
                           => n983);
   U833 : AND4_X1 port map( A1 => n319, A2 => n320, A3 => n321, A4 => n322, ZN 
                           => n984);
   U834 : AND4_X1 port map( A1 => n311, A2 => n313, A3 => n312, A4 => n314, ZN 
                           => n986);
   U835 : AOI22_X1 port map( A1 => bht_3_21_port, A2 => n1057, B1 => 
                           bht_2_21_port, B2 => n1055, ZN => n433);
   U836 : AND2_X1 port map( A1 => n844, A2 => n830, ZN => n233);
   U850 : AND2_X1 port map( A1 => n844, A2 => n826, ZN => n227);
   U851 : AND2_X1 port map( A1 => n828, A2 => n844, ZN => n229);
   U852 : CLKBUF_X1 port map( A => addr(5), Z => n987);
   U853 : AND2_X1 port map( A1 => n850, A2 => n826, ZN => n239);
   U854 : AND2_X1 port map( A1 => n830, A2 => n850, ZN => n245);
   U855 : AND2_X1 port map( A1 => n828, A2 => n850, ZN => n241);
   U856 : CLKBUF_X1 port map( A => n169, Z => n988);
   U857 : AOI22_X1 port map( A1 => bht_31_0_port, A2 => n1095, B1 => 
                           bht_30_0_port, B2 => n1091, ZN => n836);
   U858 : AOI22_X1 port map( A1 => bht_31_26_port, A2 => n1095, B1 => 
                           bht_30_26_port, B2 => n1092, ZN => n816);
   U859 : AOI22_X1 port map( A1 => n954, A2 => addr(25), B1 => n887, B2 => n959
                           , ZN => n150_port);
   U860 : INV_X1 port map( A => n281, ZN => n171);
   U861 : AOI22_X1 port map( A1 => n175, A2 => n258, B1 => n177, B2 => n257, ZN
                           => n595);
   U862 : AOI22_X1 port map( A1 => bht_1_18_port, A2 => n1051, B1 => 
                           bht_0_18_port, B2 => n1049, ZN => n331);
   U863 : AOI22_X1 port map( A1 => bht_3_18_port, A2 => n1057, B1 => 
                           bht_2_18_port, B2 => n1054, ZN => n332);
   U864 : AOI22_X1 port map( A1 => bht_7_1_port, A2 => n1069, B1 => 
                           bht_6_1_port, B2 => n1068, ZN => n226);
   U865 : AOI22_X1 port map( A1 => bht_7_16_port, A2 => n1069, B1 => 
                           bht_6_16_port, B2 => n1067, ZN => n375);
   U866 : AOI22_X1 port map( A1 => bht_7_3_port, A2 => n1069, B1 => 
                           bht_6_3_port, B2 => n1068, ZN => n520);
   U867 : AOI22_X1 port map( A1 => bht_7_17_port, A2 => n1069, B1 => 
                           bht_6_17_port, B2 => n1067, ZN => n354);
   U868 : AOI22_X1 port map( A1 => bht_7_25_port, A2 => n1069, B1 => 
                           bht_6_25_port, B2 => n1067, ZN => n505);
   U869 : AOI22_X1 port map( A1 => bht_7_20_port, A2 => n1069, B1 => 
                           bht_6_20_port, B2 => n1068, ZN => n455);
   U870 : AOI22_X1 port map( A1 => bht_7_15_port, A2 => n1069, B1 => 
                           bht_6_15_port, B2 => n1068, ZN => n395);
   U871 : AOI22_X1 port map( A1 => bht_7_21_port, A2 => n1069, B1 => 
                           bht_6_21_port, B2 => n1067, ZN => n435);
   U872 : AOI22_X1 port map( A1 => bht_7_19_port, A2 => n1069, B1 => 
                           bht_6_19_port, B2 => n1066, ZN => n475);
   U873 : AOI22_X1 port map( A1 => bht_7_11_port, A2 => n1069, B1 => 
                           bht_6_11_port, B2 => n1067, ZN => n322);
   U874 : AOI22_X1 port map( A1 => bht_7_22_port, A2 => n1069, B1 => 
                           bht_6_22_port, B2 => n1066, ZN => n415);
   U875 : AOI22_X1 port map( A1 => bht_7_18_port, A2 => n1069, B1 => 
                           bht_6_18_port, B2 => n1067, ZN => n334);
   U876 : AOI22_X1 port map( A1 => bht_29_0_port, A2 => n1087, B1 => 
                           bht_28_0_port, B2 => n1085, ZN => n835);
   U877 : AOI22_X1 port map( A1 => bht_29_3_port, A2 => n1089, B1 => 
                           bht_28_3_port, B2 => n1085, ZN => n531);
   U878 : AOI22_X1 port map( A1 => bht_29_17_port, A2 => n868, B1 => 
                           bht_28_17_port, B2 => n1086, ZN => n365);
   U879 : AOI22_X1 port map( A1 => bht_29_18_port, A2 => n1087, B1 => 
                           bht_28_18_port, B2 => n1086, ZN => n345);
   U880 : AOI22_X1 port map( A1 => bht_25_3_port, A2 => n1075, B1 => 
                           bht_24_3_port, B2 => n1009, ZN => n529);
   U881 : AOI22_X1 port map( A1 => bht_25_17_port, A2 => n1075, B1 => 
                           bht_24_17_port, B2 => n1009, ZN => n363);
   U882 : AOI22_X1 port map( A1 => bht_25_16_port, A2 => n1075, B1 => 
                           bht_24_16_port, B2 => n1009, ZN => n384);
   U883 : AOI22_X1 port map( A1 => bht_25_18_port, A2 => n1075, B1 => 
                           bht_24_18_port, B2 => n1009, ZN => n343);
   U884 : AOI22_X1 port map( A1 => bht_25_11_port, A2 => n1075, B1 => 
                           bht_24_11_port, B2 => n1009, ZN => n315);
   U885 : AND2_X1 port map( A1 => n849, A2 => n826, ZN => n240);
   U886 : AND2_X1 port map( A1 => n849, A2 => n830, ZN => n246);
   U887 : AOI22_X1 port map( A1 => bht_11_21_port, A2 => n1033, B1 => 
                           bht_10_21_port, B2 => n1031, ZN => n437);
   U888 : AOI22_X1 port map( A1 => bht_15_21_port, A2 => n1045, B1 => 
                           bht_14_21_port, B2 => n1042, ZN => n439);
   U889 : AOI22_X1 port map( A1 => bht_15_20_port, A2 => n1045, B1 => 
                           bht_14_20_port, B2 => n1042, ZN => n459);
   U890 : AOI22_X1 port map( A1 => bht_15_18_port, A2 => n1045, B1 => 
                           bht_14_18_port, B2 => n1042, ZN => n338);
   U891 : AOI22_X1 port map( A1 => bht_15_22_port, A2 => n1045, B1 => 
                           bht_14_22_port, B2 => n1042, ZN => n419);
   U892 : AOI22_X1 port map( A1 => bht_15_19_port, A2 => n1045, B1 => 
                           bht_14_19_port, B2 => n1042, ZN => n479);
   U893 : AOI22_X1 port map( A1 => bht_15_16_port, A2 => n1045, B1 => 
                           bht_14_16_port, B2 => n1042, ZN => n379);
   U894 : AND2_X1 port map( A1 => n825, A2 => n826, ZN => n989);
   U895 : AND2_X1 port map( A1 => n825, A2 => n826, ZN => n199);
   U896 : AOI22_X1 port map( A1 => bht_17_1_port, A2 => n1097, B1 => 
                           bht_16_1_port, B2 => n871, ZN => n194);
   U897 : AOI22_X1 port map( A1 => bht_17_3_port, A2 => n1098, B1 => 
                           bht_16_3_port, B2 => n869, ZN => n525);
   U898 : AOI22_X1 port map( A1 => bht_17_17_port, A2 => n1097, B1 => 
                           bht_16_17_port, B2 => n208, ZN => n359);
   U899 : AOI22_X1 port map( A1 => bht_17_15_port, A2 => n1098, B1 => 
                           bht_16_15_port, B2 => n208, ZN => n400);
   U900 : AOI22_X1 port map( A1 => n1096, A2 => bht_17_19_port, B1 => n208, B2 
                           => bht_16_19_port, ZN => n480);
   U901 : AOI22_X1 port map( A1 => bht_17_22_port, A2 => n1098, B1 => 
                           bht_16_22_port, B2 => n208, ZN => n420);
   U902 : AOI22_X1 port map( A1 => bht_17_20_port, A2 => n1097, B1 => 
                           bht_16_20_port, B2 => n871, ZN => n460);
   U903 : AOI22_X1 port map( A1 => bht_25_1_port, A2 => n1075, B1 => 
                           bht_24_1_port, B2 => n1008, ZN => n209);
   U904 : AOI22_X1 port map( A1 => bht_25_26_port, A2 => n1077, B1 => 
                           bht_24_26_port, B2 => n1008, ZN => n813);
   U905 : AOI22_X1 port map( A1 => bht_25_15_port, A2 => n1075, B1 => 
                           bht_24_15_port, B2 => n1008, ZN => n404);
   U906 : AOI22_X1 port map( A1 => bht_25_22_port, A2 => n1075, B1 => 
                           bht_24_22_port, B2 => n1008, ZN => n424);
   U907 : AOI22_X1 port map( A1 => bht_25_25_port, A2 => n1075, B1 => 
                           bht_24_25_port, B2 => n1008, ZN => n498);
   U908 : NAND2_X1 port map( A1 => n898, A2 => n276, ZN => n991);
   U909 : NAND2_X1 port map( A1 => n161, A2 => n271, ZN => n992);
   U910 : NAND2_X1 port map( A1 => n159, A2 => n266, ZN => n993);
   U911 : AND3_X1 port map( A1 => n991, A2 => n992, A3 => n993, ZN => n305);
   U912 : AOI22_X1 port map( A1 => bht_21_1_port, A2 => n1109, B1 => 
                           bht_20_1_port, B2 => n1014, ZN => n196);
   U913 : AOI22_X1 port map( A1 => bht_21_3_port, A2 => n1107, B1 => 
                           bht_20_3_port, B2 => n1106, ZN => n527);
   U914 : AOI22_X1 port map( A1 => bht_21_17_port, A2 => n1107, B1 => 
                           bht_20_17_port, B2 => n861, ZN => n361);
   U915 : AOI22_X1 port map( A1 => bht_21_22_port, A2 => n1108, B1 => 
                           bht_20_22_port, B2 => n1014, ZN => n422);
   U916 : AOI22_X1 port map( A1 => bht_21_19_port, A2 => n1108, B1 => n1105, B2
                           => bht_20_19_port, ZN => n482);
   U917 : AOI22_X1 port map( A1 => bht_21_20_port, A2 => n1107, B1 => 
                           bht_20_20_port, B2 => n1015, ZN => n462);
   U918 : AOI22_X1 port map( A1 => bht_21_21_port, A2 => n1107, B1 => n865, B2 
                           => bht_20_21_port, ZN => n442);
   U919 : NAND4_X1 port map( A1 => n994, A2 => n995, A3 => n996, A4 => n997, ZN
                           => n145_port);
   U920 : NAND2_X1 port map( A1 => n179, A2 => n263, ZN => n998);
   U921 : NAND2_X1 port map( A1 => n183, A2 => n264, ZN => n999);
   U922 : NAND2_X1 port map( A1 => n946, A2 => n298, ZN => n1000);
   U923 : AND3_X1 port map( A1 => n999, A2 => n998, A3 => n1000, ZN => n553);
   U924 : NOR4_X1 port map( A1 => n736, A2 => n739, A3 => n738, A4 => n737, ZN 
                           => n1001);
   U925 : AOI22_X1 port map( A1 => bht_17_23_port, A2 => n1096, B1 => n208, B2 
                           => bht_16_23_port, ZN => n781);
   U926 : AOI22_X1 port map( A1 => bht_31_23_port, A2 => n1095, B1 => 
                           bht_30_23_port, B2 => n1090, ZN => n788);
   U927 : AOI22_X1 port map( A1 => bht_29_16_port, A2 => n868, B1 => 
                           bht_28_16_port, B2 => n1085, ZN => n386);
   U928 : AOI22_X1 port map( A1 => bht_29_21_port, A2 => n1089, B1 => 
                           bht_28_21_port, B2 => n1085, ZN => n446);
   U929 : AOI22_X1 port map( A1 => bht_29_15_port, A2 => n1087, B1 => 
                           bht_28_15_port, B2 => n1085, ZN => n406);
   U930 : AOI22_X1 port map( A1 => bht_29_25_port, A2 => n867, B1 => 
                           bht_28_25_port, B2 => n1085, ZN => n500);
   U931 : AOI22_X1 port map( A1 => bht_29_11_port, A2 => n867, B1 => 
                           bht_28_11_port, B2 => n1086, ZN => n317);
   U932 : AOI22_X1 port map( A1 => bht_29_20_port, A2 => n1087, B1 => 
                           bht_28_20_port, B2 => n1085, ZN => n466);
   U933 : AOI22_X1 port map( A1 => bht_29_19_port, A2 => n1088, B1 => 
                           bht_28_19_port, B2 => n1084, ZN => n486);
   U934 : AOI22_X1 port map( A1 => bht_29_22_port, A2 => n868, B1 => 
                           bht_28_22_port, B2 => n1086, ZN => n426);
   U935 : AOI22_X1 port map( A1 => bht_29_26_port, A2 => n867, B1 => 
                           bht_28_26_port, B2 => n1086, ZN => n815);
   U936 : AND2_X1 port map( A1 => n844, A2 => n829, ZN => n231);
   U937 : AND2_X1 port map( A1 => n829, A2 => n850, ZN => n243);
   U938 : AOI22_X1 port map( A1 => bht_25_23_port, A2 => n1077, B1 => 
                           bht_24_23_port, B2 => n1073, ZN => n785);
   U939 : AOI22_X1 port map( A1 => bht_19_23_port, A2 => n1104, B1 => n1101, B2
                           => bht_18_23_port, ZN => n782);
   U940 : AND2_X1 port map( A1 => n1022, A2 => n1003, ZN => n1002);
   U941 : AND2_X1 port map( A1 => n1022, A2 => n1003, ZN => n249);
   U942 : AOI22_X1 port map( A1 => bht_27_23_port, A2 => n1083, B1 => 
                           bht_26_23_port, B2 => n1019, ZN => n786);
   U943 : NOR3_X1 port map( A1 => n929, A2 => n832, A3 => addr(6), ZN => n850);
   U944 : AOI22_X1 port map( A1 => bht_29_23_port, A2 => n1089, B1 => n1084, B2
                           => bht_28_23_port, ZN => n787);
   U945 : AOI22_X1 port map( A1 => bht_17_11_port, A2 => n1097, B1 => 
                           bht_16_11_port, B2 => n208, ZN => n311);
   U946 : AOI22_X1 port map( A1 => bht_17_25_port, A2 => n1097, B1 => n208, B2 
                           => bht_16_25_port, ZN => n494);
   U947 : AOI22_X1 port map( A1 => bht_17_16_port, A2 => n1097, B1 => 
                           bht_16_16_port, B2 => n208, ZN => n380);
   U948 : AOI22_X1 port map( A1 => bht_17_18_port, A2 => n1097, B1 => 
                           bht_16_18_port, B2 => n208, ZN => n339);
   U949 : AOI22_X1 port map( A1 => bht_17_21_port, A2 => n1097, B1 => 
                           bht_16_21_port, B2 => n208, ZN => n440);
   U950 : AOI22_X1 port map( A1 => bht_21_23_port, A2 => n1108, B1 => n865, B2 
                           => bht_20_23_port, ZN => n783);
   U951 : AOI22_X1 port map( A1 => bht_21_16_port, A2 => n1107, B1 => 
                           bht_20_16_port, B2 => n861, ZN => n382);
   U952 : AOI22_X1 port map( A1 => bht_21_11_port, A2 => n1109, B1 => 
                           bht_20_11_port, B2 => n865, ZN => n313);
   U953 : AOI22_X1 port map( A1 => bht_21_15_port, A2 => n1107, B1 => 
                           bht_20_15_port, B2 => n1015, ZN => n402);
   U954 : AOI22_X1 port map( A1 => bht_21_25_port, A2 => n1107, B1 => 
                           bht_20_25_port, B2 => n1015, ZN => n496);
   U955 : AOI22_X1 port map( A1 => bht_21_18_port, A2 => n1107, B1 => 
                           bht_20_18_port, B2 => n1014, ZN => n341);
   U956 : AND2_X1 port map( A1 => n1023, A2 => n1021, ZN => n1003);
   U957 : AOI22_X1 port map( A1 => n954, A2 => addr(28), B1 => n873, B2 => n959
                           , ZN => n144_port);
   U958 : AOI22_X1 port map( A1 => bht_13_1_port, A2 => n1041, B1 => 
                           bht_12_1_port, B2 => n1036, ZN => n237);
   U959 : AOI22_X1 port map( A1 => bht_13_25_port, A2 => n1039, B1 => 
                           bht_12_25_port, B2 => n1038, ZN => n508);
   U960 : AOI22_X1 port map( A1 => bht_13_3_port, A2 => n1039, B1 => 
                           bht_12_3_port, B2 => n876, ZN => n523);
   U961 : AOI22_X1 port map( A1 => bht_13_17_port, A2 => n1041, B1 => 
                           bht_12_17_port, B2 => n1038, ZN => n357);
   U962 : AOI22_X1 port map( A1 => bht_13_11_port, A2 => n1039, B1 => 
                           bht_12_11_port, B2 => n876, ZN => n325);
   U963 : AOI22_X1 port map( A1 => bht_13_19_port, A2 => n1040, B1 => 
                           bht_12_19_port, B2 => n1037, ZN => n478);
   U964 : AOI22_X1 port map( A1 => bht_13_22_port, A2 => n1041, B1 => 
                           bht_12_22_port, B2 => n876, ZN => n418);
   U965 : NAND4_X1 port map( A1 => n1004, A2 => n1005, A3 => n1006, A4 => n1007
                           , ZN => n143_port);
   U966 : AND2_X1 port map( A1 => n828, A2 => n837, ZN => n217);
   U967 : AOI22_X1 port map( A1 => bht_19_1_port, A2 => n1104, B1 => 
                           bht_18_1_port, B2 => n872, ZN => n195);
   U968 : AOI22_X1 port map( A1 => bht_19_3_port, A2 => n874, B1 => n1101, B2 
                           => bht_18_3_port, ZN => n526);
   U969 : AOI22_X1 port map( A1 => bht_19_17_port, A2 => n875, B1 => 
                           bht_18_17_port, B2 => n1101, ZN => n360);
   U970 : AOI22_X1 port map( A1 => bht_19_19_port, A2 => n1103, B1 => n1100, B2
                           => bht_18_19_port, ZN => n481);
   U971 : AOI22_X1 port map( A1 => bht_19_22_port, A2 => n1102, B1 => 
                           bht_18_22_port, B2 => n1101, ZN => n421);
   U972 : AOI22_X1 port map( A1 => bht_19_18_port, A2 => n874, B1 => 
                           bht_18_18_port, B2 => n1099, ZN => n340);
   U973 : AOI22_X1 port map( A1 => bht_19_25_port, A2 => n874, B1 => 
                           bht_18_25_port, B2 => n1101, ZN => n495);
   U974 : AOI22_X1 port map( A1 => bht_19_20_port, A2 => n1102, B1 => 
                           bht_18_20_port, B2 => n1099, ZN => n461);
   U975 : AOI22_X1 port map( A1 => bht_19_15_port, A2 => n875, B1 => 
                           bht_18_15_port, B2 => n1101, ZN => n401);
   U976 : AOI22_X1 port map( A1 => bht_19_11_port, A2 => n875, B1 => 
                           bht_18_11_port, B2 => n1099, ZN => n312);
   U977 : AOI22_X1 port map( A1 => bht_19_16_port, A2 => n1102, B1 => 
                           bht_18_16_port, B2 => n1099, ZN => n381);
   U978 : AOI22_X1 port map( A1 => bht_19_21_port, A2 => n1104, B1 => 
                           bht_18_21_port, B2 => n1099, ZN => n441);
   U979 : XNOR2_X1 port map( A => n1113, B => opcd(0), ZN => n1020);
   U980 : NAND3_X1 port map( A1 => rst, A2 => n91, A3 => opcd(2), ZN => n1010);
   U981 : NOR4_X1 port map( A1 => n1294, A2 => opcd(5), A3 => opcd(4), A4 => 
                           opcd(3), ZN => n91);
   U982 : NAND2_X1 port map( A1 => n1013, A2 => n1012, ZN => sig_brt_port);
   U983 : NAND2_X1 port map( A1 => N126, A2 => n961, ZN => n1012);
   U984 : NAND2_X1 port map( A1 => n249, A2 => n857, ZN => n1113);
   U985 : AOI22_X1 port map( A1 => bht_13_21_port, A2 => n1039, B1 => 
                           bht_12_21_port, B2 => n876, ZN => n438);
   U986 : AOI22_X1 port map( A1 => bht_13_16_port, A2 => n1041, B1 => 
                           bht_12_16_port, B2 => n1036, ZN => n378);
   U987 : AOI22_X1 port map( A1 => bht_13_15_port, A2 => n1041, B1 => 
                           bht_12_15_port, B2 => n1036, ZN => n398);
   U988 : AOI22_X1 port map( A1 => bht_13_20_port, A2 => n1039, B1 => 
                           bht_12_20_port, B2 => n876, ZN => n458);
   U989 : AOI22_X1 port map( A1 => bht_13_18_port, A2 => n1039, B1 => 
                           bht_12_18_port, B2 => n1036, ZN => n337);
   U990 : OAI222_X1 port map( A1 => n139_port, A2 => n292, B1 => n145_port, B2 
                           => n293, C1 => n878, C2 => n294, ZN => n756);
   U991 : AOI22_X1 port map( A1 => n954, A2 => addr(29), B1 => n878, B2 => n959
                           , ZN => n142_port);
   U992 : INV_X1 port map( A => n756, ZN => n248);
   U993 : AND4_X1 port map( A1 => n553, A2 => n1296, A3 => n1016, A4 => n1017, 
                           ZN => n301);
   U994 : XOR2_X1 port map( A => addr(7), B => n188_port, Z => n1016);
   U995 : XOR2_X1 port map( A => addr(8), B => n185, Z => n1017);
   U996 : AND2_X1 port map( A1 => n828, A2 => n843, ZN => n230);
   U997 : AND2_X1 port map( A1 => n830, A2 => n843, ZN => n234);
   U998 : AOI22_X1 port map( A1 => bht_27_1_port, A2 => n1081, B1 => 
                           bht_26_1_port, B2 => n1018, ZN => n210);
   U999 : AOI22_X1 port map( A1 => bht_27_3_port, A2 => n1081, B1 => 
                           bht_26_3_port, B2 => n1018, ZN => n530);
   U1000 : AOI22_X1 port map( A1 => bht_27_17_port, A2 => n1081, B1 => 
                           bht_26_17_port, B2 => n1079, ZN => n364);
   U1001 : AOI22_X1 port map( A1 => bht_27_19_port, A2 => n1081, B1 => 
                           bht_26_19_port, B2 => n1019, ZN => n485);
   U1002 : AOI22_X1 port map( A1 => bht_27_22_port, A2 => n1081, B1 => 
                           bht_26_22_port, B2 => n1080, ZN => n425);
   U1003 : AOI22_X1 port map( A1 => bht_27_18_port, A2 => n1081, B1 => 
                           bht_26_18_port, B2 => n1080, ZN => n344);
   U1004 : AOI22_X1 port map( A1 => bht_27_20_port, A2 => n1081, B1 => 
                           bht_26_20_port, B2 => n1018, ZN => n465);
   U1005 : AOI22_X1 port map( A1 => bht_27_15_port, A2 => n1081, B1 => 
                           bht_26_15_port, B2 => n1080, ZN => n405);
   U1006 : AOI22_X1 port map( A1 => bht_27_16_port, A2 => n1081, B1 => 
                           bht_26_16_port, B2 => n1018, ZN => n385);
   U1007 : AOI22_X1 port map( A1 => bht_27_21_port, A2 => n1081, B1 => 
                           bht_26_21_port, B2 => n1079, ZN => n445);
   U1008 : AOI22_X1 port map( A1 => bht_27_25_port, A2 => n1081, B1 => 
                           bht_26_25_port, B2 => n1019, ZN => n499);
   U1009 : AOI22_X1 port map( A1 => bht_27_11_port, A2 => n1081, B1 => 
                           bht_26_11_port, B2 => n1080, ZN => n316);
   U1010 : AOI22_X1 port map( A1 => bht_31_1_port, A2 => n1093, B1 => 
                           bht_30_1_port, B2 => n1092, ZN => n212);
   U1011 : AOI22_X1 port map( A1 => bht_31_3_port, A2 => n1093, B1 => 
                           bht_30_3_port, B2 => n1091, ZN => n532);
   U1012 : AOI22_X1 port map( A1 => bht_31_17_port, A2 => n1093, B1 => 
                           bht_30_17_port, B2 => n1091, ZN => n366);
   U1013 : AOI22_X1 port map( A1 => bht_31_19_port, A2 => n1093, B1 => 
                           bht_30_19_port, B2 => n1090, ZN => n487);
   U1014 : AOI22_X1 port map( A1 => bht_31_22_port, A2 => n1093, B1 => 
                           bht_30_22_port, B2 => n1091, ZN => n427);
   U1015 : AOI22_X1 port map( A1 => bht_31_18_port, A2 => n1093, B1 => 
                           bht_30_18_port, B2 => n1092, ZN => n346);
   U1016 : AOI22_X1 port map( A1 => bht_31_20_port, A2 => n1093, B1 => 
                           bht_30_20_port, B2 => n1092, ZN => n467);
   U1017 : AOI22_X1 port map( A1 => bht_31_15_port, A2 => n1093, B1 => 
                           bht_30_15_port, B2 => n1092, ZN => n407);
   U1018 : AOI22_X1 port map( A1 => bht_31_16_port, A2 => n1093, B1 => 
                           bht_30_16_port, B2 => n1091, ZN => n387);
   U1019 : AOI22_X1 port map( A1 => bht_31_21_port, A2 => n1093, B1 => 
                           bht_30_21_port, B2 => n1091, ZN => n447);
   U1020 : AOI22_X1 port map( A1 => bht_31_25_port, A2 => n1093, B1 => 
                           bht_30_25_port, B2 => n1091, ZN => n501);
   U1021 : AOI22_X1 port map( A1 => bht_31_11_port, A2 => n1093, B1 => 
                           bht_30_11_port, B2 => n1091, ZN => n318);
   U1022 : AOI22_X1 port map( A1 => bht_23_1_port, A2 => n1112, B1 => 
                           bht_22_1_port, B2 => n990, ZN => n197);
   U1023 : AOI22_X1 port map( A1 => bht_23_3_port, A2 => n1111, B1 => 
                           bht_22_3_port, B2 => n990, ZN => n528);
   U1024 : AOI22_X1 port map( A1 => bht_23_17_port, A2 => n1112, B1 => 
                           bht_22_17_port, B2 => n990, ZN => n362);
   U1025 : AOI22_X1 port map( A1 => bht_23_19_port, A2 => n1110, B1 => 
                           bht_22_19_port, B2 => n199, ZN => n483);
   U1026 : AOI22_X1 port map( A1 => bht_23_22_port, A2 => n1111, B1 => 
                           bht_22_22_port, B2 => n199, ZN => n423);
   U1027 : AOI22_X1 port map( A1 => bht_23_18_port, A2 => n1111, B1 => 
                           bht_22_18_port, B2 => n199, ZN => n342);
   U1028 : AOI22_X1 port map( A1 => bht_23_25_port, A2 => n1111, B1 => 
                           bht_22_25_port, B2 => n989, ZN => n497);
   U1029 : AOI22_X1 port map( A1 => bht_23_20_port, A2 => n1112, B1 => 
                           bht_22_20_port, B2 => n989, ZN => n463);
   U1030 : AOI22_X1 port map( A1 => bht_23_15_port, A2 => n1111, B1 => 
                           bht_22_15_port, B2 => n199, ZN => n403);
   U1031 : AOI22_X1 port map( A1 => bht_23_16_port, A2 => n1110, B1 => 
                           bht_22_16_port, B2 => n199, ZN => n383);
   U1032 : AOI22_X1 port map( A1 => bht_23_21_port, A2 => n1111, B1 => 
                           bht_22_21_port, B2 => n989, ZN => n443);
   U1033 : AOI22_X1 port map( A1 => bht_23_11_port, A2 => n1111, B1 => 
                           bht_22_11_port, B2 => n199, ZN => n314);
   U1034 : NAND4_X1 port map( A1 => n750, A2 => n749, A3 => n748, A4 => n751, 
                           ZN => n737);
   U1035 : NAND4_X1 port map( A1 => n752, A2 => n753, A3 => n754, A4 => n755, 
                           ZN => n736);
   U1036 : AOI22_X1 port map( A1 => n145_port, A2 => n293, B1 => n294, B2 => 
                           n143_port, ZN => n489);
   U1037 : AOI22_X1 port map( A1 => bht_23_23_port, A2 => n1110, B1 => 
                           bht_22_23_port, B2 => n989, ZN => n784);
   U1038 : NAND4_X1 port map( A1 => n742, A2 => n741, A3 => n740, A4 => n743, 
                           ZN => n739);
   U1039 : NAND4_X1 port map( A1 => n744, A2 => n745, A3 => n746, A4 => n747, 
                           ZN => n738);
   U1040 : OAI22_X1 port map( A1 => n956, A2 => n146_port, B1 => n147_port, B2 
                           => n954, ZN => N147);
   U1041 : AOI22_X1 port map( A1 => bht_5_1_port, A2 => n1065, B1 => 
                           bht_4_1_port, B2 => n965, ZN => n225);
   U1042 : AOI22_X1 port map( A1 => bht_5_25_port, A2 => n1064, B1 => 
                           bht_4_25_port, B2 => n1060, ZN => n504);
   U1043 : AOI22_X1 port map( A1 => bht_5_17_port, A2 => n1064, B1 => 
                           bht_4_17_port, B2 => n1061, ZN => n353);
   U1044 : AOI22_X1 port map( A1 => bht_5_19_port, A2 => n1063, B1 => 
                           bht_4_19_port, B2 => n1062, ZN => n474);
   U1045 : AOI22_X1 port map( A1 => bht_5_11_port, A2 => n1064, B1 => 
                           bht_4_11_port, B2 => n1060, ZN => n321);
   U1046 : AOI22_X1 port map( A1 => bht_5_18_port, A2 => n1064, B1 => 
                           bht_4_18_port, B2 => n1061, ZN => n333);
   U1047 : AOI22_X1 port map( A1 => bht_5_20_port, A2 => n1065, B1 => 
                           bht_4_20_port, B2 => n965, ZN => n454);
   U1048 : AOI22_X1 port map( A1 => bht_5_15_port, A2 => n1063, B1 => 
                           bht_4_15_port, B2 => n1061, ZN => n394);
   U1049 : AOI22_X1 port map( A1 => bht_5_3_port, A2 => n1064, B1 => 
                           bht_4_3_port, B2 => n1060, ZN => n519);
   U1050 : AOI22_X1 port map( A1 => bht_5_16_port, A2 => n1064, B1 => 
                           bht_4_16_port, B2 => n1060, ZN => n374);
   U1051 : AOI22_X1 port map( A1 => bht_5_21_port, A2 => n1064, B1 => 
                           bht_4_21_port, B2 => n1061, ZN => n434);
   U1052 : AOI22_X1 port map( A1 => bht_5_22_port, A2 => n1063, B1 => 
                           bht_4_22_port, B2 => n1061, ZN => n414);
   U1053 : AOI22_X1 port map( A1 => bht_13_13_port, A2 => n1039, B1 => 
                           bht_12_13_port, B2 => n1036, ZN => n654);
   U1054 : AOI22_X1 port map( A1 => bht_13_5_port, A2 => n1041, B1 => 
                           bht_12_5_port, B2 => n876, ZN => n734);
   U1055 : AOI22_X1 port map( A1 => bht_13_12_port, A2 => n1041, B1 => 
                           bht_12_12_port, B2 => n1036, ZN => n674);
   U1056 : AOI22_X1 port map( A1 => bht_13_14_port, A2 => n1041, B1 => 
                           bht_12_14_port, B2 => n1036, ZN => n714);
   U1057 : AOI22_X1 port map( A1 => bht_13_10_port, A2 => n1039, B1 => 
                           bht_12_10_port, B2 => n876, ZN => n694);
   U1058 : AOI22_X1 port map( A1 => bht_13_6_port, A2 => n1041, B1 => 
                           bht_12_6_port, B2 => n1036, ZN => n592);
   U1059 : AOI22_X1 port map( A1 => bht_13_8_port, A2 => n1039, B1 => 
                           bht_12_8_port, B2 => n1038, ZN => n634);
   U1060 : AOI22_X1 port map( A1 => bht_5_13_port, A2 => n1064, B1 => 
                           bht_4_13_port, B2 => n1060, ZN => n650);
   U1061 : AOI22_X1 port map( A1 => bht_5_5_port, A2 => n1064, B1 => 
                           bht_4_5_port, B2 => n1060, ZN => n730);
   U1062 : AOI22_X1 port map( A1 => bht_5_12_port, A2 => n1065, B1 => 
                           bht_4_12_port, B2 => n1060, ZN => n670);
   U1063 : AOI22_X1 port map( A1 => bht_5_14_port, A2 => n1065, B1 => 
                           bht_4_14_port, B2 => n1060, ZN => n710);
   U1064 : AOI22_X1 port map( A1 => bht_5_10_port, A2 => n1064, B1 => 
                           bht_4_10_port, B2 => n1060, ZN => n690);
   U1065 : AOI22_X1 port map( A1 => bht_5_6_port, A2 => n1065, B1 => 
                           bht_4_6_port, B2 => n1061, ZN => n588);
   U1066 : AOI22_X1 port map( A1 => bht_5_2_port, A2 => n1064, B1 => 
                           bht_4_2_port, B2 => n1061, ZN => n539);
   U1067 : AOI22_X1 port map( A1 => bht_5_8_port, A2 => n1064, B1 => 
                           bht_4_8_port, B2 => n1060, ZN => n630);
   U1068 : AOI22_X1 port map( A1 => bht_5_4_port, A2 => n1065, B1 => n1061, B2 
                           => bht_4_4_port, ZN => n568);
   U1069 : AOI22_X1 port map( A1 => bht_5_7_port, A2 => n1064, B1 => 
                           bht_4_7_port, B2 => n1061, ZN => n610);
   U1070 : AOI22_X1 port map( A1 => bht_5_9_port, A2 => n1063, B1 => 
                           bht_4_9_port, B2 => n1062, ZN => n742);
   U1071 : NAND2_X1 port map( A1 => n1001, A2 => n278, ZN => n1021);
   U1072 : NAND2_X1 port map( A1 => n279, A2 => n280, ZN => n1022);
   U1073 : NAND2_X1 port map( A1 => n281, A2 => n282, ZN => n1023);
   U1074 : INV_X1 port map( A => n298, ZN => n278);
   U1075 : NAND4_X1 port map( A1 => n284, A2 => n285, A3 => n286, A4 => n287, 
                           ZN => n280);
   U1076 : INV_X1 port map( A => n283, ZN => n282);
   U1077 : AOI22_X1 port map( A1 => bht_17_12_port, A2 => n1097, B1 => 
                           bht_16_12_port, B2 => n963, ZN => n660);
   U1078 : AOI22_X1 port map( A1 => bht_17_10_port, A2 => n1098, B1 => n208, B2
                           => bht_16_10_port, ZN => n680);
   U1079 : AOI22_X1 port map( A1 => bht_17_13_port, A2 => n1097, B1 => n798, B2
                           => bht_16_13_port, ZN => n640);
   U1080 : AOI22_X1 port map( A1 => bht_17_5_port, A2 => n1097, B1 => 
                           bht_16_5_port, B2 => n870, ZN => n720);
   U1081 : AOI22_X1 port map( A1 => bht_17_14_port, A2 => n1096, B1 => 
                           bht_16_14_port, B2 => n208, ZN => n700);
   U1082 : AOI22_X1 port map( A1 => bht_17_2_port, A2 => n1097, B1 => 
                           bht_16_2_port, B2 => n862, ZN => n545);
   U1083 : AOI22_X1 port map( A1 => bht_19_12_port, A2 => n1102, B1 => n1101, 
                           B2 => bht_18_12_port, ZN => n661);
   U1084 : AOI22_X1 port map( A1 => bht_19_10_port, A2 => n875, B1 => 
                           bht_18_10_port, B2 => n1099, ZN => n681);
   U1085 : AOI22_X1 port map( A1 => bht_19_13_port, A2 => n1104, B1 => 
                           bht_18_13_port, B2 => n1101, ZN => n641);
   U1086 : AOI22_X1 port map( A1 => bht_19_5_port, A2 => n874, B1 => 
                           bht_18_5_port, B2 => n1099, ZN => n721);
   U1087 : AOI22_X1 port map( A1 => bht_19_14_port, A2 => n875, B1 => n1100, B2
                           => bht_18_14_port, ZN => n701);
   U1088 : AOI22_X1 port map( A1 => bht_19_2_port, A2 => n1104, B1 => n1099, B2
                           => bht_18_2_port, ZN => n546);
   U1089 : AOI22_X1 port map( A1 => bht_19_6_port, A2 => n1104, B1 => 
                           bht_18_6_port, B2 => n1099, ZN => n579);
   U1090 : INV_X1 port map( A => addr(3), ZN => n851);
   U1091 : NOR2_X1 port map( A1 => addr(4), A2 => addr(3), ZN => n830);
   U1092 : AOI22_X1 port map( A1 => bht_13_24_port, A2 => n1041, B1 => 
                           bht_12_24_port, B2 => n1036, ZN => n775);
   U1093 : AOI22_X1 port map( A1 => bht_13_9_port, A2 => n1040, B1 => 
                           bht_12_9_port, B2 => n1037, ZN => n746);
   U1094 : AOI22_X1 port map( A1 => bht_13_7_port, A2 => n1041, B1 => 
                           bht_12_7_port, B2 => n876, ZN => n614);
   U1095 : AOI22_X1 port map( A1 => bht_13_2_port, A2 => n1041, B1 => 
                           bht_12_2_port, B2 => n876, ZN => n543);
   U1096 : AOI22_X1 port map( A1 => bht_13_4_port, A2 => n1039, B1 => 
                           bht_12_4_port, B2 => n1036, ZN => n572);
   U1097 : AOI22_X1 port map( A1 => bht_17_24_port, A2 => n1096, B1 => n208, B2
                           => bht_16_24_port, ZN => n761);
   U1098 : AOI22_X1 port map( A1 => bht_17_9_port, A2 => n1096, B1 => n208, B2 
                           => bht_16_9_port, ZN => n748);
   U1099 : AOI22_X1 port map( A1 => bht_17_7_port, A2 => n1098, B1 => 
                           bht_16_7_port, B2 => n870, ZN => n600);
   U1100 : AOI22_X1 port map( A1 => bht_17_4_port, A2 => n1097, B1 => 
                           bht_16_4_port, B2 => n208, ZN => n558);
   U1101 : AOI22_X1 port map( A1 => bht_17_8_port, A2 => n1097, B1 => 
                           bht_16_8_port, B2 => n208, ZN => n620);
   U1102 : AOI22_X1 port map( A1 => bht_25_12_port, A2 => n1076, B1 => 
                           bht_24_12_port, B2 => n1008, ZN => n664);
   U1103 : AOI22_X1 port map( A1 => bht_25_2_port, A2 => n1076, B1 => 
                           bht_24_2_port, B2 => n1074, ZN => n549);
   U1104 : AOI22_X1 port map( A1 => bht_25_6_port, A2 => n1076, B1 => 
                           bht_24_6_port, B2 => n1072, ZN => n582);
   U1105 : AOI22_X1 port map( A1 => bht_25_13_port, A2 => n1076, B1 => 
                           bht_24_13_port, B2 => n1009, ZN => n644);
   U1106 : AOI22_X1 port map( A1 => bht_25_5_port, A2 => n1076, B1 => 
                           bht_24_5_port, B2 => n1074, ZN => n724);
   U1107 : AOI22_X1 port map( A1 => bht_25_14_port, A2 => n1076, B1 => 
                           bht_24_14_port, B2 => n1072, ZN => n704);
   U1108 : AOI22_X1 port map( A1 => bht_25_10_port, A2 => n1076, B1 => 
                           bht_24_10_port, B2 => n1074, ZN => n684);
   U1109 : AOI22_X1 port map( A1 => bht_27_12_port, A2 => n1082, B1 => 
                           bht_26_12_port, B2 => n1018, ZN => n665);
   U1110 : AOI22_X1 port map( A1 => bht_27_2_port, A2 => n1082, B1 => 
                           bht_26_2_port, B2 => n1079, ZN => n550);
   U1111 : AOI22_X1 port map( A1 => bht_27_6_port, A2 => n1082, B1 => 
                           bht_26_6_port, B2 => n1018, ZN => n583);
   U1112 : AOI22_X1 port map( A1 => bht_27_13_port, A2 => n1082, B1 => 
                           bht_26_13_port, B2 => n1018, ZN => n645);
   U1113 : AOI22_X1 port map( A1 => bht_27_5_port, A2 => n1082, B1 => 
                           bht_26_5_port, B2 => n1079, ZN => n725);
   U1114 : AOI22_X1 port map( A1 => bht_27_14_port, A2 => n1082, B1 => 
                           bht_26_14_port, B2 => n1078, ZN => n705);
   U1115 : AOI22_X1 port map( A1 => bht_27_10_port, A2 => n1082, B1 => 
                           bht_26_10_port, B2 => n1080, ZN => n685);
   U1116 : AOI22_X1 port map( A1 => bht_25_24_port, A2 => n1076, B1 => n1073, 
                           B2 => bht_24_24_port, ZN => n765);
   U1117 : AOI22_X1 port map( A1 => bht_25_7_port, A2 => n1076, B1 => 
                           bht_24_7_port, B2 => n1073, ZN => n604);
   U1118 : AOI22_X1 port map( A1 => bht_25_4_port, A2 => n1076, B1 => 
                           bht_24_4_port, B2 => n1072, ZN => n562);
   U1119 : AOI22_X1 port map( A1 => bht_25_9_port, A2 => n1076, B1 => 
                           bht_24_9_port, B2 => n1072, ZN => n752);
   U1120 : AOI22_X1 port map( A1 => bht_25_8_port, A2 => n1076, B1 => 
                           bht_24_8_port, B2 => n1072, ZN => n624);
   U1121 : AOI22_X1 port map( A1 => bht_29_12_port, A2 => n1087, B1 => 
                           bht_28_12_port, B2 => n1085, ZN => n666);
   U1122 : AOI22_X1 port map( A1 => bht_29_2_port, A2 => n868, B1 => 
                           bht_28_2_port, B2 => n1086, ZN => n551);
   U1123 : AOI22_X1 port map( A1 => bht_29_6_port, A2 => n867, B1 => 
                           bht_28_6_port, B2 => n1085, ZN => n584);
   U1124 : AOI22_X1 port map( A1 => bht_29_13_port, A2 => n867, B1 => 
                           bht_28_13_port, B2 => n1085, ZN => n646);
   U1125 : AOI22_X1 port map( A1 => bht_29_5_port, A2 => n868, B1 => 
                           bht_28_5_port, B2 => n1085, ZN => n726);
   U1126 : AOI22_X1 port map( A1 => bht_29_14_port, A2 => n1088, B1 => 
                           bht_28_14_port, B2 => n1084, ZN => n706);
   U1127 : AOI22_X1 port map( A1 => bht_5_24_port, A2 => n1063, B1 => 
                           bht_4_24_port, B2 => n1061, ZN => n771);
   U1128 : AOI22_X1 port map( A1 => bht_31_12_port, A2 => n1094, B1 => 
                           bht_30_12_port, B2 => n1092, ZN => n667);
   U1129 : AOI22_X1 port map( A1 => bht_31_2_port, A2 => n1094, B1 => 
                           bht_30_2_port, B2 => n1091, ZN => n552);
   U1130 : AOI22_X1 port map( A1 => bht_31_6_port, A2 => n1094, B1 => 
                           bht_30_6_port, B2 => n1092, ZN => n585);
   U1131 : AOI22_X1 port map( A1 => bht_31_13_port, A2 => n1094, B1 => 
                           bht_30_13_port, B2 => n1091, ZN => n647);
   U1132 : AOI22_X1 port map( A1 => bht_31_5_port, A2 => n1094, B1 => 
                           bht_30_5_port, B2 => n1092, ZN => n727);
   U1133 : AOI22_X1 port map( A1 => bht_31_14_port, A2 => n1094, B1 => 
                           bht_30_14_port, B2 => n1090, ZN => n707);
   U1134 : AOI22_X1 port map( A1 => bht_31_10_port, A2 => n1094, B1 => 
                           bht_30_10_port, B2 => n1091, ZN => n687);
   U1135 : AOI22_X1 port map( A1 => bht_23_12_port, A2 => n1111, B1 => 
                           bht_22_12_port, B2 => n990, ZN => n663);
   U1136 : AOI22_X1 port map( A1 => bht_23_10_port, A2 => n1111, B1 => 
                           bht_22_10_port, B2 => n989, ZN => n683);
   U1137 : AOI22_X1 port map( A1 => bht_23_13_port, A2 => n1112, B1 => 
                           bht_22_13_port, B2 => n990, ZN => n643);
   U1138 : AOI22_X1 port map( A1 => bht_23_5_port, A2 => n1111, B1 => 
                           bht_22_5_port, B2 => n990, ZN => n723);
   U1139 : AOI22_X1 port map( A1 => bht_23_14_port, A2 => n1110, B1 => 
                           bht_22_14_port, B2 => n990, ZN => n703);
   U1140 : AOI22_X1 port map( A1 => bht_23_2_port, A2 => n1111, B1 => 
                           bht_22_2_port, B2 => n990, ZN => n548);
   U1141 : AOI22_X1 port map( A1 => bht_23_6_port, A2 => n1112, B1 => 
                           bht_22_6_port, B2 => n199, ZN => n581);
   U1142 : AOI22_X1 port map( A1 => bht_19_24_port, A2 => n1103, B1 => n1099, 
                           B2 => bht_18_24_port, ZN => n762);
   U1143 : AOI22_X1 port map( A1 => bht_19_9_port, A2 => n1103, B1 => n1100, B2
                           => bht_18_9_port, ZN => n749);
   U1144 : AOI22_X1 port map( A1 => bht_19_7_port, A2 => n875, B1 => 
                           bht_18_7_port, B2 => n1101, ZN => n601);
   U1145 : AOI22_X1 port map( A1 => bht_19_4_port, A2 => n1102, B1 => n1101, B2
                           => bht_18_4_port, ZN => n559);
   U1146 : AOI22_X1 port map( A1 => bht_19_8_port, A2 => n874, B1 => 
                           bht_18_8_port, B2 => n1101, ZN => n621);
   U1147 : AOI22_X1 port map( A1 => bht_27_24_port, A2 => n1082, B1 => n1019, 
                           B2 => bht_26_24_port, ZN => n766);
   U1148 : AOI22_X1 port map( A1 => bht_27_9_port, A2 => n1082, B1 => 
                           bht_26_9_port, B2 => n1079, ZN => n753);
   U1149 : AOI22_X1 port map( A1 => bht_27_4_port, A2 => n1082, B1 => 
                           bht_26_4_port, B2 => n1078, ZN => n563);
   U1150 : AOI22_X1 port map( A1 => bht_27_7_port, A2 => n1082, B1 => 
                           bht_26_7_port, B2 => n1079, ZN => n605);
   U1151 : AOI22_X1 port map( A1 => bht_27_8_port, A2 => n1082, B1 => 
                           bht_26_8_port, B2 => n1078, ZN => n625);
   U1152 : AOI22_X1 port map( A1 => bht_21_12_port, A2 => n1109, B1 => 
                           bht_20_12_port, B2 => n861, ZN => n662);
   U1153 : AOI22_X1 port map( A1 => bht_21_10_port, A2 => n1107, B1 => 
                           bht_20_10_port, B2 => n861, ZN => n682);
   U1154 : AOI22_X1 port map( A1 => bht_21_13_port, A2 => n1109, B1 => 
                           bht_20_13_port, B2 => n1015, ZN => n642);
   U1155 : AOI22_X1 port map( A1 => bht_21_5_port, A2 => n1107, B1 => 
                           bht_20_5_port, B2 => n1014, ZN => n722);
   U1156 : AOI22_X1 port map( A1 => bht_21_14_port, A2 => n1108, B1 => 
                           bht_20_14_port, B2 => n1105, ZN => n702);
   U1157 : AOI22_X1 port map( A1 => bht_21_2_port, A2 => n1107, B1 => 
                           bht_20_2_port, B2 => n1014, ZN => n547);
   U1158 : AOI22_X1 port map( A1 => bht_21_6_port, A2 => n1109, B1 => 
                           bht_20_6_port, B2 => n861, ZN => n580);
   U1159 : AOI22_X1 port map( A1 => bht_31_24_port, A2 => n1094, B1 => 
                           bht_30_24_port, B2 => n1090, ZN => n768);
   U1160 : AOI22_X1 port map( A1 => bht_31_9_port, A2 => n1094, B1 => 
                           bht_30_9_port, B2 => n1090, ZN => n755);
   U1161 : AOI22_X1 port map( A1 => bht_31_4_port, A2 => n1094, B1 => 
                           bht_30_4_port, B2 => n1091, ZN => n565);
   U1162 : AOI22_X1 port map( A1 => bht_31_7_port, A2 => n1094, B1 => 
                           bht_30_7_port, B2 => n1091, ZN => n607);
   U1163 : AOI22_X1 port map( A1 => bht_31_8_port, A2 => n1094, B1 => 
                           bht_30_8_port, B2 => n1090, ZN => n627);
   U1164 : AOI22_X1 port map( A1 => bht_23_24_port, A2 => n1110, B1 => 
                           bht_22_24_port, B2 => n199, ZN => n764);
   U1165 : AOI22_X1 port map( A1 => bht_23_9_port, A2 => n1110, B1 => 
                           bht_22_9_port, B2 => n990, ZN => n751);
   U1166 : AOI22_X1 port map( A1 => bht_23_4_port, A2 => n1111, B1 => 
                           bht_22_4_port, B2 => n199, ZN => n561);
   U1167 : AOI22_X1 port map( A1 => bht_23_7_port, A2 => n1111, B1 => 
                           bht_22_7_port, B2 => n989, ZN => n603);
   U1168 : AOI22_X1 port map( A1 => bht_23_8_port, A2 => n1111, B1 => 
                           bht_22_8_port, B2 => n989, ZN => n623);
   U1169 : AOI22_X1 port map( A1 => bht_29_24_port, A2 => n1088, B1 => 
                           bht_28_24_port, B2 => n1084, ZN => n767);
   U1170 : AOI22_X1 port map( A1 => bht_29_9_port, A2 => n1088, B1 => 
                           bht_28_9_port, B2 => n1084, ZN => n754);
   U1171 : AOI22_X1 port map( A1 => bht_29_4_port, A2 => n1087, B1 => 
                           bht_28_4_port, B2 => n1086, ZN => n564);
   U1172 : AOI22_X1 port map( A1 => bht_29_7_port, A2 => n1089, B1 => 
                           bht_28_7_port, B2 => n1086, ZN => n606);
   U1173 : AOI22_X1 port map( A1 => bht_29_8_port, A2 => n1088, B1 => 
                           bht_28_8_port, B2 => n1084, ZN => n626);
   U1174 : AOI22_X1 port map( A1 => bht_21_24_port, A2 => n1108, B1 => n1106, 
                           B2 => bht_20_24_port, ZN => n763);
   U1175 : AOI22_X1 port map( A1 => bht_21_9_port, A2 => n1108, B1 => n1105, B2
                           => bht_20_9_port, ZN => n750);
   U1176 : AOI22_X1 port map( A1 => bht_21_4_port, A2 => n1109, B1 => 
                           bht_20_4_port, B2 => n865, ZN => n560);
   U1177 : AOI22_X1 port map( A1 => bht_21_7_port, A2 => n1107, B1 => 
                           bht_20_7_port, B2 => n1106, ZN => n602);
   U1178 : AOI22_X1 port map( A1 => bht_21_8_port, A2 => n1108, B1 => 
                           bht_20_8_port, B2 => n1106, ZN => n622);
   U1179 : AND3_X1 port map( A1 => n831, A2 => n987, A3 => addr(6), ZN => n837)
                           ;
   U1180 : NOR3_X1 port map( A1 => n929, A2 => addr(6), A3 => addr(5), ZN => 
                           n844);
   U1181 : AOI22_X1 port map( A1 => n953, A2 => addr(31), B1 => n139_port, B2 
                           => n958, ZN => n137_port);
   U1182 : AOI22_X1 port map( A1 => n953, A2 => addr(16), B1 => n988, B2 => 
                           n958, ZN => n168);
   U1183 : AOI22_X1 port map( A1 => n953, A2 => addr(17), B1 => n167, B2 => 
                           n957, ZN => n166);
   U1184 : AOI22_X1 port map( A1 => n953, A2 => addr(9), B1 => n183, B2 => n958
                           , ZN => n182);
   U1185 : AOI22_X1 port map( A1 => n953, A2 => addr(18), B1 => n165, B2 => 
                           n957, ZN => n164);
   U1186 : AOI22_X1 port map( A1 => n953, A2 => addr(19), B1 => n163, B2 => 
                           n958, ZN => n162);
   U1187 : AOI22_X1 port map( A1 => n953, A2 => addr(10), B1 => n181, B2 => 
                           n957, ZN => n180);
   U1188 : AOI22_X1 port map( A1 => n953, A2 => addr(13), B1 => n175, B2 => 
                           n957, ZN => n174);
   U1189 : AOI22_X1 port map( A1 => n953, A2 => addr(11), B1 => n179, B2 => 
                           n956, ZN => n178);
   U1190 : AOI22_X1 port map( A1 => n953, A2 => addr(12), B1 => n177, B2 => 
                           n957, ZN => n176);
   U1191 : AOI22_X1 port map( A1 => n953, A2 => addr(14), B1 => n907, B2 => 
                           n959, ZN => n172);
   U1192 : AOI22_X1 port map( A1 => n953, A2 => addr(15), B1 => n171, B2 => 
                           n958, ZN => n170);
   U1193 : NOR3_X1 port map( A1 => n832, A2 => addr(6), A3 => addr(2), ZN => 
                           n849);
   U1194 : NOR3_X1 port map( A1 => addr(6), A2 => addr(5), A3 => addr(2), ZN =>
                           n843);
   U1195 : AND3_X1 port map( A1 => addr(2), A2 => addr(5), A3 => addr(6), ZN =>
                           n838);
   U1196 : INV_X1 port map( A => addr(2), ZN => n831);
   U1197 : AND4_X1 port map( A1 => n303, A2 => n304, A3 => n305, A4 => n306, ZN
                           => n302);
   U1198 : NAND4_X1 port map( A1 => n301, A2 => n302, A3 => n300, A4 => n299, 
                           ZN => n279);
   U1199 : INV_X1 port map( A => addr(5), ZN => n832);

end SYN_branch_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity StallGenerator_CWRD_SIZE20 is

   port( rst, clk, sig_ral, sig_bpw, sig_jral, sig_mul, sig_div, sig_sqrt : in 
         std_logic;  stall_flag : out std_logic_vector (4 downto 0));

end StallGenerator_CWRD_SIZE20;

architecture SYN_stall_generator_arch of StallGenerator_CWRD_SIZE20 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component StallGenerator_CWRD_SIZE20_DW01_inc_5
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component StallGenerator_CWRD_SIZE20_DW01_inc_4
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component StallGenerator_CWRD_SIZE20_DW01_inc_3
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component StallGenerator_CWRD_SIZE20_DW01_inc_2
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component StallGenerator_CWRD_SIZE20_DW01_inc_1
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component StallGenerator_CWRD_SIZE20_DW01_inc_0
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal stall_flag_3_port, stall_flag_2_port, stall_flag_1_port, 
      stall_flag_0_port, n_state_ral_31_port, n_state_ral_30_port, 
      n_state_ral_29_port, n_state_ral_28_port, n_state_ral_27_port, 
      n_state_ral_26_port, n_state_ral_25_port, n_state_ral_24_port, 
      n_state_ral_23_port, n_state_ral_22_port, n_state_ral_21_port, 
      n_state_ral_20_port, n_state_ral_19_port, n_state_ral_18_port, 
      n_state_ral_17_port, n_state_ral_16_port, n_state_ral_15_port, 
      n_state_ral_14_port, n_state_ral_13_port, n_state_ral_12_port, 
      n_state_ral_11_port, n_state_ral_10_port, n_state_ral_9_port, 
      n_state_ral_8_port, n_state_ral_7_port, n_state_ral_6_port, 
      n_state_ral_5_port, n_state_ral_4_port, n_state_ral_3_port, 
      n_state_ral_2_port, n_state_ral_1_port, n_state_ral_0_port, 
      c_state_ral_31_port, c_state_ral_30_port, c_state_ral_29_port, 
      c_state_ral_28_port, c_state_ral_27_port, c_state_ral_26_port, 
      c_state_ral_25_port, c_state_ral_24_port, c_state_ral_23_port, 
      c_state_ral_22_port, c_state_ral_21_port, c_state_ral_20_port, 
      c_state_ral_19_port, c_state_ral_18_port, c_state_ral_17_port, 
      c_state_ral_16_port, c_state_ral_15_port, c_state_ral_14_port, 
      c_state_ral_13_port, c_state_ral_12_port, c_state_ral_11_port, 
      c_state_ral_10_port, c_state_ral_9_port, c_state_ral_8_port, 
      c_state_ral_7_port, c_state_ral_6_port, c_state_ral_5_port, 
      c_state_ral_4_port, c_state_ral_3_port, c_state_ral_2_port, 
      c_state_ral_1_port, c_state_ral_0_port, N46, N47, N48, N49, N50, N51, N52
      , N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, 
      N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, 
      n_state_bpw_31_port, n_state_bpw_30_port, n_state_bpw_29_port, 
      n_state_bpw_28_port, n_state_bpw_27_port, n_state_bpw_26_port, 
      n_state_bpw_25_port, n_state_bpw_24_port, n_state_bpw_23_port, 
      n_state_bpw_22_port, n_state_bpw_21_port, n_state_bpw_20_port, 
      n_state_bpw_19_port, n_state_bpw_18_port, n_state_bpw_17_port, 
      n_state_bpw_16_port, n_state_bpw_15_port, n_state_bpw_14_port, 
      n_state_bpw_13_port, n_state_bpw_12_port, n_state_bpw_11_port, 
      n_state_bpw_10_port, n_state_bpw_9_port, n_state_bpw_8_port, 
      n_state_bpw_7_port, n_state_bpw_6_port, n_state_bpw_5_port, 
      n_state_bpw_4_port, n_state_bpw_3_port, n_state_bpw_2_port, 
      n_state_bpw_1_port, n_state_bpw_0_port, c_state_bpw_31_port, 
      c_state_bpw_30_port, c_state_bpw_29_port, c_state_bpw_28_port, 
      c_state_bpw_27_port, c_state_bpw_26_port, c_state_bpw_25_port, 
      c_state_bpw_24_port, c_state_bpw_23_port, c_state_bpw_22_port, 
      c_state_bpw_21_port, c_state_bpw_20_port, c_state_bpw_19_port, 
      c_state_bpw_18_port, c_state_bpw_17_port, c_state_bpw_16_port, 
      c_state_bpw_15_port, c_state_bpw_14_port, c_state_bpw_13_port, 
      c_state_bpw_12_port, c_state_bpw_11_port, c_state_bpw_10_port, 
      c_state_bpw_9_port, c_state_bpw_8_port, c_state_bpw_7_port, 
      c_state_bpw_6_port, c_state_bpw_5_port, c_state_bpw_4_port, 
      c_state_bpw_3_port, c_state_bpw_2_port, c_state_bpw_1_port, 
      c_state_bpw_0_port, N119, N120, N121, N122, N123, N124, N125, N126, N127,
      N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139, 
      N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, 
      c_state_mul_31_port, c_state_mul_30_port, c_state_mul_29_port, 
      c_state_mul_28_port, c_state_mul_27_port, c_state_mul_26_port, 
      c_state_mul_25_port, c_state_mul_24_port, c_state_mul_23_port, 
      c_state_mul_22_port, c_state_mul_21_port, c_state_mul_20_port, 
      c_state_mul_19_port, c_state_mul_18_port, c_state_mul_17_port, 
      c_state_mul_16_port, c_state_mul_15_port, c_state_mul_14_port, 
      c_state_mul_13_port, c_state_mul_12_port, c_state_mul_11_port, 
      c_state_mul_10_port, c_state_mul_9_port, c_state_mul_8_port, 
      c_state_mul_7_port, c_state_mul_6_port, c_state_mul_5_port, 
      c_state_mul_4_port, c_state_mul_3_port, c_state_mul_2_port, 
      c_state_mul_1_port, c_state_mul_0_port, n_state_mul_31_port, 
      n_state_mul_30_port, n_state_mul_29_port, n_state_mul_28_port, 
      n_state_mul_27_port, n_state_mul_26_port, n_state_mul_25_port, 
      n_state_mul_24_port, n_state_mul_23_port, n_state_mul_22_port, 
      n_state_mul_21_port, n_state_mul_20_port, n_state_mul_19_port, 
      n_state_mul_18_port, n_state_mul_17_port, n_state_mul_16_port, 
      n_state_mul_15_port, n_state_mul_14_port, n_state_mul_13_port, 
      n_state_mul_12_port, n_state_mul_11_port, n_state_mul_10_port, 
      n_state_mul_9_port, n_state_mul_8_port, n_state_mul_7_port, 
      n_state_mul_6_port, n_state_mul_5_port, n_state_mul_4_port, 
      n_state_mul_3_port, n_state_mul_2_port, n_state_mul_1_port, 
      n_state_mul_0_port, N193, N194, N195, N196, N197, N198, N199, N200, N201,
      N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, 
      N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, 
      c_state_div_31_port, c_state_div_30_port, c_state_div_29_port, 
      c_state_div_28_port, c_state_div_27_port, c_state_div_26_port, 
      c_state_div_25_port, c_state_div_24_port, c_state_div_23_port, 
      c_state_div_22_port, c_state_div_21_port, c_state_div_20_port, 
      c_state_div_19_port, c_state_div_18_port, c_state_div_17_port, 
      c_state_div_16_port, c_state_div_15_port, c_state_div_14_port, 
      c_state_div_13_port, c_state_div_12_port, c_state_div_11_port, 
      c_state_div_10_port, c_state_div_9_port, c_state_div_8_port, 
      c_state_div_7_port, c_state_div_6_port, c_state_div_5_port, 
      c_state_div_4_port, c_state_div_3_port, c_state_div_2_port, 
      c_state_div_1_port, c_state_div_0_port, n_state_div_31_port, 
      n_state_div_30_port, n_state_div_29_port, n_state_div_28_port, 
      n_state_div_27_port, n_state_div_26_port, n_state_div_25_port, 
      n_state_div_24_port, n_state_div_23_port, n_state_div_22_port, 
      n_state_div_21_port, n_state_div_20_port, n_state_div_19_port, 
      n_state_div_18_port, n_state_div_17_port, n_state_div_16_port, 
      n_state_div_15_port, n_state_div_14_port, n_state_div_13_port, 
      n_state_div_12_port, n_state_div_11_port, n_state_div_10_port, 
      n_state_div_9_port, n_state_div_8_port, n_state_div_7_port, 
      n_state_div_6_port, n_state_div_5_port, n_state_div_4_port, 
      n_state_div_3_port, n_state_div_2_port, n_state_div_1_port, 
      n_state_div_0_port, N278, N279, N280, N281, N282, N283, N284, N285, N286,
      N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, 
      N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N309, 
      c_state_sqrt_31_port, c_state_sqrt_30_port, c_state_sqrt_29_port, 
      c_state_sqrt_28_port, c_state_sqrt_27_port, c_state_sqrt_26_port, 
      c_state_sqrt_25_port, c_state_sqrt_24_port, c_state_sqrt_23_port, 
      c_state_sqrt_22_port, c_state_sqrt_21_port, c_state_sqrt_20_port, 
      c_state_sqrt_19_port, c_state_sqrt_18_port, c_state_sqrt_17_port, 
      c_state_sqrt_16_port, c_state_sqrt_15_port, c_state_sqrt_14_port, 
      c_state_sqrt_13_port, c_state_sqrt_12_port, c_state_sqrt_11_port, 
      c_state_sqrt_10_port, c_state_sqrt_9_port, c_state_sqrt_8_port, 
      c_state_sqrt_7_port, c_state_sqrt_6_port, c_state_sqrt_5_port, 
      c_state_sqrt_4_port, c_state_sqrt_3_port, c_state_sqrt_2_port, 
      c_state_sqrt_1_port, c_state_sqrt_0_port, n_state_sqrt_31_port, 
      n_state_sqrt_30_port, n_state_sqrt_29_port, n_state_sqrt_28_port, 
      n_state_sqrt_27_port, n_state_sqrt_26_port, n_state_sqrt_25_port, 
      n_state_sqrt_24_port, n_state_sqrt_23_port, n_state_sqrt_22_port, 
      n_state_sqrt_21_port, n_state_sqrt_20_port, n_state_sqrt_19_port, 
      n_state_sqrt_18_port, n_state_sqrt_17_port, n_state_sqrt_16_port, 
      n_state_sqrt_15_port, n_state_sqrt_14_port, n_state_sqrt_13_port, 
      n_state_sqrt_12_port, n_state_sqrt_11_port, n_state_sqrt_10_port, 
      n_state_sqrt_9_port, n_state_sqrt_8_port, n_state_sqrt_7_port, 
      n_state_sqrt_6_port, n_state_sqrt_5_port, n_state_sqrt_4_port, 
      n_state_sqrt_3_port, n_state_sqrt_2_port, n_state_sqrt_1_port, 
      n_state_sqrt_0_port, N363, N364, N365, N366, N367, N368, N369, N370, N371
      , N372, N373, N374, N375, N376, N377, N378, N379, N380, N381, N382, N383,
      N384, N385, N386, N387, N388, N389, N390, N391, N392, N393, N394, 
      c_state_stu_31_port, c_state_stu_30_port, c_state_stu_29_port, 
      c_state_stu_28_port, c_state_stu_27_port, c_state_stu_26_port, 
      c_state_stu_25_port, c_state_stu_24_port, c_state_stu_23_port, 
      c_state_stu_22_port, c_state_stu_21_port, c_state_stu_20_port, 
      c_state_stu_19_port, c_state_stu_18_port, c_state_stu_17_port, 
      c_state_stu_16_port, c_state_stu_15_port, c_state_stu_14_port, 
      c_state_stu_13_port, c_state_stu_12_port, c_state_stu_11_port, 
      c_state_stu_10_port, c_state_stu_9_port, c_state_stu_8_port, 
      c_state_stu_7_port, c_state_stu_6_port, c_state_stu_5_port, 
      c_state_stu_4_port, c_state_stu_3_port, c_state_stu_2_port, 
      c_state_stu_1_port, c_state_stu_0_port, n_state_stu_31_port, 
      n_state_stu_30_port, n_state_stu_29_port, n_state_stu_28_port, 
      n_state_stu_27_port, n_state_stu_26_port, n_state_stu_25_port, 
      n_state_stu_24_port, n_state_stu_23_port, n_state_stu_22_port, 
      n_state_stu_21_port, n_state_stu_20_port, n_state_stu_19_port, 
      n_state_stu_18_port, n_state_stu_17_port, n_state_stu_16_port, 
      n_state_stu_15_port, n_state_stu_14_port, n_state_stu_13_port, 
      n_state_stu_12_port, n_state_stu_11_port, n_state_stu_10_port, 
      n_state_stu_9_port, n_state_stu_8_port, n_state_stu_7_port, 
      n_state_stu_6_port, n_state_stu_5_port, n_state_stu_4_port, 
      n_state_stu_3_port, n_state_stu_2_port, n_state_stu_1_port, 
      n_state_stu_0_port, N444, N445, N446, N447, N448, N449, N450, N451, N452,
      N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, 
      N465, N466, N467, N468, N469, N470, N471, N472, N473, N474, N475, n192, 
      n194_port, n195_port, n197_port, n214_port, n222_port, n230, n231, n232, 
      n247, n261, n262, n263, n266, n276, n294_port, n307_port, n308_port, 
      n309_port, n310, n311, n312, n342, n343, n344, n347, n348, n155, n157, 
      n158, n159, n160, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n180, n181, n182, n183, n185, n186, n187, 
      n188, n189, n190, n191, n193_port, n196_port, n198_port, n199_port, 
      n200_port, n201_port, n205_port, n206_port, n207_port, n208_port, 
      n210_port, n211_port, n212_port, n213_port, n218_port, n219_port, 
      n220_port, n221_port, n226, n227, n228, n229, n233, n234, n235, n239, 
      n240, n241, n242, n243, n244, n249, net107995, net107996, net107997, 
      net107998, net107999, net108000, net108001, net108002, net108003, 
      net108004, net108005, net108006, net108007, net108008, net108009, 
      net108010, net108011, net108012, net108013, net108014, net108015, 
      net108016, net108017, net108018, net108019, net108020, net108021, 
      net108022, net108023, net108024, net108025, net108026, net108027, 
      net108028, net108029, net108030, net108031, net108032, net108033, 
      net108034, net108035, net108036, net108037, net108038, net108039, 
      net108040, net108041, net108042, net108043, net108044, net108045, 
      net108046, net108047, net108048, net108049, net108050, net108051, 
      net108052, net108053, net108054, net108055, net108056, net108057, 
      net108058, net108059, net108060, net108061, net108062, net108063, n37, 
      n38, n39, n41, n42, n43, n44, n45, n46_port, n47_port, n48_port, n49_port
      , n50_port, n52_port, n53_port, n54_port, n55_port, n56_port, n57_port, 
      n58_port, n59_port, n60_port, n62_port, n63_port, n65_port, n66_port, 
      n67_port, n68_port, n69_port, n70_port, n71_port, n72_port, n75_port, 
      n76_port, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90
      , n94, n95, n96, n100, n101, n102, n103, n104, n105, n107, n108, n109, 
      n110, n111, n112, n113, n114, n115, n116, n117, n118, n119_port, 
      n120_port, n122_port, n123_port, n124_port, n125_port, n126_port, 
      n127_port, n128_port, n129_port, n130_port, n131_port, n132_port, 
      n133_port, n134_port, n135_port, n137_port, n138_port, n139_port, 
      n140_port, n141_port, n142_port, n143_port, n144_port, n145_port, 
      n146_port, n147_port, n148_port, n149_port, n150_port, n151, n152, n153, 
      n154, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, 
      n265, n268, n269, n270, n272, n273, n274, n275, n277, n278_port, 
      n279_port, n280_port, n281_port, n282_port, n283_port, n284_port, 
      n285_port, n286_port, n287_port, n288_port, n289_port, n290_port, n264, 
      n267, n271, n291_port, n292_port, n293_port, n295_port, n296_port, 
      n297_port, n298_port, n299_port, n300_port, n301_port, n302_port, 
      n303_port, n304_port, n305_port, n306_port, n313, n314, n315, n316, n317,
      n318, n319, n320, n321, n322, n323, n324, n325, net163713, net163714, 
      net163715, net163716, net163717, net163718, net163719, net163720, 
      net163721, net163722, net163723, net163724, net163725, net163726, 
      net163727, net163728, net163729, net163730, net163731, net163732, 
      net163733, net163734, net163735, net163736, net163737, net163738, 
      net163739, net163740, net163741, net163742, net163743, net163744, 
      net163745, net163746 : std_logic;

begin
   stall_flag <= ( stall_flag_3_port, stall_flag_3_port, stall_flag_2_port, 
      stall_flag_1_port, stall_flag_0_port );
   
   c_state_ral_reg_0_inst : DFFR_X1 port map( D => n_state_ral_0_port, CK => 
                           clk, RN => n317, Q => c_state_ral_0_port, QN => 
                           n195_port);
   c_state_ral_reg_10_inst : DFFR_X1 port map( D => n_state_ral_10_port, CK => 
                           clk, RN => n316, Q => c_state_ral_10_port, QN => 
                           net108063);
   c_state_ral_reg_1_inst : DFFR_X1 port map( D => n_state_ral_1_port, CK => 
                           clk, RN => n315, Q => c_state_ral_1_port, QN => n231
                           );
   c_state_ral_reg_2_inst : DFFR_X1 port map( D => n_state_ral_2_port, CK => 
                           clk, RN => n315, Q => c_state_ral_2_port, QN => 
                           net108062);
   c_state_ral_reg_3_inst : DFFR_X1 port map( D => n_state_ral_3_port, CK => 
                           clk, RN => n315, Q => c_state_ral_3_port, QN => 
                           net108061);
   c_state_ral_reg_4_inst : DFFR_X1 port map( D => n_state_ral_4_port, CK => 
                           clk, RN => n315, Q => c_state_ral_4_port, QN => 
                           net163746);
   c_state_ral_reg_5_inst : DFFR_X1 port map( D => n_state_ral_5_port, CK => 
                           clk, RN => n315, Q => c_state_ral_5_port, QN => 
                           n208_port);
   c_state_ral_reg_6_inst : DFFR_X1 port map( D => n_state_ral_6_port, CK => 
                           clk, RN => n315, Q => c_state_ral_6_port, QN => 
                           n207_port);
   c_state_ral_reg_7_inst : DFFR_X1 port map( D => n_state_ral_7_port, CK => 
                           clk, RN => n315, Q => c_state_ral_7_port, QN => 
                           n206_port);
   c_state_ral_reg_8_inst : DFFR_X1 port map( D => n_state_ral_8_port, CK => 
                           clk, RN => n315, Q => c_state_ral_8_port, QN => 
                           net108060);
   c_state_ral_reg_9_inst : DFFR_X1 port map( D => n_state_ral_9_port, CK => 
                           clk, RN => n317, Q => c_state_ral_9_port, QN => 
                           net108059);
   c_state_ral_reg_11_inst : DFFR_X1 port map( D => n_state_ral_11_port, CK => 
                           clk, RN => n316, Q => c_state_ral_11_port, QN => 
                           net108058);
   c_state_ral_reg_12_inst : DFFR_X1 port map( D => n_state_ral_12_port, CK => 
                           clk, RN => n316, Q => c_state_ral_12_port, QN => 
                           n205_port);
   c_state_ral_reg_13_inst : DFFR_X1 port map( D => n_state_ral_13_port, CK => 
                           clk, RN => n316, Q => c_state_ral_13_port, QN => 
                           net163745);
   c_state_ral_reg_14_inst : DFFR_X1 port map( D => n_state_ral_14_port, CK => 
                           clk, RN => n316, Q => c_state_ral_14_port, QN => 
                           net163744);
   c_state_ral_reg_15_inst : DFFR_X1 port map( D => n_state_ral_15_port, CK => 
                           clk, RN => n316, Q => c_state_ral_15_port, QN => 
                           net163743);
   c_state_ral_reg_16_inst : DFFR_X1 port map( D => n_state_ral_16_port, CK => 
                           clk, RN => n316, Q => c_state_ral_16_port, QN => 
                           net108057);
   c_state_ral_reg_17_inst : DFFR_X1 port map( D => n_state_ral_17_port, CK => 
                           clk, RN => n316, Q => c_state_ral_17_port, QN => 
                           net108056);
   c_state_ral_reg_18_inst : DFFR_X1 port map( D => n_state_ral_18_port, CK => 
                           clk, RN => n316, Q => c_state_ral_18_port, QN => 
                           net108055);
   c_state_ral_reg_19_inst : DFFR_X1 port map( D => n_state_ral_19_port, CK => 
                           clk, RN => n316, Q => c_state_ral_19_port, QN => 
                           n201_port);
   c_state_ral_reg_20_inst : DFFR_X1 port map( D => n_state_ral_20_port, CK => 
                           clk, RN => n316, Q => c_state_ral_20_port, QN => 
                           n200_port);
   c_state_ral_reg_21_inst : DFFR_X1 port map( D => n_state_ral_21_port, CK => 
                           clk, RN => n316, Q => c_state_ral_21_port, QN => 
                           n199_port);
   c_state_ral_reg_22_inst : DFFR_X1 port map( D => n_state_ral_22_port, CK => 
                           clk, RN => n317, Q => c_state_ral_22_port, QN => 
                           n198_port);
   c_state_ral_reg_23_inst : DFFR_X1 port map( D => n_state_ral_23_port, CK => 
                           clk, RN => n317, Q => c_state_ral_23_port, QN => 
                           n196_port);
   c_state_ral_reg_24_inst : DFFR_X1 port map( D => n_state_ral_24_port, CK => 
                           clk, RN => n317, Q => c_state_ral_24_port, QN => 
                           n193_port);
   c_state_ral_reg_25_inst : DFFR_X1 port map( D => n_state_ral_25_port, CK => 
                           clk, RN => n317, Q => c_state_ral_25_port, QN => 
                           n191);
   c_state_ral_reg_26_inst : DFFR_X1 port map( D => n_state_ral_26_port, CK => 
                           clk, RN => n317, Q => c_state_ral_26_port, QN => 
                           n190);
   c_state_ral_reg_27_inst : DFFR_X1 port map( D => n_state_ral_27_port, CK => 
                           clk, RN => n317, Q => c_state_ral_27_port, QN => 
                           n189);
   c_state_ral_reg_28_inst : DFFR_X1 port map( D => n_state_ral_28_port, CK => 
                           clk, RN => n317, Q => c_state_ral_28_port, QN => 
                           n188);
   c_state_ral_reg_29_inst : DFFR_X1 port map( D => n_state_ral_29_port, CK => 
                           clk, RN => n317, Q => c_state_ral_29_port, QN => 
                           n187);
   c_state_ral_reg_30_inst : DFFR_X1 port map( D => n_state_ral_30_port, CK => 
                           clk, RN => n317, Q => c_state_ral_30_port, QN => 
                           n186);
   c_state_ral_reg_31_inst : DFFR_X1 port map( D => n_state_ral_31_port, CK => 
                           clk, RN => n317, Q => c_state_ral_31_port, QN => 
                           n185);
   c_state_bpw_reg_0_inst : DFFR_X1 port map( D => n_state_bpw_0_port, CK => 
                           clk, RN => n306_port, Q => c_state_bpw_0_port, QN =>
                           n197_port);
   c_state_bpw_reg_10_inst : DFFR_X1 port map( D => n_state_bpw_10_port, CK => 
                           clk, RN => n304_port, Q => c_state_bpw_10_port, QN 
                           => net108054);
   c_state_bpw_reg_1_inst : DFFR_X1 port map( D => n_state_bpw_1_port, CK => 
                           clk, RN => n304_port, Q => c_state_bpw_1_port, QN =>
                           n232);
   c_state_bpw_reg_2_inst : DFFR_X1 port map( D => n_state_bpw_2_port, CK => 
                           clk, RN => n304_port, Q => c_state_bpw_2_port, QN =>
                           net108053);
   c_state_bpw_reg_3_inst : DFFR_X1 port map( D => n_state_bpw_3_port, CK => 
                           clk, RN => n304_port, Q => c_state_bpw_3_port, QN =>
                           net108052);
   c_state_bpw_reg_4_inst : DFFR_X1 port map( D => n_state_bpw_4_port, CK => 
                           clk, RN => n304_port, Q => c_state_bpw_4_port, QN =>
                           net163742);
   c_state_bpw_reg_5_inst : DFFR_X1 port map( D => n_state_bpw_5_port, CK => 
                           clk, RN => n304_port, Q => c_state_bpw_5_port, QN =>
                           n183);
   c_state_bpw_reg_6_inst : DFFR_X1 port map( D => n_state_bpw_6_port, CK => 
                           clk, RN => n304_port, Q => c_state_bpw_6_port, QN =>
                           n182);
   c_state_bpw_reg_7_inst : DFFR_X1 port map( D => n_state_bpw_7_port, CK => 
                           clk, RN => n304_port, Q => c_state_bpw_7_port, QN =>
                           n181);
   c_state_bpw_reg_8_inst : DFFR_X1 port map( D => n_state_bpw_8_port, CK => 
                           clk, RN => n304_port, Q => c_state_bpw_8_port, QN =>
                           net108051);
   c_state_bpw_reg_9_inst : DFFR_X1 port map( D => n_state_bpw_9_port, CK => 
                           clk, RN => n306_port, Q => c_state_bpw_9_port, QN =>
                           net108050);
   c_state_bpw_reg_11_inst : DFFR_X1 port map( D => n_state_bpw_11_port, CK => 
                           clk, RN => n304_port, Q => c_state_bpw_11_port, QN 
                           => net108049);
   c_state_bpw_reg_12_inst : DFFR_X1 port map( D => n_state_bpw_12_port, CK => 
                           clk, RN => n304_port, Q => c_state_bpw_12_port, QN 
                           => n180);
   c_state_bpw_reg_13_inst : DFFR_X1 port map( D => n_state_bpw_13_port, CK => 
                           clk, RN => n304_port, Q => c_state_bpw_13_port, QN 
                           => net163741);
   c_state_bpw_reg_14_inst : DFFR_X1 port map( D => n_state_bpw_14_port, CK => 
                           clk, RN => n305_port, Q => c_state_bpw_14_port, QN 
                           => net163740);
   c_state_bpw_reg_15_inst : DFFR_X1 port map( D => n_state_bpw_15_port, CK => 
                           clk, RN => n305_port, Q => c_state_bpw_15_port, QN 
                           => net163739);
   c_state_bpw_reg_16_inst : DFFR_X1 port map( D => n_state_bpw_16_port, CK => 
                           clk, RN => n305_port, Q => c_state_bpw_16_port, QN 
                           => net108048);
   c_state_bpw_reg_17_inst : DFFR_X1 port map( D => n_state_bpw_17_port, CK => 
                           clk, RN => n305_port, Q => c_state_bpw_17_port, QN 
                           => net108047);
   c_state_bpw_reg_18_inst : DFFR_X1 port map( D => n_state_bpw_18_port, CK => 
                           clk, RN => n305_port, Q => c_state_bpw_18_port, QN 
                           => net108046);
   c_state_bpw_reg_19_inst : DFFR_X1 port map( D => n_state_bpw_19_port, CK => 
                           clk, RN => n305_port, Q => c_state_bpw_19_port, QN 
                           => n176);
   c_state_bpw_reg_20_inst : DFFR_X1 port map( D => n_state_bpw_20_port, CK => 
                           clk, RN => n305_port, Q => c_state_bpw_20_port, QN 
                           => n175);
   c_state_bpw_reg_21_inst : DFFR_X1 port map( D => n_state_bpw_21_port, CK => 
                           clk, RN => n305_port, Q => c_state_bpw_21_port, QN 
                           => n174);
   c_state_bpw_reg_22_inst : DFFR_X1 port map( D => n_state_bpw_22_port, CK => 
                           clk, RN => n305_port, Q => c_state_bpw_22_port, QN 
                           => n173);
   c_state_bpw_reg_23_inst : DFFR_X1 port map( D => n_state_bpw_23_port, CK => 
                           clk, RN => n305_port, Q => c_state_bpw_23_port, QN 
                           => n172);
   c_state_bpw_reg_24_inst : DFFR_X1 port map( D => n_state_bpw_24_port, CK => 
                           clk, RN => n305_port, Q => c_state_bpw_24_port, QN 
                           => n171);
   c_state_bpw_reg_25_inst : DFFR_X1 port map( D => n_state_bpw_25_port, CK => 
                           clk, RN => n305_port, Q => c_state_bpw_25_port, QN 
                           => n170);
   c_state_bpw_reg_26_inst : DFFR_X1 port map( D => n_state_bpw_26_port, CK => 
                           clk, RN => n306_port, Q => c_state_bpw_26_port, QN 
                           => n169);
   c_state_bpw_reg_27_inst : DFFR_X1 port map( D => n_state_bpw_27_port, CK => 
                           clk, RN => n306_port, Q => c_state_bpw_27_port, QN 
                           => n168);
   c_state_bpw_reg_28_inst : DFFR_X1 port map( D => n_state_bpw_28_port, CK => 
                           clk, RN => n306_port, Q => c_state_bpw_28_port, QN 
                           => n167);
   c_state_bpw_reg_29_inst : DFFR_X1 port map( D => n_state_bpw_29_port, CK => 
                           clk, RN => n306_port, Q => c_state_bpw_29_port, QN 
                           => n166);
   c_state_bpw_reg_30_inst : DFFR_X1 port map( D => n_state_bpw_30_port, CK => 
                           clk, RN => n306_port, Q => c_state_bpw_30_port, QN 
                           => n165);
   c_state_bpw_reg_31_inst : DFFR_X1 port map( D => n_state_bpw_31_port, CK => 
                           clk, RN => n306_port, Q => c_state_bpw_31_port, QN 
                           => n164);
   c_state_mul_reg_0_inst : DFFR_X1 port map( D => n_state_mul_0_port, CK => 
                           clk, RN => n320, Q => c_state_mul_0_port, QN => 
                           n294_port);
   c_state_mul_reg_10_inst : DFFR_X1 port map( D => n_state_mul_10_port, CK => 
                           clk, RN => n318, Q => c_state_mul_10_port, QN => 
                           net163738);
   c_state_mul_reg_1_inst : DFFR_X1 port map( D => n_state_mul_1_port, CK => 
                           clk, RN => n320, Q => c_state_mul_1_port, QN => n163
                           );
   c_state_mul_reg_2_inst : DFFR_X1 port map( D => n_state_mul_2_port, CK => 
                           clk, RN => n320, Q => c_state_mul_2_port, QN => n310
                           );
   c_state_mul_reg_3_inst : DFFR_X1 port map( D => n_state_mul_3_port, CK => 
                           clk, RN => n320, Q => c_state_mul_3_port, QN => 
                           n222_port);
   c_state_mul_reg_4_inst : DFFR_X1 port map( D => n_state_mul_4_port, CK => 
                           clk, RN => n320, Q => c_state_mul_4_port, QN => 
                           net108045);
   c_state_mul_reg_5_inst : DFFR_X1 port map( D => n_state_mul_5_port, CK => 
                           clk, RN => n320, Q => c_state_mul_5_port, QN => 
                           net108044);
   c_state_mul_reg_6_inst : DFFR_X1 port map( D => n_state_mul_6_port, CK => 
                           clk, RN => n320, Q => c_state_mul_6_port, QN => 
                           net108043);
   c_state_mul_reg_7_inst : DFFR_X1 port map( D => n_state_mul_7_port, CK => 
                           clk, RN => n320, Q => c_state_mul_7_port, QN => 
                           net163737);
   c_state_mul_reg_8_inst : DFFR_X1 port map( D => n_state_mul_8_port, CK => 
                           clk, RN => n319, Q => c_state_mul_8_port, QN => 
                           net163736);
   c_state_mul_reg_9_inst : DFFR_X1 port map( D => n_state_mul_9_port, CK => 
                           clk, RN => n319, Q => c_state_mul_9_port, QN => 
                           net163735);
   c_state_mul_reg_11_inst : DFFR_X1 port map( D => n_state_mul_11_port, CK => 
                           clk, RN => n318, Q => c_state_mul_11_port, QN => 
                           net108042);
   c_state_mul_reg_12_inst : DFFR_X1 port map( D => n_state_mul_12_port, CK => 
                           clk, RN => n318, Q => c_state_mul_12_port, QN => 
                           net108041);
   c_state_mul_reg_13_inst : DFFR_X1 port map( D => n_state_mul_13_port, CK => 
                           clk, RN => n318, Q => c_state_mul_13_port, QN => 
                           net108040);
   c_state_mul_reg_14_inst : DFFR_X1 port map( D => n_state_mul_14_port, CK => 
                           clk, RN => n318, Q => c_state_mul_14_port, QN => 
                           net163734);
   c_state_mul_reg_15_inst : DFFR_X1 port map( D => n_state_mul_15_port, CK => 
                           clk, RN => n318, Q => c_state_mul_15_port, QN => 
                           net163733);
   c_state_mul_reg_16_inst : DFFR_X1 port map( D => n_state_mul_16_port, CK => 
                           clk, RN => n318, Q => c_state_mul_16_port, QN => 
                           n160);
   c_state_mul_reg_17_inst : DFFR_X1 port map( D => n_state_mul_17_port, CK => 
                           clk, RN => n318, Q => c_state_mul_17_port, QN => 
                           net108039);
   c_state_mul_reg_18_inst : DFFR_X1 port map( D => n_state_mul_18_port, CK => 
                           clk, RN => n318, Q => c_state_mul_18_port, QN => 
                           net108038);
   c_state_mul_reg_19_inst : DFFR_X1 port map( D => n_state_mul_19_port, CK => 
                           clk, RN => n318, Q => c_state_mul_19_port, QN => 
                           net108037);
   c_state_mul_reg_20_inst : DFFR_X1 port map( D => n_state_mul_20_port, CK => 
                           clk, RN => n318, Q => c_state_mul_20_port, QN => 
                           n159);
   c_state_mul_reg_21_inst : DFFR_X1 port map( D => n_state_mul_21_port, CK => 
                           clk, RN => n318, Q => c_state_mul_21_port, QN => 
                           n158);
   c_state_mul_reg_22_inst : DFFR_X1 port map( D => n_state_mul_22_port, CK => 
                           clk, RN => n319, Q => c_state_mul_22_port, QN => 
                           n157);
   c_state_mul_reg_23_inst : DFFR_X1 port map( D => n_state_mul_23_port, CK => 
                           clk, RN => n319, Q => c_state_mul_23_port, QN => 
                           net163732);
   c_state_mul_reg_24_inst : DFFR_X1 port map( D => n_state_mul_24_port, CK => 
                           clk, RN => n319, Q => c_state_mul_24_port, QN => 
                           net108036);
   c_state_mul_reg_25_inst : DFFR_X1 port map( D => n_state_mul_25_port, CK => 
                           clk, RN => n319, Q => c_state_mul_25_port, QN => 
                           net108035);
   c_state_mul_reg_26_inst : DFFR_X1 port map( D => n_state_mul_26_port, CK => 
                           clk, RN => n319, Q => c_state_mul_26_port, QN => 
                           net108034);
   c_state_mul_reg_27_inst : DFFR_X1 port map( D => n_state_mul_27_port, CK => 
                           clk, RN => n319, Q => c_state_mul_27_port, QN => 
                           n307_port);
   c_state_mul_reg_28_inst : DFFR_X1 port map( D => n_state_mul_28_port, CK => 
                           clk, RN => n319, Q => c_state_mul_28_port, QN => 
                           n308_port);
   c_state_mul_reg_29_inst : DFFR_X1 port map( D => n_state_mul_29_port, CK => 
                           clk, RN => n319, Q => c_state_mul_29_port, QN => 
                           n309_port);
   c_state_mul_reg_30_inst : DFFR_X1 port map( D => n_state_mul_30_port, CK => 
                           clk, RN => n319, Q => c_state_mul_30_port, QN => 
                           n311);
   c_state_mul_reg_31_inst : DFFR_X1 port map( D => n_state_mul_31_port, CK => 
                           clk, RN => n319, Q => c_state_mul_31_port, QN => 
                           n312);
   c_state_div_reg_0_inst : DFFR_X1 port map( D => n_state_div_0_port, CK => 
                           clk, RN => n323, Q => c_state_div_0_port, QN => 
                           net163731);
   c_state_div_reg_10_inst : DFFR_X1 port map( D => n_state_div_10_port, CK => 
                           clk, RN => n320, Q => c_state_div_10_port, QN => 
                           net163730);
   c_state_div_reg_1_inst : DFFR_X1 port map( D => n_state_div_1_port, CK => 
                           clk, RN => n323, Q => c_state_div_1_port, QN => n155
                           );
   c_state_div_reg_2_inst : DFFR_X1 port map( D => n_state_div_2_port, CK => 
                           clk, RN => n323, Q => c_state_div_2_port, QN => n344
                           );
   c_state_div_reg_3_inst : DFFR_X1 port map( D => n_state_div_3_port, CK => 
                           clk, RN => n323, Q => c_state_div_3_port, QN => n347
                           );
   c_state_div_reg_4_inst : DFFR_X1 port map( D => n_state_div_4_port, CK => 
                           clk, RN => n322, Q => c_state_div_4_port, QN => n348
                           );
   c_state_div_reg_5_inst : DFFR_X1 port map( D => n_state_div_5_port, CK => 
                           clk, RN => n322, Q => c_state_div_5_port, QN => n230
                           );
   c_state_div_reg_6_inst : DFFR_X1 port map( D => n_state_div_6_port, CK => 
                           clk, RN => n322, Q => c_state_div_6_port, QN => 
                           net108033);
   c_state_div_reg_7_inst : DFFR_X1 port map( D => n_state_div_7_port, CK => 
                           clk, RN => n322, Q => c_state_div_7_port, QN => 
                           net108032);
   c_state_div_reg_8_inst : DFFR_X1 port map( D => n_state_div_8_port, CK => 
                           clk, RN => n322, Q => c_state_div_8_port, QN => 
                           net108031);
   c_state_div_reg_9_inst : DFFR_X1 port map( D => n_state_div_9_port, CK => 
                           clk, RN => n322, Q => c_state_div_9_port, QN => 
                           net163729);
   c_state_div_reg_11_inst : DFFR_X1 port map( D => n_state_div_11_port, CK => 
                           clk, RN => n320, Q => c_state_div_11_port, QN => 
                           net108030);
   c_state_div_reg_12_inst : DFFR_X1 port map( D => n_state_div_12_port, CK => 
                           clk, RN => n320, Q => c_state_div_12_port, QN => 
                           net108029);
   c_state_div_reg_13_inst : DFFR_X1 port map( D => n_state_div_13_port, CK => 
                           clk, RN => n320, Q => c_state_div_13_port, QN => 
                           n249);
   c_state_div_reg_14_inst : DFFR_X1 port map( D => n_state_div_14_port, CK => 
                           clk, RN => n321, Q => c_state_div_14_port, QN => 
                           net163728);
   c_state_div_reg_15_inst : DFFR_X1 port map( D => n_state_div_15_port, CK => 
                           clk, RN => n321, Q => c_state_div_15_port, QN => 
                           net163727);
   c_state_div_reg_16_inst : DFFR_X1 port map( D => n_state_div_16_port, CK => 
                           clk, RN => n321, Q => c_state_div_16_port, QN => 
                           net108028);
   c_state_div_reg_17_inst : DFFR_X1 port map( D => n_state_div_17_port, CK => 
                           clk, RN => n321, Q => c_state_div_17_port, QN => 
                           net108027);
   c_state_div_reg_18_inst : DFFR_X1 port map( D => n_state_div_18_port, CK => 
                           clk, RN => n321, Q => c_state_div_18_port, QN => 
                           net108026);
   c_state_div_reg_19_inst : DFFR_X1 port map( D => n_state_div_19_port, CK => 
                           clk, RN => n321, Q => c_state_div_19_port, QN => 
                           net163726);
   c_state_div_reg_20_inst : DFFR_X1 port map( D => n_state_div_20_port, CK => 
                           clk, RN => n321, Q => c_state_div_20_port, QN => 
                           n244);
   c_state_div_reg_21_inst : DFFR_X1 port map( D => n_state_div_21_port, CK => 
                           clk, RN => n321, Q => c_state_div_21_port, QN => 
                           n243);
   c_state_div_reg_22_inst : DFFR_X1 port map( D => n_state_div_22_port, CK => 
                           clk, RN => n321, Q => c_state_div_22_port, QN => 
                           net108025);
   c_state_div_reg_23_inst : DFFR_X1 port map( D => n_state_div_23_port, CK => 
                           clk, RN => n321, Q => c_state_div_23_port, QN => 
                           net108024);
   c_state_div_reg_24_inst : DFFR_X1 port map( D => n_state_div_24_port, CK => 
                           clk, RN => n321, Q => c_state_div_24_port, QN => 
                           net108023);
   c_state_div_reg_25_inst : DFFR_X1 port map( D => n_state_div_25_port, CK => 
                           clk, RN => n321, Q => c_state_div_25_port, QN => 
                           n242);
   c_state_div_reg_26_inst : DFFR_X1 port map( D => n_state_div_26_port, CK => 
                           clk, RN => n322, Q => c_state_div_26_port, QN => 
                           n241);
   c_state_div_reg_27_inst : DFFR_X1 port map( D => n_state_div_27_port, CK => 
                           clk, RN => n322, Q => c_state_div_27_port, QN => 
                           net108022);
   c_state_div_reg_28_inst : DFFR_X1 port map( D => n_state_div_28_port, CK => 
                           clk, RN => n322, Q => c_state_div_28_port, QN => 
                           n342);
   c_state_div_reg_29_inst : DFFR_X1 port map( D => n_state_div_29_port, CK => 
                           clk, RN => n322, Q => c_state_div_29_port, QN => 
                           n343);
   c_state_div_reg_30_inst : DFFR_X1 port map( D => n_state_div_30_port, CK => 
                           clk, RN => n322, Q => c_state_div_30_port, QN => 
                           net163725);
   c_state_div_reg_31_inst : DFFR_X1 port map( D => n_state_div_31_port, CK => 
                           clk, RN => n322, Q => c_state_div_31_port, QN => 
                           net108021);
   c_state_sqrt_reg_0_inst : DFFR_X1 port map( D => n_state_sqrt_0_port, CK => 
                           clk, RN => n315, Q => c_state_sqrt_0_port, QN => 
                           n247);
   c_state_sqrt_reg_10_inst : DFFR_X1 port map( D => n_state_sqrt_10_port, CK 
                           => clk, RN => n306_port, Q => c_state_sqrt_10_port, 
                           QN => n276);
   c_state_sqrt_reg_1_inst : DFFR_X1 port map( D => n_state_sqrt_1_port, CK => 
                           clk, RN => n315, Q => c_state_sqrt_1_port, QN => 
                           n240);
   c_state_sqrt_reg_2_inst : DFFR_X1 port map( D => n_state_sqrt_2_port, CK => 
                           clk, RN => n315, Q => c_state_sqrt_2_port, QN => 
                           n263);
   c_state_sqrt_reg_3_inst : DFFR_X1 port map( D => n_state_sqrt_3_port, CK => 
                           clk, RN => n315, Q => c_state_sqrt_3_port, QN => 
                           n266);
   c_state_sqrt_reg_4_inst : DFFR_X1 port map( D => n_state_sqrt_4_port, CK => 
                           clk, RN => n314, Q => c_state_sqrt_4_port, QN => 
                           net108020);
   c_state_sqrt_reg_5_inst : DFFR_X1 port map( D => n_state_sqrt_5_port, CK => 
                           clk, RN => n314, Q => c_state_sqrt_5_port, QN => 
                           net163724);
   c_state_sqrt_reg_6_inst : DFFR_X1 port map( D => n_state_sqrt_6_port, CK => 
                           clk, RN => n314, Q => c_state_sqrt_6_port, QN => 
                           net108019);
   c_state_sqrt_reg_7_inst : DFFR_X1 port map( D => n_state_sqrt_7_port, CK => 
                           clk, RN => n314, Q => c_state_sqrt_7_port, QN => 
                           net108018);
   c_state_sqrt_reg_8_inst : DFFR_X1 port map( D => n_state_sqrt_8_port, CK => 
                           clk, RN => n314, Q => c_state_sqrt_8_port, QN => 
                           net108017);
   c_state_sqrt_reg_9_inst : DFFR_X1 port map( D => n_state_sqrt_9_port, CK => 
                           clk, RN => n314, Q => c_state_sqrt_9_port, QN => 
                           net163723);
   c_state_sqrt_reg_11_inst : DFFR_X1 port map( D => n_state_sqrt_11_port, CK 
                           => clk, RN => n306_port, Q => c_state_sqrt_11_port, 
                           QN => net108016);
   c_state_sqrt_reg_12_inst : DFFR_X1 port map( D => n_state_sqrt_12_port, CK 
                           => clk, RN => n306_port, Q => c_state_sqrt_12_port, 
                           QN => net108015);
   c_state_sqrt_reg_13_inst : DFFR_X1 port map( D => n_state_sqrt_13_port, CK 
                           => clk, RN => n306_port, Q => c_state_sqrt_13_port, 
                           QN => n239);
   c_state_sqrt_reg_14_inst : DFFR_X1 port map( D => n_state_sqrt_14_port, CK 
                           => clk, RN => n313, Q => c_state_sqrt_14_port, QN =>
                           net163722);
   c_state_sqrt_reg_15_inst : DFFR_X1 port map( D => n_state_sqrt_15_port, CK 
                           => clk, RN => n313, Q => c_state_sqrt_15_port, QN =>
                           net163721);
   c_state_sqrt_reg_16_inst : DFFR_X1 port map( D => n_state_sqrt_16_port, CK 
                           => clk, RN => n313, Q => c_state_sqrt_16_port, QN =>
                           net108014);
   c_state_sqrt_reg_17_inst : DFFR_X1 port map( D => n_state_sqrt_17_port, CK 
                           => clk, RN => n313, Q => c_state_sqrt_17_port, QN =>
                           net108013);
   c_state_sqrt_reg_18_inst : DFFR_X1 port map( D => n_state_sqrt_18_port, CK 
                           => clk, RN => n313, Q => c_state_sqrt_18_port, QN =>
                           net108012);
   c_state_sqrt_reg_19_inst : DFFR_X1 port map( D => n_state_sqrt_19_port, CK 
                           => clk, RN => n313, Q => c_state_sqrt_19_port, QN =>
                           net163720);
   c_state_sqrt_reg_20_inst : DFFR_X1 port map( D => n_state_sqrt_20_port, CK 
                           => clk, RN => n313, Q => c_state_sqrt_20_port, QN =>
                           n235);
   c_state_sqrt_reg_21_inst : DFFR_X1 port map( D => n_state_sqrt_21_port, CK 
                           => clk, RN => n313, Q => c_state_sqrt_21_port, QN =>
                           n234);
   c_state_sqrt_reg_22_inst : DFFR_X1 port map( D => n_state_sqrt_22_port, CK 
                           => clk, RN => n313, Q => c_state_sqrt_22_port, QN =>
                           net108011);
   c_state_sqrt_reg_23_inst : DFFR_X1 port map( D => n_state_sqrt_23_port, CK 
                           => clk, RN => n313, Q => c_state_sqrt_23_port, QN =>
                           net108010);
   c_state_sqrt_reg_24_inst : DFFR_X1 port map( D => n_state_sqrt_24_port, CK 
                           => clk, RN => n313, Q => c_state_sqrt_24_port, QN =>
                           net108009);
   c_state_sqrt_reg_25_inst : DFFR_X1 port map( D => n_state_sqrt_25_port, CK 
                           => clk, RN => n313, Q => c_state_sqrt_25_port, QN =>
                           n233);
   c_state_sqrt_reg_26_inst : DFFR_X1 port map( D => n_state_sqrt_26_port, CK 
                           => clk, RN => n314, Q => c_state_sqrt_26_port, QN =>
                           n229);
   c_state_sqrt_reg_27_inst : DFFR_X1 port map( D => n_state_sqrt_27_port, CK 
                           => clk, RN => n314, Q => c_state_sqrt_27_port, QN =>
                           net108008);
   c_state_sqrt_reg_28_inst : DFFR_X1 port map( D => n_state_sqrt_28_port, CK 
                           => clk, RN => n314, Q => c_state_sqrt_28_port, QN =>
                           n261);
   c_state_sqrt_reg_29_inst : DFFR_X1 port map( D => n_state_sqrt_29_port, CK 
                           => clk, RN => n314, Q => c_state_sqrt_29_port, QN =>
                           n262);
   c_state_sqrt_reg_30_inst : DFFR_X1 port map( D => n_state_sqrt_30_port, CK 
                           => clk, RN => n314, Q => c_state_sqrt_30_port, QN =>
                           net163719);
   c_state_sqrt_reg_31_inst : DFFR_X1 port map( D => n_state_sqrt_31_port, CK 
                           => clk, RN => n314, Q => c_state_sqrt_31_port, QN =>
                           net108007);
   c_state_stu_reg_0_inst : DFFR_X1 port map( D => n_state_stu_0_port, CK => 
                           clk, RN => n325, Q => c_state_stu_0_port, QN => n192
                           );
   c_state_stu_reg_31_inst : DFFR_X1 port map( D => n_state_stu_31_port, CK => 
                           clk, RN => n325, Q => c_state_stu_31_port, QN => 
                           n228);
   c_state_stu_reg_2_inst : DFFR_X1 port map( D => n_state_stu_2_port, CK => 
                           clk, RN => n325, Q => c_state_stu_2_port, QN => 
                           n214_port);
   c_state_stu_reg_9_inst : DFFR_X1 port map( D => n_state_stu_9_port, CK => 
                           clk, RN => n325, Q => c_state_stu_9_port, QN => 
                           net108006);
   c_state_stu_reg_8_inst : DFFR_X1 port map( D => n_state_stu_8_port, CK => 
                           clk, RN => n325, Q => c_state_stu_8_port, QN => 
                           net108005);
   c_state_stu_reg_7_inst : DFFR_X1 port map( D => n_state_stu_7_port, CK => 
                           clk, RN => n325, Q => c_state_stu_7_port, QN => 
                           net108004);
   c_state_stu_reg_6_inst : DFFR_X1 port map( D => n_state_stu_6_port, CK => 
                           clk, RN => n325, Q => c_state_stu_6_port, QN => n227
                           );
   c_state_stu_reg_5_inst : DFFR_X1 port map( D => n_state_stu_5_port, CK => 
                           clk, RN => n325, Q => c_state_stu_5_port, QN => n226
                           );
   c_state_stu_reg_4_inst : DFFR_X1 port map( D => n_state_stu_4_port, CK => 
                           clk, RN => n325, Q => c_state_stu_4_port, QN => 
                           net163718);
   c_state_stu_reg_3_inst : DFFR_X1 port map( D => n_state_stu_3_port, CK => 
                           clk, RN => n325, Q => c_state_stu_3_port, QN => 
                           net163717);
   c_state_stu_reg_30_inst : DFFR_X1 port map( D => n_state_stu_30_port, CK => 
                           clk, RN => n325, Q => c_state_stu_30_port, QN => 
                           net108003);
   c_state_stu_reg_29_inst : DFFR_X1 port map( D => n_state_stu_29_port, CK => 
                           clk, RN => n324, Q => c_state_stu_29_port, QN => 
                           net108002);
   c_state_stu_reg_28_inst : DFFR_X1 port map( D => n_state_stu_28_port, CK => 
                           clk, RN => n324, Q => c_state_stu_28_port, QN => 
                           net108001);
   c_state_stu_reg_27_inst : DFFR_X1 port map( D => n_state_stu_27_port, CK => 
                           clk, RN => n324, Q => c_state_stu_27_port, QN => 
                           net163716);
   c_state_stu_reg_26_inst : DFFR_X1 port map( D => n_state_stu_26_port, CK => 
                           clk, RN => n324, Q => c_state_stu_26_port, QN => 
                           n221_port);
   c_state_stu_reg_25_inst : DFFR_X1 port map( D => n_state_stu_25_port, CK => 
                           clk, RN => n324, Q => c_state_stu_25_port, QN => 
                           n220_port);
   c_state_stu_reg_24_inst : DFFR_X1 port map( D => n_state_stu_24_port, CK => 
                           clk, RN => n324, Q => c_state_stu_24_port, QN => 
                           n219_port);
   c_state_stu_reg_23_inst : DFFR_X1 port map( D => n_state_stu_23_port, CK => 
                           clk, RN => n324, Q => c_state_stu_23_port, QN => 
                           net108000);
   c_state_stu_reg_22_inst : DFFR_X1 port map( D => n_state_stu_22_port, CK => 
                           clk, RN => n324, Q => c_state_stu_22_port, QN => 
                           net107999);
   c_state_stu_reg_21_inst : DFFR_X1 port map( D => n_state_stu_21_port, CK => 
                           clk, RN => n324, Q => c_state_stu_21_port, QN => 
                           net107998);
   c_state_stu_reg_20_inst : DFFR_X1 port map( D => n_state_stu_20_port, CK => 
                           clk, RN => n324, Q => c_state_stu_20_port, QN => 
                           n218_port);
   c_state_stu_reg_1_inst : DFFR_X1 port map( D => n_state_stu_1_port, CK => 
                           clk, RN => n325, Q => c_state_stu_1_port, QN => 
                           n194_port);
   c_state_stu_reg_19_inst : DFFR_X1 port map( D => n_state_stu_19_port, CK => 
                           clk, RN => n324, Q => c_state_stu_19_port, QN => 
                           net163715);
   c_state_stu_reg_18_inst : DFFR_X1 port map( D => n_state_stu_18_port, CK => 
                           clk, RN => n324, Q => c_state_stu_18_port, QN => 
                           net163714);
   c_state_stu_reg_17_inst : DFFR_X1 port map( D => n_state_stu_17_port, CK => 
                           clk, RN => n323, Q => c_state_stu_17_port, QN => 
                           net163713);
   c_state_stu_reg_16_inst : DFFR_X1 port map( D => n_state_stu_16_port, CK => 
                           clk, RN => n323, Q => c_state_stu_16_port, QN => 
                           net107997);
   c_state_stu_reg_15_inst : DFFR_X1 port map( D => n_state_stu_15_port, CK => 
                           clk, RN => n323, Q => c_state_stu_15_port, QN => 
                           net107996);
   c_state_stu_reg_14_inst : DFFR_X1 port map( D => n_state_stu_14_port, CK => 
                           clk, RN => n323, Q => c_state_stu_14_port, QN => 
                           net107995);
   c_state_stu_reg_13_inst : DFFR_X1 port map( D => n_state_stu_13_port, CK => 
                           clk, RN => n323, Q => c_state_stu_13_port, QN => 
                           n213_port);
   c_state_stu_reg_12_inst : DFFR_X1 port map( D => n_state_stu_12_port, CK => 
                           clk, RN => n323, Q => c_state_stu_12_port, QN => 
                           n212_port);
   c_state_stu_reg_11_inst : DFFR_X1 port map( D => n_state_stu_11_port, CK => 
                           clk, RN => n323, Q => c_state_stu_11_port, QN => 
                           n211_port);
   c_state_stu_reg_10_inst : DFFR_X1 port map( D => n_state_stu_10_port, CK => 
                           clk, RN => n323, Q => c_state_stu_10_port, QN => 
                           n210_port);
   U333 : NAND3_X1 port map( A1 => n39, A2 => n300_port, A3 => n38, ZN => 
                           stall_flag_2_port);
   U334 : NAND3_X1 port map( A1 => n44, A2 => n45, A3 => n46_port, ZN => n43);
   U335 : NAND3_X1 port map( A1 => n78, A2 => n79, A3 => n80, ZN => 
                           stall_flag_0_port);
   U336 : NAND3_X1 port map( A1 => n214_port, A2 => n86, A3 => n228, ZN => 
                           n75_port);
   U337 : NAND3_X1 port map( A1 => n88, A2 => n312, A3 => n89, ZN => n66_port);
   U338 : OAI33_X1 port map( A1 => c_state_sqrt_0_port, A2 => net108020, A3 => 
                           n69_port, B1 => c_state_sqrt_4_port, B2 => n100, B3 
                           => n101, ZN => n68_port);
   U339 : OAI33_X1 port map( A1 => n102, A2 => n230, A3 => c_state_div_0_port, 
                           B1 => c_state_div_5_port, B2 => n103, B3 => n104, ZN
                           => n62_port);
   U340 : NAND3_X1 port map( A1 => n261, A2 => n239, A3 => n262, ZN => 
                           n129_port);
   U341 : NAND3_X1 port map( A1 => net108015, A2 => net108014, A3 => net108016,
                           ZN => n131_port);
   U342 : NAND3_X1 port map( A1 => n133_port, A2 => n96, A3 => N46, ZN => 
                           n134_port);
   U343 : NAND3_X1 port map( A1 => n185, A2 => n76_port, A3 => n195_port, ZN =>
                           n96);
   U344 : NAND3_X1 port map( A1 => net108035, A2 => net108034, A3 => net108036,
                           ZN => n254);
   U345 : NAND3_X1 port map( A1 => n342, A2 => n249, A3 => n343, ZN => n274);
   U346 : NAND3_X1 port map( A1 => net108023, A2 => net108022, A3 => net108024,
                           ZN => n275);
   U347 : NAND3_X1 port map( A1 => net108029, A2 => net108028, A3 => net108030,
                           ZN => n277);
   U348 : NAND3_X1 port map( A1 => n279_port, A2 => n85, A3 => N119, ZN => 
                           n280_port);
   U349 : NAND3_X1 port map( A1 => n164, A2 => n281_port, A3 => n197_port, ZN 
                           => n85);
   add_319 : StallGenerator_CWRD_SIZE20_DW01_inc_0 port map( A(31) => 
                           c_state_stu_31_port, A(30) => c_state_stu_30_port, 
                           A(29) => c_state_stu_29_port, A(28) => 
                           c_state_stu_28_port, A(27) => c_state_stu_27_port, 
                           A(26) => c_state_stu_26_port, A(25) => 
                           c_state_stu_25_port, A(24) => c_state_stu_24_port, 
                           A(23) => c_state_stu_23_port, A(22) => 
                           c_state_stu_22_port, A(21) => c_state_stu_21_port, 
                           A(20) => c_state_stu_20_port, A(19) => 
                           c_state_stu_19_port, A(18) => c_state_stu_18_port, 
                           A(17) => c_state_stu_17_port, A(16) => 
                           c_state_stu_16_port, A(15) => c_state_stu_15_port, 
                           A(14) => c_state_stu_14_port, A(13) => 
                           c_state_stu_13_port, A(12) => c_state_stu_12_port, 
                           A(11) => c_state_stu_11_port, A(10) => 
                           c_state_stu_10_port, A(9) => c_state_stu_9_port, 
                           A(8) => c_state_stu_8_port, A(7) => 
                           c_state_stu_7_port, A(6) => c_state_stu_6_port, A(5)
                           => c_state_stu_5_port, A(4) => c_state_stu_4_port, 
                           A(3) => c_state_stu_3_port, A(2) => 
                           c_state_stu_2_port, A(1) => c_state_stu_1_port, A(0)
                           => c_state_stu_0_port, SUM(31) => N475, SUM(30) => 
                           N474, SUM(29) => N473, SUM(28) => N472, SUM(27) => 
                           N471, SUM(26) => N470, SUM(25) => N469, SUM(24) => 
                           N468, SUM(23) => N467, SUM(22) => N466, SUM(21) => 
                           N465, SUM(20) => N464, SUM(19) => N463, SUM(18) => 
                           N462, SUM(17) => N461, SUM(16) => N460, SUM(15) => 
                           N459, SUM(14) => N458, SUM(13) => N457, SUM(12) => 
                           N456, SUM(11) => N455, SUM(10) => N454, SUM(9) => 
                           N453, SUM(8) => N452, SUM(7) => N451, SUM(6) => N450
                           , SUM(5) => N449, SUM(4) => N448, SUM(3) => N447, 
                           SUM(2) => N446, SUM(1) => N445, SUM(0) => N444);
   add_277 : StallGenerator_CWRD_SIZE20_DW01_inc_1 port map( A(31) => 
                           c_state_sqrt_31_port, A(30) => c_state_sqrt_30_port,
                           A(29) => c_state_sqrt_29_port, A(28) => 
                           c_state_sqrt_28_port, A(27) => c_state_sqrt_27_port,
                           A(26) => c_state_sqrt_26_port, A(25) => 
                           c_state_sqrt_25_port, A(24) => c_state_sqrt_24_port,
                           A(23) => c_state_sqrt_23_port, A(22) => 
                           c_state_sqrt_22_port, A(21) => c_state_sqrt_21_port,
                           A(20) => c_state_sqrt_20_port, A(19) => 
                           c_state_sqrt_19_port, A(18) => c_state_sqrt_18_port,
                           A(17) => c_state_sqrt_17_port, A(16) => 
                           c_state_sqrt_16_port, A(15) => c_state_sqrt_15_port,
                           A(14) => c_state_sqrt_14_port, A(13) => 
                           c_state_sqrt_13_port, A(12) => c_state_sqrt_12_port,
                           A(11) => c_state_sqrt_11_port, A(10) => 
                           c_state_sqrt_10_port, A(9) => c_state_sqrt_9_port, 
                           A(8) => c_state_sqrt_8_port, A(7) => 
                           c_state_sqrt_7_port, A(6) => c_state_sqrt_6_port, 
                           A(5) => c_state_sqrt_5_port, A(4) => 
                           c_state_sqrt_4_port, A(3) => c_state_sqrt_3_port, 
                           A(2) => c_state_sqrt_2_port, A(1) => 
                           c_state_sqrt_1_port, A(0) => c_state_sqrt_0_port, 
                           SUM(31) => N394, SUM(30) => N393, SUM(29) => N392, 
                           SUM(28) => N391, SUM(27) => N390, SUM(26) => N389, 
                           SUM(25) => N388, SUM(24) => N387, SUM(23) => N386, 
                           SUM(22) => N385, SUM(21) => N384, SUM(20) => N383, 
                           SUM(19) => N382, SUM(18) => N381, SUM(17) => N380, 
                           SUM(16) => N379, SUM(15) => N378, SUM(14) => N377, 
                           SUM(13) => N376, SUM(12) => N375, SUM(11) => N374, 
                           SUM(10) => N373, SUM(9) => N372, SUM(8) => N371, 
                           SUM(7) => N370, SUM(6) => N369, SUM(5) => N368, 
                           SUM(4) => N367, SUM(3) => N366, SUM(2) => N365, 
                           SUM(1) => N364, SUM(0) => N363);
   add_232 : StallGenerator_CWRD_SIZE20_DW01_inc_2 port map( A(31) => 
                           c_state_div_31_port, A(30) => c_state_div_30_port, 
                           A(29) => c_state_div_29_port, A(28) => 
                           c_state_div_28_port, A(27) => c_state_div_27_port, 
                           A(26) => c_state_div_26_port, A(25) => 
                           c_state_div_25_port, A(24) => c_state_div_24_port, 
                           A(23) => c_state_div_23_port, A(22) => 
                           c_state_div_22_port, A(21) => c_state_div_21_port, 
                           A(20) => c_state_div_20_port, A(19) => 
                           c_state_div_19_port, A(18) => c_state_div_18_port, 
                           A(17) => c_state_div_17_port, A(16) => 
                           c_state_div_16_port, A(15) => c_state_div_15_port, 
                           A(14) => c_state_div_14_port, A(13) => 
                           c_state_div_13_port, A(12) => c_state_div_12_port, 
                           A(11) => c_state_div_11_port, A(10) => 
                           c_state_div_10_port, A(9) => c_state_div_9_port, 
                           A(8) => c_state_div_8_port, A(7) => 
                           c_state_div_7_port, A(6) => c_state_div_6_port, A(5)
                           => c_state_div_5_port, A(4) => c_state_div_4_port, 
                           A(3) => c_state_div_3_port, A(2) => 
                           c_state_div_2_port, A(1) => c_state_div_1_port, A(0)
                           => c_state_div_0_port, SUM(31) => N309, SUM(30) => 
                           N308, SUM(29) => N307, SUM(28) => N306, SUM(27) => 
                           N305, SUM(26) => N304, SUM(25) => N303, SUM(24) => 
                           N302, SUM(23) => N301, SUM(22) => N300, SUM(21) => 
                           N299, SUM(20) => N298, SUM(19) => N297, SUM(18) => 
                           N296, SUM(17) => N295, SUM(16) => N294, SUM(15) => 
                           N293, SUM(14) => N292, SUM(13) => N291, SUM(12) => 
                           N290, SUM(11) => N289, SUM(10) => N288, SUM(9) => 
                           N287, SUM(8) => N286, SUM(7) => N285, SUM(6) => N284
                           , SUM(5) => N283, SUM(4) => N282, SUM(3) => N281, 
                           SUM(2) => N280, SUM(1) => N279, SUM(0) => N278);
   add_187 : StallGenerator_CWRD_SIZE20_DW01_inc_3 port map( A(31) => 
                           c_state_mul_31_port, A(30) => c_state_mul_30_port, 
                           A(29) => c_state_mul_29_port, A(28) => 
                           c_state_mul_28_port, A(27) => c_state_mul_27_port, 
                           A(26) => c_state_mul_26_port, A(25) => 
                           c_state_mul_25_port, A(24) => c_state_mul_24_port, 
                           A(23) => c_state_mul_23_port, A(22) => 
                           c_state_mul_22_port, A(21) => c_state_mul_21_port, 
                           A(20) => c_state_mul_20_port, A(19) => 
                           c_state_mul_19_port, A(18) => c_state_mul_18_port, 
                           A(17) => c_state_mul_17_port, A(16) => 
                           c_state_mul_16_port, A(15) => c_state_mul_15_port, 
                           A(14) => c_state_mul_14_port, A(13) => 
                           c_state_mul_13_port, A(12) => c_state_mul_12_port, 
                           A(11) => c_state_mul_11_port, A(10) => 
                           c_state_mul_10_port, A(9) => c_state_mul_9_port, 
                           A(8) => c_state_mul_8_port, A(7) => 
                           c_state_mul_7_port, A(6) => c_state_mul_6_port, A(5)
                           => c_state_mul_5_port, A(4) => c_state_mul_4_port, 
                           A(3) => c_state_mul_3_port, A(2) => 
                           c_state_mul_2_port, A(1) => c_state_mul_1_port, A(0)
                           => c_state_mul_0_port, SUM(31) => N224, SUM(30) => 
                           N223, SUM(29) => N222, SUM(28) => N221, SUM(27) => 
                           N220, SUM(26) => N219, SUM(25) => N218, SUM(24) => 
                           N217, SUM(23) => N216, SUM(22) => N215, SUM(21) => 
                           N214, SUM(20) => N213, SUM(19) => N212, SUM(18) => 
                           N211, SUM(17) => N210, SUM(16) => N209, SUM(15) => 
                           N208, SUM(14) => N207, SUM(13) => N206, SUM(12) => 
                           N205, SUM(11) => N204, SUM(10) => N203, SUM(9) => 
                           N202, SUM(8) => N201, SUM(7) => N200, SUM(6) => N199
                           , SUM(5) => N198, SUM(4) => N197, SUM(3) => N196, 
                           SUM(2) => N195, SUM(1) => N194, SUM(0) => N193);
   add_109 : StallGenerator_CWRD_SIZE20_DW01_inc_4 port map( A(31) => 
                           c_state_bpw_31_port, A(30) => c_state_bpw_30_port, 
                           A(29) => c_state_bpw_29_port, A(28) => 
                           c_state_bpw_28_port, A(27) => c_state_bpw_27_port, 
                           A(26) => c_state_bpw_26_port, A(25) => 
                           c_state_bpw_25_port, A(24) => c_state_bpw_24_port, 
                           A(23) => c_state_bpw_23_port, A(22) => 
                           c_state_bpw_22_port, A(21) => c_state_bpw_21_port, 
                           A(20) => c_state_bpw_20_port, A(19) => 
                           c_state_bpw_19_port, A(18) => c_state_bpw_18_port, 
                           A(17) => c_state_bpw_17_port, A(16) => 
                           c_state_bpw_16_port, A(15) => c_state_bpw_15_port, 
                           A(14) => c_state_bpw_14_port, A(13) => 
                           c_state_bpw_13_port, A(12) => c_state_bpw_12_port, 
                           A(11) => c_state_bpw_11_port, A(10) => 
                           c_state_bpw_10_port, A(9) => c_state_bpw_9_port, 
                           A(8) => c_state_bpw_8_port, A(7) => 
                           c_state_bpw_7_port, A(6) => c_state_bpw_6_port, A(5)
                           => c_state_bpw_5_port, A(4) => c_state_bpw_4_port, 
                           A(3) => c_state_bpw_3_port, A(2) => 
                           c_state_bpw_2_port, A(1) => c_state_bpw_1_port, A(0)
                           => c_state_bpw_0_port, SUM(31) => N150, SUM(30) => 
                           N149, SUM(29) => N148, SUM(28) => N147, SUM(27) => 
                           N146, SUM(26) => N145, SUM(25) => N144, SUM(24) => 
                           N143, SUM(23) => N142, SUM(22) => N141, SUM(21) => 
                           N140, SUM(20) => N139, SUM(19) => N138, SUM(18) => 
                           N137, SUM(17) => N136, SUM(16) => N135, SUM(15) => 
                           N134, SUM(14) => N133, SUM(13) => N132, SUM(12) => 
                           N131, SUM(11) => N130, SUM(10) => N129, SUM(9) => 
                           N128, SUM(8) => N127, SUM(7) => N126, SUM(6) => N125
                           , SUM(5) => N124, SUM(4) => N123, SUM(3) => N122, 
                           SUM(2) => N121, SUM(1) => N120, SUM(0) => N119);
   add_69 : StallGenerator_CWRD_SIZE20_DW01_inc_5 port map( A(31) => 
                           c_state_ral_31_port, A(30) => c_state_ral_30_port, 
                           A(29) => c_state_ral_29_port, A(28) => 
                           c_state_ral_28_port, A(27) => c_state_ral_27_port, 
                           A(26) => c_state_ral_26_port, A(25) => 
                           c_state_ral_25_port, A(24) => c_state_ral_24_port, 
                           A(23) => c_state_ral_23_port, A(22) => 
                           c_state_ral_22_port, A(21) => c_state_ral_21_port, 
                           A(20) => c_state_ral_20_port, A(19) => 
                           c_state_ral_19_port, A(18) => c_state_ral_18_port, 
                           A(17) => c_state_ral_17_port, A(16) => 
                           c_state_ral_16_port, A(15) => c_state_ral_15_port, 
                           A(14) => c_state_ral_14_port, A(13) => 
                           c_state_ral_13_port, A(12) => c_state_ral_12_port, 
                           A(11) => c_state_ral_11_port, A(10) => 
                           c_state_ral_10_port, A(9) => c_state_ral_9_port, 
                           A(8) => c_state_ral_8_port, A(7) => 
                           c_state_ral_7_port, A(6) => c_state_ral_6_port, A(5)
                           => c_state_ral_5_port, A(4) => c_state_ral_4_port, 
                           A(3) => c_state_ral_3_port, A(2) => 
                           c_state_ral_2_port, A(1) => c_state_ral_1_port, A(0)
                           => c_state_ral_0_port, SUM(31) => N77, SUM(30) => 
                           N76, SUM(29) => N75, SUM(28) => N74, SUM(27) => N73,
                           SUM(26) => N72, SUM(25) => N71, SUM(24) => N70, 
                           SUM(23) => N69, SUM(22) => N68, SUM(21) => N67, 
                           SUM(20) => N66, SUM(19) => N65, SUM(18) => N64, 
                           SUM(17) => N63, SUM(16) => N62, SUM(15) => N61, 
                           SUM(14) => N60, SUM(13) => N59, SUM(12) => N58, 
                           SUM(11) => N57, SUM(10) => N56, SUM(9) => N55, 
                           SUM(8) => N54, SUM(7) => N53, SUM(6) => N52, SUM(5) 
                           => N51, SUM(4) => N50, SUM(3) => N49, SUM(2) => N48,
                           SUM(1) => N47, SUM(0) => N46);
   U3 : AND3_X1 port map( A1 => n263, A2 => n240, A3 => n266, ZN => n100);
   U4 : NOR3_X1 port map( A1 => c_state_sqrt_0_port, A2 => n69_port, A3 => 
                           c_state_sqrt_4_port, ZN => n53_port);
   U5 : NOR3_X1 port map( A1 => n102, A2 => c_state_div_0_port, A3 => 
                           c_state_div_5_port, ZN => n60_port);
   U6 : NOR3_X1 port map( A1 => n65_port, A2 => c_state_mul_0_port, A3 => 
                           c_state_mul_3_port, ZN => n55_port);
   U7 : NOR2_X1 port map( A1 => n260, A2 => n104, ZN => n50_port);
   U8 : INV_X1 port map( A => n50_port, ZN => n102);
   U9 : INV_X1 port map( A => n69_port, ZN => n67_port);
   U10 : NOR3_X1 port map( A1 => n41, A2 => n42, A3 => n43, ZN => n38);
   U11 : OAI211_X1 port map( C1 => n83, C2 => n60_port, A => n45, B => sig_div,
                           ZN => n46_port);
   U12 : OAI211_X1 port map( C1 => n84, C2 => n55_port, A => n45, B => sig_mul,
                           ZN => n44);
   U13 : NAND2_X1 port map( A1 => n119_port, A2 => n100, ZN => n69_port);
   U14 : NAND2_X1 port map( A1 => n150_port, A2 => n151, ZN => n94);
   U15 : OAI21_X1 port map( B1 => c_state_mul_2_port, B2 => c_state_mul_1_port,
                           A => c_state_mul_3_port, ZN => n151);
   U16 : OAI21_X1 port map( B1 => c_state_mul_3_port, B2 => n65_port, A => 
                           n66_port, ZN => n63_port);
   U17 : INV_X1 port map( A => n118, ZN => n42);
   U18 : INV_X1 port map( A => n75_port, ZN => n70_port);
   U19 : INV_X1 port map( A => n260, ZN => n103);
   U20 : INV_X1 port map( A => n101, ZN => n119_port);
   U21 : AND2_X1 port map( A1 => N308, A2 => n291_port, ZN => 
                           n_state_div_30_port);
   U22 : AND2_X1 port map( A1 => N306, A2 => n291_port, ZN => 
                           n_state_div_28_port);
   U23 : AND2_X1 port map( A1 => N303, A2 => n291_port, ZN => 
                           n_state_div_25_port);
   U24 : AND2_X1 port map( A1 => N300, A2 => n291_port, ZN => 
                           n_state_div_22_port);
   U25 : AND2_X1 port map( A1 => N223, A2 => n293_port, ZN => 
                           n_state_mul_30_port);
   U26 : AND2_X1 port map( A1 => N221, A2 => n293_port, ZN => 
                           n_state_mul_28_port);
   U27 : AND2_X1 port map( A1 => N218, A2 => n293_port, ZN => 
                           n_state_mul_25_port);
   U28 : AND2_X1 port map( A1 => N215, A2 => n293_port, ZN => 
                           n_state_mul_22_port);
   U29 : AND2_X1 port map( A1 => N393, A2 => n297_port, ZN => 
                           n_state_sqrt_30_port);
   U30 : AND2_X1 port map( A1 => N391, A2 => n297_port, ZN => 
                           n_state_sqrt_28_port);
   U31 : AND2_X1 port map( A1 => N388, A2 => n297_port, ZN => 
                           n_state_sqrt_25_port);
   U32 : AND2_X1 port map( A1 => N385, A2 => n297_port, ZN => 
                           n_state_sqrt_22_port);
   U33 : AND2_X1 port map( A1 => N390, A2 => n296_port, ZN => 
                           n_state_sqrt_27_port);
   U34 : AND2_X1 port map( A1 => N387, A2 => n296_port, ZN => 
                           n_state_sqrt_24_port);
   U35 : AND2_X1 port map( A1 => N305, A2 => n271, ZN => n_state_div_27_port);
   U36 : AND2_X1 port map( A1 => N302, A2 => n271, ZN => n_state_div_24_port);
   U37 : AND2_X1 port map( A1 => N220, A2 => n292_port, ZN => 
                           n_state_mul_27_port);
   U38 : AND2_X1 port map( A1 => N217, A2 => n292_port, ZN => 
                           n_state_mul_24_port);
   U39 : AND2_X1 port map( A1 => N392, A2 => n116, ZN => n_state_sqrt_29_port);
   U40 : AND2_X1 port map( A1 => N389, A2 => n116, ZN => n_state_sqrt_26_port);
   U41 : AND2_X1 port map( A1 => N386, A2 => n116, ZN => n_state_sqrt_23_port);
   U42 : AND2_X1 port map( A1 => N307, A2 => n255, ZN => n_state_div_29_port);
   U43 : AND2_X1 port map( A1 => N304, A2 => n255, ZN => n_state_div_26_port);
   U44 : AND2_X1 port map( A1 => N301, A2 => n255, ZN => n_state_div_23_port);
   U45 : AND2_X1 port map( A1 => N222, A2 => n146_port, ZN => 
                           n_state_mul_29_port);
   U46 : AND2_X1 port map( A1 => N219, A2 => n146_port, ZN => 
                           n_state_mul_26_port);
   U47 : AND2_X1 port map( A1 => N216, A2 => n146_port, ZN => 
                           n_state_mul_23_port);
   U48 : AND2_X1 port map( A1 => N74, A2 => n132_port, ZN => 
                           n_state_ral_28_port);
   U49 : AND2_X1 port map( A1 => N72, A2 => n132_port, ZN => 
                           n_state_ral_26_port);
   U50 : AND2_X1 port map( A1 => N70, A2 => n132_port, ZN => 
                           n_state_ral_24_port);
   U51 : AND2_X1 port map( A1 => N68, A2 => n132_port, ZN => 
                           n_state_ral_22_port);
   U52 : AND2_X1 port map( A1 => N466, A2 => n105, ZN => n_state_stu_22_port);
   U53 : AND2_X1 port map( A1 => N467, A2 => n105, ZN => n_state_stu_23_port);
   U54 : AND2_X1 port map( A1 => N468, A2 => n105, ZN => n_state_stu_24_port);
   U55 : AND2_X1 port map( A1 => N469, A2 => n105, ZN => n_state_stu_25_port);
   U56 : AND2_X1 port map( A1 => N470, A2 => n105, ZN => n_state_stu_26_port);
   U57 : AND2_X1 port map( A1 => N471, A2 => n105, ZN => n_state_stu_27_port);
   U58 : AND2_X1 port map( A1 => N472, A2 => n105, ZN => n_state_stu_28_port);
   U59 : AND2_X1 port map( A1 => N473, A2 => n105, ZN => n_state_stu_29_port);
   U60 : AND2_X1 port map( A1 => N474, A2 => n105, ZN => n_state_stu_30_port);
   U61 : AND2_X1 port map( A1 => N146, A2 => n264, ZN => n_state_bpw_27_port);
   U62 : AND2_X1 port map( A1 => N143, A2 => n264, ZN => n_state_bpw_24_port);
   U63 : AND2_X1 port map( A1 => N149, A2 => n267, ZN => n_state_bpw_30_port);
   U64 : AND2_X1 port map( A1 => N148, A2 => n278_port, ZN => 
                           n_state_bpw_29_port);
   U65 : AND2_X1 port map( A1 => N147, A2 => n267, ZN => n_state_bpw_28_port);
   U66 : AND2_X1 port map( A1 => N145, A2 => n278_port, ZN => 
                           n_state_bpw_26_port);
   U67 : AND2_X1 port map( A1 => N144, A2 => n267, ZN => n_state_bpw_25_port);
   U68 : AND2_X1 port map( A1 => N142, A2 => n278_port, ZN => 
                           n_state_bpw_23_port);
   U69 : AND2_X1 port map( A1 => N141, A2 => n267, ZN => n_state_bpw_22_port);
   U70 : AND2_X1 port map( A1 => N76, A2 => n295_port, ZN => 
                           n_state_ral_30_port);
   U71 : AND2_X1 port map( A1 => N75, A2 => n295_port, ZN => 
                           n_state_ral_29_port);
   U72 : AND2_X1 port map( A1 => N73, A2 => n295_port, ZN => 
                           n_state_ral_27_port);
   U73 : AND2_X1 port map( A1 => N71, A2 => n295_port, ZN => 
                           n_state_ral_25_port);
   U74 : AND2_X1 port map( A1 => N69, A2 => n295_port, ZN => 
                           n_state_ral_23_port);
   U75 : AND3_X1 port map( A1 => n96, A2 => n45, A3 => n133_port, ZN => 
                           n132_port);
   U76 : INV_X1 port map( A => n299_port, ZN => n298_port);
   U77 : AND3_X1 port map( A1 => n85, A2 => n300_port, A3 => n279_port, ZN => 
                           n264);
   U78 : AND3_X1 port map( A1 => n85, A2 => n300_port, A3 => n279_port, ZN => 
                           n278_port);
   U79 : AND3_X1 port map( A1 => n85, A2 => n300_port, A3 => n279_port, ZN => 
                           n267);
   U80 : AND3_X1 port map( A1 => n96, A2 => n45, A3 => n133_port, ZN => 
                           n295_port);
   U81 : INV_X1 port map( A => n135_port, ZN => n76_port);
   U82 : AND2_X1 port map( A1 => N295, A2 => n291_port, ZN => 
                           n_state_div_17_port);
   U83 : AND2_X1 port map( A1 => N292, A2 => n291_port, ZN => 
                           n_state_div_14_port);
   U84 : AND2_X1 port map( A1 => N289, A2 => n291_port, ZN => 
                           n_state_div_11_port);
   U85 : AND2_X1 port map( A1 => N285, A2 => n291_port, ZN => 
                           n_state_div_7_port);
   U86 : AND2_X1 port map( A1 => N282, A2 => n291_port, ZN => 
                           n_state_div_4_port);
   U87 : AND2_X1 port map( A1 => N279, A2 => n291_port, ZN => 
                           n_state_div_1_port);
   U88 : AND2_X1 port map( A1 => N210, A2 => n293_port, ZN => 
                           n_state_mul_17_port);
   U89 : AND2_X1 port map( A1 => N207, A2 => n293_port, ZN => 
                           n_state_mul_14_port);
   U90 : AND2_X1 port map( A1 => N204, A2 => n293_port, ZN => 
                           n_state_mul_11_port);
   U91 : AND2_X1 port map( A1 => N200, A2 => n293_port, ZN => 
                           n_state_mul_7_port);
   U92 : AND2_X1 port map( A1 => N197, A2 => n293_port, ZN => 
                           n_state_mul_4_port);
   U93 : AND2_X1 port map( A1 => N194, A2 => n293_port, ZN => 
                           n_state_mul_1_port);
   U94 : AND2_X1 port map( A1 => N380, A2 => n297_port, ZN => 
                           n_state_sqrt_17_port);
   U95 : AND2_X1 port map( A1 => N377, A2 => n297_port, ZN => 
                           n_state_sqrt_14_port);
   U96 : AND2_X1 port map( A1 => N374, A2 => n297_port, ZN => 
                           n_state_sqrt_11_port);
   U97 : AND2_X1 port map( A1 => N370, A2 => n297_port, ZN => 
                           n_state_sqrt_7_port);
   U98 : AND2_X1 port map( A1 => N367, A2 => n297_port, ZN => 
                           n_state_sqrt_4_port);
   U99 : AND2_X1 port map( A1 => N364, A2 => n297_port, ZN => 
                           n_state_sqrt_1_port);
   U100 : AND2_X1 port map( A1 => N384, A2 => n296_port, ZN => 
                           n_state_sqrt_21_port);
   U101 : AND2_X1 port map( A1 => N382, A2 => n296_port, ZN => 
                           n_state_sqrt_19_port);
   U102 : AND2_X1 port map( A1 => N379, A2 => n296_port, ZN => 
                           n_state_sqrt_16_port);
   U103 : AND2_X1 port map( A1 => N376, A2 => n296_port, ZN => 
                           n_state_sqrt_13_port);
   U104 : AND2_X1 port map( A1 => N372, A2 => n296_port, ZN => 
                           n_state_sqrt_9_port);
   U105 : AND2_X1 port map( A1 => N369, A2 => n296_port, ZN => 
                           n_state_sqrt_6_port);
   U106 : AND2_X1 port map( A1 => N366, A2 => n296_port, ZN => 
                           n_state_sqrt_3_port);
   U107 : AND2_X1 port map( A1 => N365, A2 => n296_port, ZN => 
                           n_state_sqrt_2_port);
   U108 : AND2_X1 port map( A1 => N373, A2 => n296_port, ZN => 
                           n_state_sqrt_10_port);
   U109 : AND2_X1 port map( A1 => N299, A2 => n271, ZN => n_state_div_21_port);
   U110 : AND2_X1 port map( A1 => N297, A2 => n271, ZN => n_state_div_19_port);
   U111 : AND2_X1 port map( A1 => N294, A2 => n271, ZN => n_state_div_16_port);
   U112 : AND2_X1 port map( A1 => N291, A2 => n271, ZN => n_state_div_13_port);
   U113 : AND2_X1 port map( A1 => N287, A2 => n271, ZN => n_state_div_9_port);
   U114 : AND2_X1 port map( A1 => N284, A2 => n271, ZN => n_state_div_6_port);
   U115 : AND2_X1 port map( A1 => N281, A2 => n271, ZN => n_state_div_3_port);
   U116 : AND2_X1 port map( A1 => N280, A2 => n271, ZN => n_state_div_2_port);
   U117 : AND2_X1 port map( A1 => N288, A2 => n271, ZN => n_state_div_10_port);
   U118 : AND2_X1 port map( A1 => N214, A2 => n292_port, ZN => 
                           n_state_mul_21_port);
   U119 : AND2_X1 port map( A1 => N212, A2 => n292_port, ZN => 
                           n_state_mul_19_port);
   U120 : AND2_X1 port map( A1 => N209, A2 => n292_port, ZN => 
                           n_state_mul_16_port);
   U121 : AND2_X1 port map( A1 => N206, A2 => n292_port, ZN => 
                           n_state_mul_13_port);
   U122 : AND2_X1 port map( A1 => N202, A2 => n292_port, ZN => 
                           n_state_mul_9_port);
   U123 : AND2_X1 port map( A1 => N199, A2 => n292_port, ZN => 
                           n_state_mul_6_port);
   U124 : AND2_X1 port map( A1 => N196, A2 => n292_port, ZN => 
                           n_state_mul_3_port);
   U125 : AND2_X1 port map( A1 => N195, A2 => n292_port, ZN => 
                           n_state_mul_2_port);
   U126 : AND2_X1 port map( A1 => N203, A2 => n292_port, ZN => 
                           n_state_mul_10_port);
   U127 : AND2_X1 port map( A1 => N383, A2 => n116, ZN => n_state_sqrt_20_port)
                           ;
   U128 : AND2_X1 port map( A1 => N381, A2 => n116, ZN => n_state_sqrt_18_port)
                           ;
   U129 : AND2_X1 port map( A1 => N378, A2 => n116, ZN => n_state_sqrt_15_port)
                           ;
   U130 : AND2_X1 port map( A1 => N375, A2 => n116, ZN => n_state_sqrt_12_port)
                           ;
   U131 : AND2_X1 port map( A1 => N371, A2 => n116, ZN => n_state_sqrt_8_port);
   U132 : AND2_X1 port map( A1 => N368, A2 => n116, ZN => n_state_sqrt_5_port);
   U133 : AND2_X1 port map( A1 => N298, A2 => n255, ZN => n_state_div_20_port);
   U134 : AND2_X1 port map( A1 => N296, A2 => n255, ZN => n_state_div_18_port);
   U135 : AND2_X1 port map( A1 => N293, A2 => n255, ZN => n_state_div_15_port);
   U136 : AND2_X1 port map( A1 => N290, A2 => n255, ZN => n_state_div_12_port);
   U137 : AND2_X1 port map( A1 => N286, A2 => n255, ZN => n_state_div_8_port);
   U138 : AND2_X1 port map( A1 => N283, A2 => n255, ZN => n_state_div_5_port);
   U139 : AND2_X1 port map( A1 => N213, A2 => n146_port, ZN => 
                           n_state_mul_20_port);
   U140 : AND2_X1 port map( A1 => N211, A2 => n146_port, ZN => 
                           n_state_mul_18_port);
   U141 : AND2_X1 port map( A1 => N208, A2 => n146_port, ZN => 
                           n_state_mul_15_port);
   U142 : AND2_X1 port map( A1 => N205, A2 => n146_port, ZN => 
                           n_state_mul_12_port);
   U143 : AND2_X1 port map( A1 => N201, A2 => n146_port, ZN => 
                           n_state_mul_8_port);
   U144 : AND2_X1 port map( A1 => N198, A2 => n146_port, ZN => 
                           n_state_mul_5_port);
   U145 : AND2_X1 port map( A1 => N66, A2 => n132_port, ZN => 
                           n_state_ral_20_port);
   U146 : AND2_X1 port map( A1 => N65, A2 => n132_port, ZN => 
                           n_state_ral_19_port);
   U147 : AND2_X1 port map( A1 => N63, A2 => n132_port, ZN => 
                           n_state_ral_17_port);
   U148 : AND2_X1 port map( A1 => N61, A2 => n132_port, ZN => 
                           n_state_ral_15_port);
   U149 : AND2_X1 port map( A1 => N59, A2 => n132_port, ZN => 
                           n_state_ral_13_port);
   U150 : AND2_X1 port map( A1 => N57, A2 => n132_port, ZN => 
                           n_state_ral_11_port);
   U151 : AND2_X1 port map( A1 => N54, A2 => n132_port, ZN => 
                           n_state_ral_8_port);
   U152 : AND2_X1 port map( A1 => N52, A2 => n132_port, ZN => 
                           n_state_ral_6_port);
   U153 : AND2_X1 port map( A1 => N50, A2 => n132_port, ZN => 
                           n_state_ral_4_port);
   U154 : AND2_X1 port map( A1 => N48, A2 => n132_port, ZN => 
                           n_state_ral_2_port);
   U155 : AND2_X1 port map( A1 => N454, A2 => n298_port, ZN => 
                           n_state_stu_10_port);
   U156 : AND2_X1 port map( A1 => N455, A2 => n298_port, ZN => 
                           n_state_stu_11_port);
   U157 : AND2_X1 port map( A1 => N456, A2 => n298_port, ZN => 
                           n_state_stu_12_port);
   U158 : AND2_X1 port map( A1 => N457, A2 => n298_port, ZN => 
                           n_state_stu_13_port);
   U159 : AND2_X1 port map( A1 => N458, A2 => n298_port, ZN => 
                           n_state_stu_14_port);
   U160 : AND2_X1 port map( A1 => N459, A2 => n298_port, ZN => 
                           n_state_stu_15_port);
   U161 : AND2_X1 port map( A1 => N460, A2 => n298_port, ZN => 
                           n_state_stu_16_port);
   U162 : AND2_X1 port map( A1 => N461, A2 => n298_port, ZN => 
                           n_state_stu_17_port);
   U163 : AND2_X1 port map( A1 => N462, A2 => n298_port, ZN => 
                           n_state_stu_18_port);
   U164 : AND2_X1 port map( A1 => N463, A2 => n298_port, ZN => 
                           n_state_stu_19_port);
   U165 : AND2_X1 port map( A1 => N445, A2 => n298_port, ZN => 
                           n_state_stu_1_port);
   U166 : AND2_X1 port map( A1 => N464, A2 => n298_port, ZN => 
                           n_state_stu_20_port);
   U167 : AND2_X1 port map( A1 => N465, A2 => n105, ZN => n_state_stu_21_port);
   U168 : AND2_X1 port map( A1 => N447, A2 => n298_port, ZN => 
                           n_state_stu_3_port);
   U169 : AND2_X1 port map( A1 => N448, A2 => n105, ZN => n_state_stu_4_port);
   U170 : AND2_X1 port map( A1 => N449, A2 => n105, ZN => n_state_stu_5_port);
   U171 : AND2_X1 port map( A1 => N450, A2 => n105, ZN => n_state_stu_6_port);
   U172 : AND2_X1 port map( A1 => N451, A2 => n105, ZN => n_state_stu_7_port);
   U173 : AND2_X1 port map( A1 => N452, A2 => n298_port, ZN => 
                           n_state_stu_8_port);
   U174 : AND2_X1 port map( A1 => N453, A2 => n105, ZN => n_state_stu_9_port);
   U175 : AND2_X1 port map( A1 => N140, A2 => n264, ZN => n_state_bpw_21_port);
   U176 : AND2_X1 port map( A1 => N138, A2 => n264, ZN => n_state_bpw_19_port);
   U177 : AND2_X1 port map( A1 => N135, A2 => n264, ZN => n_state_bpw_16_port);
   U178 : AND2_X1 port map( A1 => N132, A2 => n264, ZN => n_state_bpw_13_port);
   U179 : AND2_X1 port map( A1 => N128, A2 => n264, ZN => n_state_bpw_9_port);
   U180 : AND2_X1 port map( A1 => N125, A2 => n264, ZN => n_state_bpw_6_port);
   U181 : AND2_X1 port map( A1 => N122, A2 => n264, ZN => n_state_bpw_3_port);
   U182 : AND2_X1 port map( A1 => N121, A2 => n264, ZN => n_state_bpw_2_port);
   U183 : AND2_X1 port map( A1 => N129, A2 => n264, ZN => n_state_bpw_10_port);
   U184 : AND2_X1 port map( A1 => N139, A2 => n278_port, ZN => 
                           n_state_bpw_20_port);
   U185 : AND2_X1 port map( A1 => N137, A2 => n278_port, ZN => 
                           n_state_bpw_18_port);
   U186 : AND2_X1 port map( A1 => N136, A2 => n267, ZN => n_state_bpw_17_port);
   U187 : AND2_X1 port map( A1 => N134, A2 => n278_port, ZN => 
                           n_state_bpw_15_port);
   U188 : AND2_X1 port map( A1 => N133, A2 => n267, ZN => n_state_bpw_14_port);
   U189 : AND2_X1 port map( A1 => N131, A2 => n278_port, ZN => 
                           n_state_bpw_12_port);
   U190 : AND2_X1 port map( A1 => N130, A2 => n267, ZN => n_state_bpw_11_port);
   U191 : AND2_X1 port map( A1 => N127, A2 => n278_port, ZN => 
                           n_state_bpw_8_port);
   U192 : AND2_X1 port map( A1 => N126, A2 => n267, ZN => n_state_bpw_7_port);
   U193 : AND2_X1 port map( A1 => N124, A2 => n278_port, ZN => 
                           n_state_bpw_5_port);
   U194 : AND2_X1 port map( A1 => N123, A2 => n267, ZN => n_state_bpw_4_port);
   U195 : AND2_X1 port map( A1 => N120, A2 => n267, ZN => n_state_bpw_1_port);
   U196 : AND2_X1 port map( A1 => N67, A2 => n295_port, ZN => 
                           n_state_ral_21_port);
   U197 : AND2_X1 port map( A1 => N62, A2 => n295_port, ZN => 
                           n_state_ral_16_port);
   U198 : AND2_X1 port map( A1 => N58, A2 => n295_port, ZN => 
                           n_state_ral_12_port);
   U199 : AND2_X1 port map( A1 => N55, A2 => n295_port, ZN => 
                           n_state_ral_9_port);
   U200 : AND2_X1 port map( A1 => N53, A2 => n295_port, ZN => 
                           n_state_ral_7_port);
   U201 : AND2_X1 port map( A1 => N51, A2 => n295_port, ZN => 
                           n_state_ral_5_port);
   U202 : AND2_X1 port map( A1 => N47, A2 => n295_port, ZN => 
                           n_state_ral_1_port);
   U203 : AND2_X1 port map( A1 => N64, A2 => n295_port, ZN => 
                           n_state_ral_18_port);
   U204 : AND2_X1 port map( A1 => N60, A2 => n295_port, ZN => 
                           n_state_ral_14_port);
   U205 : AND2_X1 port map( A1 => N49, A2 => n295_port, ZN => 
                           n_state_ral_3_port);
   U206 : AND2_X1 port map( A1 => N56, A2 => n295_port, ZN => 
                           n_state_ral_10_port);
   U207 : OR2_X1 port map( A1 => n299_port, A2 => N446, ZN => 
                           n_state_stu_2_port);
   U208 : AOI211_X1 port map( C1 => n50_port, C2 => c_state_div_5_port, A => 
                           n62_port, B => n68_port, ZN => n78);
   U209 : INV_X1 port map( A => sig_ral, ZN => n45);
   U210 : NAND4_X1 port map( A1 => n47_port, A2 => n39, A3 => n48_port, A4 => 
                           n49_port, ZN => stall_flag_1_port);
   U211 : OAI221_X1 port map( B1 => n53_port, B2 => n54_port, C1 => n55_port, 
                           C2 => n56_port, A => n57_port, ZN => n41);
   U212 : INV_X1 port map( A => n63_port, ZN => n56_port);
   U213 : AOI21_X1 port map( B1 => net108020, B2 => n67_port, A => n68_port, ZN
                           => n54_port);
   U214 : INV_X1 port map( A => n58_port, ZN => n57_port);
   U215 : NOR4_X1 port map( A1 => n112, A2 => c_state_stu_19_port, A3 => 
                           c_state_stu_17_port, A4 => c_state_stu_18_port, ZN 
                           => n111);
   U216 : NAND4_X1 port map( A1 => n213_port, A2 => n212_port, A3 => n211_port,
                           A4 => n210_port, ZN => n112);
   U217 : NOR4_X1 port map( A1 => n128_port, A2 => c_state_sqrt_14_port, A3 => 
                           c_state_sqrt_19_port, A4 => c_state_sqrt_15_port, ZN
                           => n127_port);
   U218 : NAND4_X1 port map( A1 => n235, A2 => n234, A3 => n233, A4 => n229, ZN
                           => n128_port);
   U219 : NOR4_X1 port map( A1 => n273, A2 => c_state_div_14_port, A3 => 
                           c_state_div_19_port, A4 => c_state_div_15_port, ZN 
                           => n272);
   U220 : NAND4_X1 port map( A1 => n244, A2 => n243, A3 => n242, A4 => n241, ZN
                           => n273);
   U221 : NOR4_X1 port map( A1 => n251, A2 => c_state_mul_10_port, A3 => 
                           c_state_mul_15_port, A4 => c_state_mul_14_port, ZN 
                           => n250);
   U222 : NAND4_X1 port map( A1 => n160, A2 => n159, A3 => n158, A4 => n157, ZN
                           => n251);
   U223 : OAI22_X1 port map( A1 => n59_port, A2 => n60_port, B1 => 
                           c_state_stu_0_port, B2 => n39, ZN => n58_port);
   U224 : AOI21_X1 port map( B1 => n50_port, B2 => n230, A => n62_port, ZN => 
                           n59_port);
   U225 : NAND4_X1 port map( A1 => n108, A2 => n109, A3 => n110, A4 => n111, ZN
                           => n87);
   U226 : NOR4_X1 port map( A1 => n115, A2 => c_state_stu_9_port, A3 => 
                           c_state_stu_7_port, A4 => c_state_stu_8_port, ZN => 
                           n108);
   U227 : NOR4_X1 port map( A1 => n114, A2 => c_state_stu_22_port, A3 => 
                           c_state_stu_16_port, A4 => c_state_stu_21_port, ZN 
                           => n109);
   U228 : NOR4_X1 port map( A1 => n113, A2 => c_state_stu_4_port, A3 => 
                           c_state_stu_27_port, A4 => c_state_stu_3_port, ZN =>
                           n110);
   U229 : AOI22_X1 port map( A1 => n90, A2 => n222_port, B1 => 
                           c_state_mul_3_port, B2 => c_state_mul_0_port, ZN => 
                           n89);
   U230 : INV_X1 port map( A => n94, ZN => n88);
   U231 : NOR2_X1 port map( A1 => c_state_mul_2_port, A2 => c_state_mul_1_port,
                           ZN => n90);
   U232 : INV_X1 port map( A => n87, ZN => n86);
   U233 : NAND4_X1 port map( A1 => n155, A2 => n348, A3 => n347, A4 => n344, ZN
                           => n260);
   U234 : NAND2_X1 port map( A1 => n163, A2 => n149_port, ZN => n65_port);
   U235 : NAND2_X1 port map( A1 => net108021, A2 => n265, ZN => n104);
   U236 : NAND4_X1 port map( A1 => net108010, A2 => net108009, A3 => net108008,
                           A4 => n276, ZN => n130_port);
   U237 : NAND4_X1 port map( A1 => net108040, A2 => net108039, A3 => net108038,
                           A4 => net108037, ZN => n252);
   U238 : NAND4_X1 port map( A1 => n311, A2 => n309_port, A3 => n308_port, A4 
                           => n307_port, ZN => n253);
   U239 : NAND4_X1 port map( A1 => n221_port, A2 => n220_port, A3 => n219_port,
                           A4 => n218_port, ZN => n113);
   U240 : NAND4_X1 port map( A1 => net107996, A2 => net107995, A3 => n227, A4 
                           => n226, ZN => n114);
   U241 : NAND4_X1 port map( A1 => net108003, A2 => net108002, A3 => net108001,
                           A4 => net108000, ZN => n115);
   U242 : NAND2_X1 port map( A1 => n194_port, A2 => n70_port, ZN => n39);
   U243 : NAND2_X1 port map( A1 => net108007, A2 => n123_port, ZN => n101);
   U244 : AND3_X1 port map( A1 => n310, A2 => n150_port, A3 => n312, ZN => 
                           n149_port);
   U245 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => stall_flag_3_port);
   U246 : INV_X1 port map( A => sig_jral, ZN => n37);
   U247 : AND4_X1 port map( A1 => n124_port, A2 => n125_port, A3 => n126_port, 
                           A4 => n127_port, ZN => n123_port);
   U248 : NOR4_X1 port map( A1 => n131_port, A2 => c_state_sqrt_6_port, A3 => 
                           c_state_sqrt_8_port, A4 => c_state_sqrt_7_port, ZN 
                           => n124_port);
   U249 : NOR4_X1 port map( A1 => n130_port, A2 => c_state_sqrt_17_port, A3 => 
                           c_state_sqrt_22_port, A4 => c_state_sqrt_18_port, ZN
                           => n125_port);
   U250 : NOR4_X1 port map( A1 => n129_port, A2 => c_state_sqrt_9_port, A3 => 
                           c_state_sqrt_30_port, A4 => c_state_sqrt_5_port, ZN 
                           => n126_port);
   U251 : AND4_X1 port map( A1 => n268, A2 => n269, A3 => n270, A4 => n272, ZN 
                           => n265);
   U252 : NOR4_X1 port map( A1 => n277, A2 => c_state_div_6_port, A3 => 
                           c_state_div_8_port, A4 => c_state_div_7_port, ZN => 
                           n268);
   U253 : NOR4_X1 port map( A1 => n275, A2 => c_state_div_17_port, A3 => 
                           c_state_div_22_port, A4 => c_state_div_18_port, ZN 
                           => n269);
   U254 : NOR4_X1 port map( A1 => n274, A2 => c_state_div_10_port, A3 => 
                           c_state_div_30_port, A4 => c_state_div_9_port, ZN =>
                           n270);
   U255 : AND4_X1 port map( A1 => n347, A2 => n344, A3 => n348, A4 => n258, ZN 
                           => n83);
   U256 : NOR4_X1 port map( A1 => n230, A2 => n155, A3 => n104, A4 => 
                           c_state_div_0_port, ZN => n258);
   U257 : AND4_X1 port map( A1 => n294_port, A2 => n149_port, A3 => 
                           c_state_mul_1_port, A4 => c_state_mul_3_port, ZN => 
                           n84);
   U258 : AND4_X1 port map( A1 => n119_port, A2 => n266, A3 => n247, A4 => 
                           n120_port, ZN => n82);
   U259 : NOR3_X1 port map( A1 => c_state_sqrt_2_port, A2 => net108020, A3 => 
                           n240, ZN => n120_port);
   U260 : AND4_X1 port map( A1 => n152, A2 => n153, A3 => n154, A4 => n250, ZN 
                           => n150_port);
   U261 : NOR4_X1 port map( A1 => n254, A2 => c_state_mul_4_port, A3 => 
                           c_state_mul_6_port, A4 => c_state_mul_5_port, ZN => 
                           n152);
   U262 : NOR4_X1 port map( A1 => n253, A2 => c_state_mul_9_port, A3 => 
                           c_state_mul_7_port, A4 => c_state_mul_8_port, ZN => 
                           n153);
   U263 : NOR4_X1 port map( A1 => n252, A2 => c_state_mul_23_port, A3 => 
                           c_state_mul_12_port, A4 => c_state_mul_11_port, ZN 
                           => n154);
   U264 : AND2_X1 port map( A1 => N394, A2 => n116, ZN => n_state_sqrt_31_port)
                           ;
   U265 : AND2_X1 port map( A1 => N309, A2 => n255, ZN => n_state_div_31_port);
   U266 : AND2_X1 port map( A1 => N224, A2 => n146_port, ZN => 
                           n_state_mul_31_port);
   U267 : AND2_X1 port map( A1 => N77, A2 => n132_port, ZN => 
                           n_state_ral_31_port);
   U268 : AND2_X1 port map( A1 => N475, A2 => n298_port, ZN => 
                           n_state_stu_31_port);
   U269 : AND2_X1 port map( A1 => N150, A2 => n278_port, ZN => 
                           n_state_bpw_31_port);
   U270 : AOI21_X1 port map( B1 => n259, B2 => net108021, A => n60_port, ZN => 
                           n291_port);
   U271 : AOI21_X1 port map( B1 => n94, B2 => n312, A => n55_port, ZN => 
                           n293_port);
   U272 : AOI21_X1 port map( B1 => n122_port, B2 => net108007, A => n53_port, 
                           ZN => n297_port);
   U273 : AOI21_X1 port map( B1 => n122_port, B2 => net108007, A => n53_port, 
                           ZN => n296_port);
   U274 : AOI21_X1 port map( B1 => n259, B2 => net108021, A => n60_port, ZN => 
                           n271);
   U275 : AOI21_X1 port map( B1 => n94, B2 => n312, A => n55_port, ZN => 
                           n292_port);
   U276 : AOI21_X1 port map( B1 => n122_port, B2 => net108007, A => n53_port, 
                           ZN => n116);
   U277 : AOI21_X1 port map( B1 => n259, B2 => net108021, A => n60_port, ZN => 
                           n255);
   U278 : AOI21_X1 port map( B1 => n94, B2 => n312, A => n55_port, ZN => 
                           n146_port);
   U279 : NOR4_X1 port map( A1 => n288_port, A2 => c_state_bpw_13_port, A3 => 
                           c_state_bpw_15_port, A4 => c_state_bpw_14_port, ZN 
                           => n284_port);
   U280 : NAND4_X1 port map( A1 => n176, A2 => n175, A3 => n174, A4 => n173, ZN
                           => n288_port);
   U281 : NOR4_X1 port map( A1 => n143_port, A2 => c_state_ral_13_port, A3 => 
                           c_state_ral_15_port, A4 => c_state_ral_14_port, ZN 
                           => n139_port);
   U282 : NAND4_X1 port map( A1 => n201_port, A2 => n200_port, A3 => n199_port,
                           A4 => n198_port, ZN => n143_port);
   U283 : INV_X1 port map( A => n72_port, ZN => n281_port);
   U284 : OAI21_X1 port map( B1 => n100, B2 => net108020, A => n123_port, ZN =>
                           n122_port);
   U285 : OAI21_X1 port map( B1 => n103, B2 => n230, A => n265, ZN => n259);
   U286 : NAND4_X1 port map( A1 => n282_port, A2 => n283_port, A3 => n284_port,
                           A4 => n285_port, ZN => n72_port);
   U287 : NOR2_X1 port map( A1 => n286_port, A2 => n287_port, ZN => n285_port);
   U288 : NOR4_X1 port map( A1 => n290_port, A2 => c_state_bpw_10_port, A3 => 
                           c_state_bpw_3_port, A4 => c_state_bpw_2_port, ZN => 
                           n282_port);
   U289 : NOR4_X1 port map( A1 => n289_port, A2 => c_state_bpw_17_port, A3 => 
                           c_state_bpw_4_port, A4 => c_state_bpw_18_port, ZN =>
                           n283_port);
   U290 : OAI21_X1 port map( B1 => n72_port, B2 => c_state_bpw_1_port, A => 
                           n164, ZN => n279_port);
   U291 : OAI21_X1 port map( B1 => n135_port, B2 => c_state_ral_1_port, A => 
                           n185, ZN => n133_port);
   U292 : NAND4_X1 port map( A1 => n137_port, A2 => n138_port, A3 => n139_port,
                           A4 => n140_port, ZN => n135_port);
   U293 : NOR2_X1 port map( A1 => n141_port, A2 => n142_port, ZN => n140_port);
   U294 : NOR4_X1 port map( A1 => n145_port, A2 => c_state_ral_10_port, A3 => 
                           c_state_ral_3_port, A4 => c_state_ral_2_port, ZN => 
                           n137_port);
   U295 : NOR4_X1 port map( A1 => n144_port, A2 => c_state_ral_17_port, A3 => 
                           c_state_ral_4_port, A4 => c_state_ral_18_port, ZN =>
                           n138_port);
   U296 : NAND2_X1 port map( A1 => n45, A2 => n134_port, ZN => 
                           n_state_ral_0_port);
   U297 : INV_X1 port map( A => n105, ZN => n299_port);
   U298 : OAI21_X1 port map( B1 => n107, B2 => n87, A => n228, ZN => n105);
   U299 : AOI21_X1 port map( B1 => n192, B2 => n194_port, A => n214_port, ZN =>
                           n107);
   U300 : NAND4_X1 port map( A1 => n183, A2 => n182, A3 => n181, A4 => n180, ZN
                           => n289_port);
   U301 : NAND4_X1 port map( A1 => net108051, A2 => net108050, A3 => net108049,
                           A4 => net108048, ZN => n290_port);
   U302 : NAND4_X1 port map( A1 => n208_port, A2 => n207_port, A3 => n206_port,
                           A4 => n205_port, ZN => n144_port);
   U303 : NAND4_X1 port map( A1 => net108060, A2 => net108059, A3 => net108058,
                           A4 => net108057, ZN => n145_port);
   U304 : NAND4_X1 port map( A1 => n172, A2 => n171, A3 => n170, A4 => n169, ZN
                           => n287_port);
   U305 : NAND4_X1 port map( A1 => n196_port, A2 => n193_port, A3 => n191, A4 
                           => n190, ZN => n142_port);
   U306 : NAND4_X1 port map( A1 => n168, A2 => n167, A3 => n166, A4 => n165, ZN
                           => n286_port);
   U307 : NAND4_X1 port map( A1 => n189, A2 => n188, A3 => n187, A4 => n186, ZN
                           => n141_port);
   U308 : OAI21_X1 port map( B1 => n256, B2 => n257, A => n46_port, ZN => 
                           n_state_div_0_port);
   U309 : INV_X1 port map( A => N278, ZN => n257);
   U310 : INV_X1 port map( A => n291_port, ZN => n256);
   U311 : OAI21_X1 port map( B1 => n147_port, B2 => n148_port, A => n44, ZN => 
                           n_state_mul_0_port);
   U312 : INV_X1 port map( A => N193, ZN => n148_port);
   U313 : INV_X1 port map( A => n293_port, ZN => n147_port);
   U314 : NAND2_X1 port map( A1 => n300_port, A2 => n280_port, ZN => 
                           n_state_bpw_0_port);
   U315 : INV_X1 port map( A => n117, ZN => n_state_sqrt_0_port);
   U316 : AOI21_X1 port map( B1 => n297_port, B2 => N363, A => n42, ZN => n117)
                           ;
   U317 : OR2_X1 port map( A1 => n299_port, A2 => N444, ZN => 
                           n_state_stu_0_port);
   U318 : AOI211_X1 port map( C1 => n50_port, C2 => c_state_div_0_port, A => 
                           n52_port, B => n41, ZN => n49_port);
   U319 : OAI22_X1 port map( A1 => n294_port, A2 => n65_port, B1 => n247, B2 =>
                           n69_port, ZN => n52_port);
   U320 : NOR4_X1 port map( A1 => n81, A2 => n82, A3 => n83, A4 => n84, ZN => 
                           n80);
   U321 : OAI211_X1 port map( C1 => n232, C2 => n85, A => n66_port, B => 
                           n75_port, ZN => n81);
   U322 : AOI21_X1 port map( B1 => n192, B2 => n70_port, A => n71_port, ZN => 
                           n48_port);
   U323 : NOR4_X1 port map( A1 => n197_port, A2 => n72_port, A3 => 
                           c_state_bpw_31_port, A4 => c_state_bpw_1_port, ZN =>
                           n71_port);
   U324 : NAND4_X1 port map( A1 => n231, A2 => n185, A3 => n76_port, A4 => 
                           c_state_ral_0_port, ZN => n47_port);
   U325 : INV_X1 port map( A => n95, ZN => n79);
   U326 : OAI222_X1 port map( A1 => n65_port, A2 => n222_port, B1 => n96, B2 =>
                           n231, C1 => n69_port, C2 => net108020, ZN => n95);
   U327 : BUF_X1 port map( A => rst, Z => n301_port);
   U328 : BUF_X1 port map( A => rst, Z => n302_port);
   U329 : BUF_X1 port map( A => rst, Z => n303_port);
   U330 : OAI211_X1 port map( C1 => n53_port, C2 => n82, A => n45, B => 
                           sig_sqrt, ZN => n118);
   U331 : INV_X1 port map( A => sig_bpw, ZN => n300_port);
   U332 : CLKBUF_X1 port map( A => n301_port, Z => n304_port);
   U350 : CLKBUF_X1 port map( A => n301_port, Z => n305_port);
   U351 : CLKBUF_X1 port map( A => n301_port, Z => n306_port);
   U352 : CLKBUF_X1 port map( A => n301_port, Z => n313);
   U353 : CLKBUF_X1 port map( A => n301_port, Z => n314);
   U354 : CLKBUF_X1 port map( A => n301_port, Z => n315);
   U355 : CLKBUF_X1 port map( A => n302_port, Z => n316);
   U356 : CLKBUF_X1 port map( A => n302_port, Z => n317);
   U357 : CLKBUF_X1 port map( A => n302_port, Z => n318);
   U358 : CLKBUF_X1 port map( A => n302_port, Z => n319);
   U359 : CLKBUF_X1 port map( A => n302_port, Z => n320);
   U360 : CLKBUF_X1 port map( A => n302_port, Z => n321);
   U361 : CLKBUF_X1 port map( A => n303_port, Z => n322);
   U362 : CLKBUF_X1 port map( A => n303_port, Z => n323);
   U363 : CLKBUF_X1 port map( A => n303_port, Z => n324);
   U364 : CLKBUF_X1 port map( A => n303_port, Z => n325);

end SYN_stall_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity CwGenerator_DATA_SIZE32_OPCD_SIZE6_FUNC_SIZE11_CWRD_SIZE20_CALU_SIZE5 is

   port( clk, rst : in std_logic;  opcd : in std_logic_vector (5 downto 0);  
         func : in std_logic_vector (10 downto 0);  stall_flag : in 
         std_logic_vector (4 downto 0);  taken : in std_logic;  cw : out 
         std_logic_vector (19 downto 0);  calu : out std_logic_vector (4 downto
         0));

end CwGenerator_DATA_SIZE32_OPCD_SIZE6_FUNC_SIZE11_CWRD_SIZE20_CALU_SIZE5;

architecture SYN_cw_generator_arch of 
   CwGenerator_DATA_SIZE32_OPCD_SIZE6_FUNC_SIZE11_CWRD_SIZE20_CALU_SIZE5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal cw_0_port, calu_4_port, calu_3_port, calu_2_port, calu_1_port, n12, 
      cw_2_port, cw_1_port, net107993, n4, n5, calu_0_port, n7, n8, n9, n10, 
      n11 : std_logic;

begin
   cw <= ( cw_2_port, cw_2_port, cw_2_port, cw_2_port, cw_2_port, cw_2_port, 
      cw_2_port, cw_2_port, cw_2_port, cw_2_port, cw_2_port, cw_2_port, 
      cw_2_port, cw_2_port, cw_2_port, cw_2_port, cw_2_port, cw_2_port, 
      cw_1_port, cw_0_port );
   calu <= ( calu_4_port, calu_3_port, calu_2_port, calu_1_port, calu_0_port );
   
   calu_reg_3_inst : DFF_X1 port map( D => n10, CK => clk, Q => calu_3_port, QN
                           => n9);
   calu_reg_2_inst : DFF_X1 port map( D => calu_2_port, CK => clk, Q => 
                           calu_2_port, QN => net107993);
   cw_2_port <= '0';
   calu_reg_4_inst : DFF_X1 port map( D => n8, CK => clk, Q => calu_4_port, QN 
                           => n7);
   calu_reg_1_inst : DFF_X1 port map( D => calu_1_port, CK => clk, Q => 
                           calu_1_port, QN => n11);
   calu_reg_0_inst : DFF_X1 port map( D => n12, CK => clk, Q => n12, QN => n5);
   U3 : NOR2_X1 port map( A1 => n4, A2 => stall_flag(3), ZN => cw_1_port);
   U4 : INV_X1 port map( A => taken, ZN => n4);
   U5 : INV_X2 port map( A => n5, ZN => calu_0_port);
   U7 : INV_X1 port map( A => n7, ZN => n8);
   U8 : INV_X1 port map( A => n9, ZN => n10);
   U9 : INV_X1 port map( A => stall_flag(4), ZN => cw_0_port);

end SYN_cw_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity 
   DataPath_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_OPCD_SIZE6_IMME_SIZE16_CWRD_SIZE20_CALU_SIZE5_DRCW_SIZE4 
   is

   port( clk, rst : in std_logic;  istr_addr : out std_logic_vector (31 downto 
         0);  istr_val : in std_logic_vector (31 downto 0);  ir_out, pc_out, 
         reg_a_out, ld_a_out, data_addr : out std_logic_vector (31 downto 0);  
         data_i_val : in std_logic_vector (31 downto 0);  data_o_val : out 
         std_logic_vector (31 downto 0);  cw : in std_logic_vector (19 downto 
         0);  dr_cw : out std_logic_vector (3 downto 0);  calu : in 
         std_logic_vector (4 downto 0);  sig_bal : out std_logic;  sig_bpw : in
         std_logic;  sig_jral, sig_ral, sig_mul, sig_div, sig_sqrt : out 
         std_logic);

end 
   DataPath_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_OPCD_SIZE6_IMME_SIZE16_CWRD_SIZE20_CALU_SIZE5_DRCW_SIZE4;

architecture SYN_data_path_arch of 
   DataPath_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_OPCD_SIZE6_IMME_SIZE16_CWRD_SIZE20_CALU_SIZE5_DRCW_SIZE4 
   is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component Reg_DATA_SIZE5_1
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 
            0);  dout : out std_logic_vector (4 downto 0));
   end component;
   
   component Reg_DATA_SIZE32_2
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 
            0);  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Reg_DATA_SIZE5_2
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 
            0);  dout : out std_logic_vector (4 downto 0));
   end component;
   
   component Reg_DATA_SIZE32_3
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 
            0);  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Mux_DATA_SIZE32_2
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0)
            ;  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_1
      port( reg_c, reg_f, reg_ff : in std_logic_vector (31 downto 0);  addr_c, 
            addr_f, addr_ff : in std_logic_vector (4 downto 0);  valid_f, 
            valid_ff, dirty_f, dirty_ff, en : in std_logic;  output : out 
            std_logic_vector (31 downto 0);  match_dirty_f, match_dirty_ff : 
            out std_logic);
   end component;
   
   component Reg_DATA_SIZE32_4
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 
            0);  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Reg_DATA_SIZE32_5
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 
            0);  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Reg_DATA_SIZE5_3
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 
            0);  dout : out std_logic_vector (4 downto 0));
   end component;
   
   component Reg_DATA_SIZE5_4
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 
            0);  dout : out std_logic_vector (4 downto 0));
   end component;
   
   component Reg_DATA_SIZE32_6
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 
            0);  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Reg_DATA_SIZE32_7
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 
            0);  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Mux4_DATA_SIZE32
      port( sel : in std_logic_vector (1 downto 0);  din0, din1, din2, din3 : 
            in std_logic_vector (31 downto 0);  dout : out std_logic_vector (31
            downto 0));
   end component;
   
   component Div_DATA_SIZE32_DIV_STAGE34_SQRT_STAGE18
      port( rst, clk, en, lock, sign, func : in std_logic;  a, b : in 
            std_logic_vector (31 downto 0);  o : out std_logic_vector (31 
            downto 0));
   end component;
   
   component Mul_DATA_SIZE16_STAGE10
      port( rst, clk, en, lock, sign : in std_logic;  a, b : in 
            std_logic_vector (15 downto 0);  o : out std_logic_vector (31 
            downto 0));
   end component;
   
   component Alu_DATA_SIZE32
      port( f : in std_logic_vector (4 downto 0);  a, b : in std_logic_vector 
            (31 downto 0);  o : out std_logic_vector (31 downto 0));
   end component;
   
   component Mux_DATA_SIZE32_3
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0)
            ;  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_2
      port( reg_c, reg_f, reg_ff : in std_logic_vector (31 downto 0);  addr_c, 
            addr_f, addr_ff : in std_logic_vector (4 downto 0);  valid_f, 
            valid_ff, dirty_f, dirty_ff, en : in std_logic;  output : out 
            std_logic_vector (31 downto 0);  match_dirty_f, match_dirty_ff : 
            out std_logic);
   end component;
   
   component FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_3
      port( reg_c, reg_f, reg_ff : in std_logic_vector (31 downto 0);  addr_c, 
            addr_f, addr_ff : in std_logic_vector (4 downto 0);  valid_f, 
            valid_ff, dirty_f, dirty_ff, en : in std_logic;  output : out 
            std_logic_vector (31 downto 0);  match_dirty_f, match_dirty_ff : 
            out std_logic);
   end component;
   
   component Mux_DATA_SIZE32_4
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0)
            ;  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Mux_DATA_SIZE32_5
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0)
            ;  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Reg_DATA_SIZE32_8
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 
            0);  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Reg_DATA_SIZE5_5
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 
            0);  dout : out std_logic_vector (4 downto 0));
   end component;
   
   component Reg_DATA_SIZE5_6
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 
            0);  dout : out std_logic_vector (4 downto 0));
   end component;
   
   component Reg_DATA_SIZE5_0
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 
            0);  dout : out std_logic_vector (4 downto 0));
   end component;
   
   component Reg_DATA_SIZE32_9
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 
            0);  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Reg_DATA_SIZE32_10
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 
            0);  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Reg_DATA_SIZE32_11
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 
            0);  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_4
      port( reg_c, reg_f, reg_ff : in std_logic_vector (31 downto 0);  addr_c, 
            addr_f, addr_ff : in std_logic_vector (4 downto 0);  valid_f, 
            valid_ff, dirty_f, dirty_ff, en : in std_logic;  output : out 
            std_logic_vector (31 downto 0);  match_dirty_f, match_dirty_ff : 
            out std_logic);
   end component;
   
   component FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_0
      port( reg_c, reg_f, reg_ff : in std_logic_vector (31 downto 0);  addr_c, 
            addr_f, addr_ff : in std_logic_vector (4 downto 0);  valid_f, 
            valid_ff, dirty_f, dirty_ff, en : in std_logic;  output : out 
            std_logic_vector (31 downto 0);  match_dirty_f, match_dirty_ff : 
            out std_logic);
   end component;
   
   component Mux_DATA_SIZE32_6
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0)
            ;  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Adder_DATA_SIZE32_7
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;
   
   component Mux_DATA_SIZE32_7
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0)
            ;  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component RegisterFile_DATA_SIZE32_REG_NUM32
      port( clk, rst, en, rd1_en, rd2_en, wr_en, link_en : in std_logic;  
            rd1_addr, rd2_addr, wr_addr : in std_logic_vector (4 downto 0);  
            d_out1, d_out2 : out std_logic_vector (31 downto 0);  d_in, d_link 
            : in std_logic_vector (31 downto 0));
   end component;
   
   component Extender_SRC_SIZE26_DEST_SIZE32
      port( s : in std_logic;  i : in std_logic_vector (25 downto 0);  o : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component Extender_SRC_SIZE16_DEST_SIZE32
      port( s : in std_logic;  i : in std_logic_vector (15 downto 0);  o : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component Mux_DATA_SIZE5
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (4 downto 0);
            dout : out std_logic_vector (4 downto 0));
   end component;
   
   component Mux_DATA_SIZE32_8
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0)
            ;  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Mux_DATA_SIZE32_9
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0)
            ;  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Reg_DATA_SIZE32_12
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 
            0);  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Reg_DATA_SIZE32_0
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 
            0);  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Mux_DATA_SIZE32_0
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0)
            ;  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Adder_DATA_SIZE32_0
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, istr_addr_31_port, istr_addr_30_port, 
      istr_addr_29_port, n120, istr_addr_27_port, istr_addr_26_port, 
      istr_addr_25_port, istr_addr_24_port, istr_addr_23_port, 
      istr_addr_22_port, istr_addr_21_port, istr_addr_20_port, 
      istr_addr_19_port, istr_addr_18_port, istr_addr_17_port, 
      istr_addr_16_port, istr_addr_15_port, istr_addr_14_port, 
      istr_addr_13_port, istr_addr_12_port, istr_addr_11_port, 
      istr_addr_10_port, istr_addr_9_port, istr_addr_8_port, istr_addr_7_port, 
      istr_addr_6_port, istr_addr_5_port, istr_addr_4_port, istr_addr_3_port, 
      n121, n122, n123, data_addr_31_port, data_addr_30_port, data_addr_29_port
      , data_addr_28_port, data_addr_27_port, data_addr_26_port, 
      data_addr_25_port, data_addr_24_port, data_addr_23_port, 
      data_addr_22_port, data_addr_21_port, data_addr_20_port, 
      data_addr_19_port, data_addr_18_port, data_addr_17_port, 
      data_addr_16_port, data_addr_15_port, data_addr_14_port, 
      data_addr_13_port, data_addr_12_port, data_addr_11_port, 
      data_addr_10_port, data_addr_9_port, data_addr_8_port, data_addr_7_port, 
      data_addr_6_port, data_addr_5_port, data_addr_4_port, data_addr_3_port, 
      data_addr_2_port, data_addr_1_port, data_addr_0_port, sig_ral_port, 
      sig_div_port, s1_npc_31_port, s1_npc_30_port, s1_npc_29_port, 
      s1_npc_28_port, s1_npc_27_port, s1_npc_26_port, s1_npc_25_port, 
      s1_npc_24_port, s1_npc_23_port, s1_npc_22_port, s1_npc_21_port, 
      s1_npc_20_port, s1_npc_19_port, s1_npc_18_port, s1_npc_17_port, 
      s1_npc_16_port, s1_npc_15_port, s1_npc_14_port, s1_npc_13_port, 
      s1_npc_12_port, s1_npc_11_port, s1_npc_10_port, s1_npc_9_port, 
      s1_npc_8_port, s1_npc_7_port, s1_npc_6_port, s1_npc_5_port, s1_npc_4_port
      , s1_npc_3_port, s1_npc_2_port, s1_npc_1_port, s1_npc_0_port, 
      s2_pc_sel_31_port, s2_pc_sel_30_port, s2_pc_sel_29_port, 
      s2_pc_sel_28_port, s2_pc_sel_27_port, s2_pc_sel_26_port, 
      s2_pc_sel_25_port, s2_pc_sel_24_port, s2_pc_sel_23_port, 
      s2_pc_sel_22_port, s2_pc_sel_21_port, s2_pc_sel_20_port, 
      s2_pc_sel_19_port, s2_pc_sel_18_port, s2_pc_sel_17_port, 
      s2_pc_sel_16_port, s2_pc_sel_15_port, s2_pc_sel_14_port, 
      s2_pc_sel_13_port, s2_pc_sel_12_port, s2_pc_sel_11_port, 
      s2_pc_sel_10_port, s2_pc_sel_9_port, s2_pc_sel_8_port, s2_pc_sel_7_port, 
      s2_pc_sel_6_port, s2_pc_sel_5_port, s2_pc_sel_4_port, s2_pc_sel_3_port, 
      s2_pc_sel_2_port, s2_pc_sel_1_port, s2_pc_sel_0_port, 
      s3_pc_notsel_31_port, s3_pc_notsel_30_port, s3_pc_notsel_29_port, 
      s3_pc_notsel_28_port, s3_pc_notsel_27_port, s3_pc_notsel_26_port, 
      s3_pc_notsel_25_port, s3_pc_notsel_24_port, s3_pc_notsel_23_port, 
      s3_pc_notsel_22_port, s3_pc_notsel_21_port, s3_pc_notsel_20_port, 
      s3_pc_notsel_19_port, s3_pc_notsel_18_port, s3_pc_notsel_17_port, 
      s3_pc_notsel_16_port, s3_pc_notsel_15_port, s3_pc_notsel_14_port, 
      s3_pc_notsel_13_port, s3_pc_notsel_12_port, s3_pc_notsel_11_port, 
      s3_pc_notsel_10_port, s3_pc_notsel_9_port, s3_pc_notsel_8_port, 
      s3_pc_notsel_7_port, s3_pc_notsel_6_port, s3_pc_notsel_5_port, 
      s3_pc_notsel_4_port, s3_pc_notsel_3_port, s3_pc_notsel_2_port, 
      s3_pc_notsel_1_port, s3_pc_notsel_0_port, s2_npc_31_port, s2_npc_30_port,
      s2_npc_29_port, s2_npc_28_port, s2_npc_27_port, s2_npc_26_port, 
      s2_npc_25_port, s2_npc_24_port, s2_npc_23_port, s2_npc_22_port, 
      s2_npc_21_port, s2_npc_20_port, s2_npc_19_port, s2_npc_18_port, 
      s2_npc_17_port, s2_npc_16_port, s2_npc_15_port, s2_npc_14_port, 
      s2_npc_13_port, s2_npc_12_port, s2_npc_11_port, s2_npc_10_port, 
      s2_npc_9_port, s2_npc_8_port, s2_npc_7_port, s2_npc_6_port, s2_npc_5_port
      , s2_npc_4_port, s2_npc_3_port, s2_npc_2_port, s2_npc_1_port, 
      s2_npc_0_port, s2_jpc_30_port, s2_jpc_29_port, s2_jpc_28_port, 
      s2_jpc_27_port, s2_jpc_26_port, s2_jpc_25_port, s2_jpc_24_port, 
      s2_jpc_23_port, s2_jpc_22_port, s2_jpc_21_port, s2_jpc_20_port, 
      s2_jpc_19_port, s2_jpc_18_port, s2_jpc_17_port, s2_jpc_16_port, 
      s2_jpc_15_port, s2_jpc_14_port, s2_jpc_13_port, s2_jpc_12_port, 
      s2_jpc_11_port, s2_jpc_10_port, s2_jpc_9_port, s2_jpc_8_port, 
      s2_jpc_7_port, s2_jpc_6_port, s2_jpc_5_port, s2_jpc_4_port, s2_jpc_3_port
      , s2_jpc_2_port, s2_jpc_1_port, s2_jpc_0_port, s2_pc_notsel_31_port, 
      s2_pc_notsel_30_port, s2_pc_notsel_29_port, s2_pc_notsel_28_port, 
      s2_pc_notsel_27_port, s2_pc_notsel_26_port, s2_pc_notsel_25_port, 
      s2_pc_notsel_24_port, s2_pc_notsel_23_port, s2_pc_notsel_22_port, 
      s2_pc_notsel_21_port, s2_pc_notsel_20_port, s2_pc_notsel_19_port, 
      s2_pc_notsel_18_port, s2_pc_notsel_17_port, s2_pc_notsel_16_port, 
      s2_pc_notsel_15_port, s2_pc_notsel_14_port, s2_pc_notsel_13_port, 
      s2_pc_notsel_12_port, s2_pc_notsel_11_port, s2_pc_notsel_10_port, 
      s2_pc_notsel_9_port, s2_pc_notsel_8_port, s2_pc_notsel_7_port, 
      s2_pc_notsel_6_port, s2_pc_notsel_5_port, s2_pc_notsel_4_port, 
      s2_pc_notsel_3_port, s2_pc_notsel_2_port, s2_pc_notsel_1_port, 
      s2_pc_notsel_0_port, s2_wr_addr_sel, s2_wr_addr_4_port, s2_wr_addr_3_port
      , s2_wr_addr_2_port, s2_wr_addr_1_port, s2_wr_addr_0_port, 
      s2_imm_l_ext_31_port, s2_imm_l_ext_15_port, s2_imm_l_ext_14_port, 
      s2_imm_l_ext_13_port, s2_imm_l_ext_12_port, s2_imm_l_ext_11_port, 
      s2_imm_l_ext_10_port, s2_imm_l_ext_9_port, s2_imm_l_ext_8_port, 
      s2_imm_l_ext_7_port, s2_imm_l_ext_6_port, s2_imm_l_ext_5_port, 
      s2_imm_l_ext_4_port, s2_imm_l_ext_3_port, s2_imm_l_ext_2_port, 
      s2_imm_l_ext_1_port, s2_imm_l_ext_0_port, s2_imm_j_ext_31_port, 
      s2_imm_j_ext_30_port, s2_imm_j_ext_29_port, s2_imm_j_ext_28_port, 
      s2_imm_j_ext_27_port, s2_imm_j_ext_26_port, s2_imm_j_ext_25_port, 
      s2_imm_j_ext_24_port, s2_imm_j_ext_23_port, s2_imm_j_ext_22_port, 
      s2_imm_j_ext_21_port, s2_imm_j_ext_20_port, s2_imm_j_ext_19_port, 
      s2_imm_j_ext_18_port, s2_imm_j_ext_17_port, s2_imm_j_ext_16_port, 
      s2_imm_j_ext_15_port, s2_imm_j_ext_14_port, s2_imm_j_ext_13_port, 
      s2_imm_j_ext_12_port, s2_imm_j_ext_11_port, s2_imm_j_ext_10_port, 
      s2_imm_j_ext_9_port, s2_imm_j_ext_8_port, s2_imm_j_ext_7_port, 
      s2_imm_j_ext_6_port, s2_imm_j_ext_5_port, s2_imm_j_ext_4_port, 
      s2_imm_j_ext_3_port, s2_imm_j_ext_2_port, s2_imm_j_ext_1_port, 
      s2_imm_j_ext_0_port, s2_imm_i_ext_31_port, s2_imm_i_ext_30_port, 
      s2_imm_i_ext_29_port, s2_imm_i_ext_28_port, s2_imm_i_ext_27_port, 
      s2_imm_i_ext_26_port, s2_imm_i_ext_25_port, s2_imm_i_ext_24_port, 
      s2_imm_i_ext_23_port, s2_imm_i_ext_22_port, s2_imm_i_ext_21_port, 
      s2_imm_i_ext_20_port, s2_imm_i_ext_19_port, s2_imm_i_ext_18_port, 
      s2_imm_i_ext_17_port, s2_imm_i_ext_16_port, s2_imm_i_ext_15_port, 
      s2_imm_i_ext_14_port, s2_imm_i_ext_13_port, s2_imm_i_ext_12_port, 
      s2_imm_i_ext_11_port, s2_imm_i_ext_10_port, s2_imm_i_ext_9_port, 
      s2_imm_i_ext_8_port, s2_imm_i_ext_7_port, s2_imm_i_ext_6_port, 
      s2_imm_i_ext_5_port, s2_imm_i_ext_4_port, s2_imm_i_ext_3_port, 
      s2_imm_i_ext_2_port, s2_imm_i_ext_1_port, s2_imm_i_ext_0_port, s2_rf_en, 
      s5_wr_addr_4_port, s5_wr_addr_3_port, s5_wr_addr_2_port, 
      s5_wr_addr_1_port, s5_wr_addr_0_port, s2_a_31_port, s2_a_30_port, 
      s2_a_29_port, s2_a_28_port, s2_a_27_port, s2_a_26_port, s2_a_25_port, 
      s2_a_24_port, s2_a_23_port, s2_a_22_port, s2_a_21_port, s2_a_20_port, 
      s2_a_19_port, s2_a_18_port, s2_a_17_port, s2_a_16_port, s2_a_15_port, 
      s2_a_14_port, s2_a_13_port, s2_a_12_port, s2_a_11_port, s2_a_10_port, 
      s2_a_9_port, s2_a_8_port, s2_a_7_port, s2_a_6_port, s2_a_5_port, 
      s2_a_4_port, s2_a_3_port, s2_a_2_port, s2_a_1_port, s2_a_0_port, 
      s2_b_31_port, s2_b_30_port, s2_b_29_port, s2_b_28_port, s2_b_27_port, 
      s2_b_26_port, s2_b_25_port, s2_b_24_port, s2_b_23_port, s2_b_22_port, 
      s2_b_21_port, s2_b_20_port, s2_b_19_port, s2_b_18_port, s2_b_17_port, 
      s2_b_16_port, s2_b_15_port, s2_b_14_port, s2_b_13_port, s2_b_12_port, 
      s2_b_11_port, s2_b_10_port, s2_b_9_port, s2_b_8_port, s2_b_7_port, 
      s2_b_6_port, s2_b_5_port, s2_b_4_port, s2_b_3_port, s2_b_2_port, 
      s2_b_1_port, s2_b_0_port, s5_result_31_port, s5_result_30_port, 
      s5_result_29_port, s5_result_28_port, s5_result_27_port, 
      s5_result_26_port, s5_result_25_port, s5_result_24_port, 
      s5_result_23_port, s5_result_22_port, s5_result_21_port, 
      s5_result_20_port, s5_result_19_port, s5_result_18_port, 
      s5_result_17_port, s5_result_16_port, s5_result_15_port, 
      s5_result_14_port, s5_result_13_port, s5_result_12_port, 
      s5_result_11_port, s5_result_10_port, s5_result_9_port, s5_result_8_port,
      s5_result_7_port, s5_result_6_port, s5_result_5_port, s5_result_4_port, 
      s5_result_3_port, s5_result_2_port, s5_result_1_port, s5_result_0_port, 
      s2_jump_addr_imm_31_port, s2_jump_addr_imm_30_port, 
      s2_jump_addr_imm_29_port, s2_jump_addr_imm_28_port, 
      s2_jump_addr_imm_27_port, s2_jump_addr_imm_26_port, 
      s2_jump_addr_imm_25_port, s2_jump_addr_imm_24_port, 
      s2_jump_addr_imm_23_port, s2_jump_addr_imm_22_port, 
      s2_jump_addr_imm_21_port, s2_jump_addr_imm_20_port, 
      s2_jump_addr_imm_19_port, s2_jump_addr_imm_18_port, 
      s2_jump_addr_imm_17_port, s2_jump_addr_imm_16_port, 
      s2_jump_addr_imm_15_port, s2_jump_addr_imm_14_port, 
      s2_jump_addr_imm_13_port, s2_jump_addr_imm_12_port, 
      s2_jump_addr_imm_11_port, s2_jump_addr_imm_10_port, 
      s2_jump_addr_imm_9_port, s2_jump_addr_imm_8_port, s2_jump_addr_imm_7_port
      , s2_jump_addr_imm_6_port, s2_jump_addr_imm_5_port, 
      s2_jump_addr_imm_4_port, s2_jump_addr_imm_3_port, s2_jump_addr_imm_2_port
      , s2_jump_addr_imm_1_port, s2_jump_addr_imm_0_port, 
      s2_jump_addr_rel_31_port, s2_jump_addr_rel_30_port, 
      s2_jump_addr_rel_29_port, s2_jump_addr_rel_28_port, 
      s2_jump_addr_rel_27_port, s2_jump_addr_rel_26_port, 
      s2_jump_addr_rel_25_port, s2_jump_addr_rel_24_port, 
      s2_jump_addr_rel_23_port, s2_jump_addr_rel_22_port, 
      s2_jump_addr_rel_21_port, s2_jump_addr_rel_20_port, 
      s2_jump_addr_rel_19_port, s2_jump_addr_rel_18_port, 
      s2_jump_addr_rel_17_port, s2_jump_addr_rel_16_port, 
      s2_jump_addr_rel_15_port, s2_jump_addr_rel_14_port, 
      s2_jump_addr_rel_13_port, s2_jump_addr_rel_12_port, 
      s2_jump_addr_rel_11_port, s2_jump_addr_rel_10_port, 
      s2_jump_addr_rel_9_port, s2_jump_addr_rel_8_port, s2_jump_addr_rel_7_port
      , s2_jump_addr_rel_6_port, s2_jump_addr_rel_5_port, 
      s2_jump_addr_rel_4_port, s2_jump_addr_rel_3_port, s2_jump_addr_rel_2_port
      , s2_jump_addr_rel_1_port, s2_jump_addr_rel_0_port, 
      s2_jump_addr_reg_31_port, s2_jump_addr_reg_30_port, 
      s2_jump_addr_reg_29_port, s2_jump_addr_reg_28_port, 
      s2_jump_addr_reg_27_port, s2_jump_addr_reg_26_port, 
      s2_jump_addr_reg_25_port, s2_jump_addr_reg_24_port, 
      s2_jump_addr_reg_23_port, s2_jump_addr_reg_22_port, 
      s2_jump_addr_reg_21_port, s2_jump_addr_reg_20_port, 
      s2_jump_addr_reg_19_port, s2_jump_addr_reg_18_port, 
      s2_jump_addr_reg_17_port, s2_jump_addr_reg_16_port, 
      s2_jump_addr_reg_15_port, s2_jump_addr_reg_14_port, 
      s2_jump_addr_reg_13_port, s2_jump_addr_reg_12_port, 
      s2_jump_addr_reg_11_port, s2_jump_addr_reg_10_port, 
      s2_jump_addr_reg_9_port, s2_jump_addr_reg_8_port, s2_jump_addr_reg_7_port
      , s2_jump_addr_reg_6_port, s2_jump_addr_reg_5_port, 
      s2_jump_addr_reg_4_port, s2_jump_addr_reg_3_port, s2_jump_addr_reg_2_port
      , s2_jump_addr_reg_1_port, s2_jump_addr_reg_0_port, s2_a_f_b_en, 
      s2_a_ff_b_en, s3_exe_out_31_port, s3_exe_out_30_port, s3_exe_out_29_port,
      s3_exe_out_28_port, s3_exe_out_27_port, s3_exe_out_26_port, 
      s3_exe_out_25_port, s3_exe_out_24_port, s3_exe_out_23_port, 
      s3_exe_out_22_port, s3_exe_out_21_port, s3_exe_out_20_port, 
      s3_exe_out_19_port, s3_exe_out_18_port, s3_exe_out_17_port, 
      s3_exe_out_16_port, s3_exe_out_15_port, s3_exe_out_14_port, 
      s3_exe_out_13_port, s3_exe_out_12_port, s3_exe_out_11_port, 
      s3_exe_out_10_port, s3_exe_out_9_port, s3_exe_out_8_port, 
      s3_exe_out_7_port, s3_exe_out_6_port, s3_exe_out_5_port, 
      s3_exe_out_4_port, s3_exe_out_3_port, s3_exe_out_2_port, 
      s3_exe_out_1_port, s3_exe_out_0_port, s4_result_31_port, 
      s4_result_30_port, s4_result_29_port, s4_result_28_port, 
      s4_result_27_port, s4_result_26_port, s4_result_25_port, 
      s4_result_24_port, s4_result_23_port, s4_result_22_port, 
      s4_result_21_port, s4_result_20_port, s4_result_19_port, 
      s4_result_18_port, s4_result_17_port, s4_result_16_port, 
      s4_result_15_port, s4_result_14_port, s4_result_13_port, 
      s4_result_12_port, s4_result_11_port, s4_result_10_port, s4_result_9_port
      , s4_result_8_port, s4_result_7_port, s4_result_6_port, s4_result_5_port,
      s4_result_4_port, s4_result_3_port, s4_result_2_port, s4_result_1_port, 
      s4_result_0_port, s3_wr_addr_4_port, s3_wr_addr_3_port, s3_wr_addr_2_port
      , s3_wr_addr_1_port, s3_wr_addr_0_port, s4_wr_addr_4_port, 
      s4_wr_addr_3_port, s4_wr_addr_2_port, s4_wr_addr_1_port, 
      s4_wr_addr_0_port, s2_a_f_j_en, s2_a_ff_j_en, s3_a_31_port, s3_a_30_port,
      s3_a_29_port, s3_a_28_port, s3_a_27_port, s3_a_26_port, s3_a_25_port, 
      s3_a_24_port, s3_a_23_port, s3_a_22_port, s3_a_21_port, s3_a_20_port, 
      s3_a_19_port, s3_a_18_port, s3_a_17_port, s3_a_16_port, s3_a_15_port, 
      s3_a_14_port, s3_a_13_port, s3_a_12_port, s3_a_11_port, s3_a_10_port, 
      s3_a_9_port, s3_a_8_port, s3_a_7_port, s3_a_6_port, s3_a_5_port, 
      s3_a_4_port, s3_a_3_port, s3_a_2_port, s3_a_1_port, s3_a_0_port, 
      s3_b_31_port, s3_b_30_port, s3_b_29_port, s3_b_28_port, s3_b_27_port, 
      s3_b_26_port, s3_b_25_port, s3_b_24_port, s3_b_23_port, s3_b_22_port, 
      s3_b_21_port, s3_b_20_port, s3_b_19_port, s3_b_18_port, s3_b_17_port, 
      s3_b_16_port, s3_b_15_port, s3_b_14_port, s3_b_13_port, s3_b_12_port, 
      s3_b_11_port, s3_b_10_port, s3_b_9_port, s3_b_8_port, s3_b_7_port, 
      s3_b_6_port, s3_b_5_port, s3_b_4_port, s3_b_3_port, s3_b_2_port, 
      s3_b_1_port, s3_b_0_port, s3_imm_i_ext_31_port, s3_imm_i_ext_30_port, 
      s3_imm_i_ext_29_port, s3_imm_i_ext_28_port, s3_imm_i_ext_27_port, 
      s3_imm_i_ext_26_port, s3_imm_i_ext_25_port, s3_imm_i_ext_24_port, 
      s3_imm_i_ext_23_port, s3_imm_i_ext_22_port, s3_imm_i_ext_21_port, 
      s3_imm_i_ext_20_port, s3_imm_i_ext_19_port, s3_imm_i_ext_18_port, 
      s3_imm_i_ext_17_port, s3_imm_i_ext_16_port, s3_imm_i_ext_15_port, 
      s3_imm_i_ext_14_port, s3_imm_i_ext_13_port, s3_imm_i_ext_12_port, 
      s3_imm_i_ext_11_port, s3_imm_i_ext_10_port, s3_imm_i_ext_9_port, 
      s3_imm_i_ext_8_port, s3_imm_i_ext_7_port, s3_imm_i_ext_6_port, 
      s3_imm_i_ext_5_port, s3_imm_i_ext_4_port, s3_imm_i_ext_3_port, 
      s3_imm_i_ext_2_port, s3_imm_i_ext_1_port, s3_imm_i_ext_0_port, 
      s3_rd1_addr_4_port, s3_rd1_addr_3_port, s3_rd1_addr_2_port, 
      s3_rd1_addr_1_port, s3_rd1_addr_0_port, s3_rd2_addr_4_port, 
      s3_rd2_addr_3_port, s3_rd2_addr_2_port, s3_rd2_addr_1_port, 
      s3_rd2_addr_0_port, s4_reg_b_wait, s4_a_31_port, s4_a_30_port, 
      s4_a_29_port, s4_a_28_port, s4_a_27_port, s4_a_26_port, s4_a_25_port, 
      s4_a_24_port, s4_a_23_port, s4_a_22_port, s4_a_21_port, s4_a_20_port, 
      s4_a_19_port, s4_a_18_port, s4_a_17_port, s4_a_16_port, s4_a_15_port, 
      s4_a_14_port, s4_a_13_port, s4_a_12_port, s4_a_11_port, s4_a_10_port, 
      s4_a_9_port, s4_a_8_port, s4_a_7_port, s4_a_6_port, s4_a_5_port, 
      s4_a_4_port, s4_a_3_port, s4_a_2_port, s4_a_1_port, s4_a_0_port, 
      s3_a_keep_31_port, s3_a_keep_30_port, s3_a_keep_29_port, 
      s3_a_keep_28_port, s3_a_keep_27_port, s3_a_keep_26_port, 
      s3_a_keep_25_port, s3_a_keep_24_port, s3_a_keep_23_port, 
      s3_a_keep_22_port, s3_a_keep_21_port, s3_a_keep_20_port, 
      s3_a_keep_19_port, s3_a_keep_18_port, s3_a_keep_17_port, 
      s3_a_keep_16_port, s3_a_keep_15_port, s3_a_keep_14_port, 
      s3_a_keep_13_port, s3_a_keep_12_port, s3_a_keep_11_port, 
      s3_a_keep_10_port, s3_a_keep_9_port, s3_a_keep_8_port, s3_a_keep_7_port, 
      s3_a_keep_6_port, s3_a_keep_5_port, s3_a_keep_4_port, s3_a_keep_3_port, 
      s3_a_keep_2_port, s3_a_keep_1_port, s3_a_keep_0_port, s4_reg_a_wait, 
      s4_b_31_port, s4_b_30_port, s4_b_29_port, s4_b_28_port, s4_b_27_port, 
      s4_b_26_port, s4_b_25_port, s4_b_24_port, s4_b_23_port, s4_b_22_port, 
      s4_b_21_port, s4_b_20_port, s4_b_19_port, s4_b_18_port, s4_b_17_port, 
      s4_b_16_port, s4_b_15_port, s4_b_14_port, s4_b_13_port, s4_b_12_port, 
      s4_b_11_port, s4_b_10_port, s4_b_9_port, s4_b_8_port, s4_b_7_port, 
      s4_b_6_port, s4_b_5_port, s4_b_4_port, s4_b_3_port, s4_b_2_port, 
      s4_b_1_port, s4_b_0_port, s3_b_keep_31_port, s3_b_keep_30_port, 
      s3_b_keep_29_port, s3_b_keep_28_port, s3_b_keep_27_port, 
      s3_b_keep_26_port, s3_b_keep_25_port, s3_b_keep_24_port, 
      s3_b_keep_23_port, s3_b_keep_22_port, s3_b_keep_21_port, 
      s3_b_keep_20_port, s3_b_keep_19_port, s3_b_keep_18_port, 
      s3_b_keep_17_port, s3_b_keep_16_port, s3_b_keep_15_port, 
      s3_b_keep_14_port, s3_b_keep_13_port, s3_b_keep_12_port, 
      s3_b_keep_11_port, s3_b_keep_10_port, s3_b_keep_9_port, s3_b_keep_8_port,
      s3_b_keep_7_port, s3_b_keep_6_port, s3_b_keep_5_port, s3_b_keep_4_port, 
      s3_b_keep_3_port, s3_b_keep_2_port, s3_b_keep_1_port, s3_b_keep_0_port, 
      s3_a_sel_f_en, s3_a_sel_ff_en, s3_a_sel_31_port, s3_a_sel_30_port, 
      s3_a_sel_29_port, s3_a_sel_28_port, s3_a_sel_27_port, s3_a_sel_26_port, 
      s3_a_sel_25_port, s3_a_sel_24_port, s3_a_sel_23_port, s3_a_sel_22_port, 
      s3_a_sel_21_port, s3_a_sel_20_port, s3_a_sel_19_port, s3_a_sel_18_port, 
      s3_a_sel_17_port, s3_a_sel_16_port, s3_a_sel_15_port, s3_a_sel_14_port, 
      s3_a_sel_13_port, s3_a_sel_12_port, s3_a_sel_11_port, s3_a_sel_10_port, 
      s3_a_sel_9_port, s3_a_sel_8_port, s3_a_sel_7_port, s3_a_sel_6_port, 
      s3_a_sel_5_port, s3_a_sel_4_port, s3_a_sel_3_port, s3_a_sel_2_port, 
      s3_a_sel_1_port, s3_a_sel_0_port, s3_reg_a_wait, s3_b_sel_f_en, 
      s3_b_sel_ff_en, s3_b_fwd_31_port, s3_b_fwd_30_port, s3_b_fwd_29_port, 
      s3_b_fwd_28_port, s3_b_fwd_27_port, s3_b_fwd_26_port, s3_b_fwd_25_port, 
      s3_b_fwd_24_port, s3_b_fwd_23_port, s3_b_fwd_22_port, s3_b_fwd_21_port, 
      s3_b_fwd_20_port, s3_b_fwd_19_port, s3_b_fwd_18_port, s3_b_fwd_17_port, 
      s3_b_fwd_16_port, s3_b_fwd_15_port, s3_b_fwd_14_port, s3_b_fwd_13_port, 
      s3_b_fwd_12_port, s3_b_fwd_11_port, s3_b_fwd_10_port, s3_b_fwd_9_port, 
      s3_b_fwd_8_port, s3_b_fwd_7_port, s3_b_fwd_6_port, s3_b_fwd_5_port, 
      s3_b_fwd_4_port, s3_b_fwd_3_port, s3_b_fwd_2_port, s3_b_fwd_1_port, 
      s3_b_fwd_0_port, s3_reg_b_wait, s3_b_sel_31_port, s3_b_sel_30_port, 
      s3_b_sel_29_port, s3_b_sel_28_port, s3_b_sel_27_port, s3_b_sel_26_port, 
      s3_b_sel_25_port, s3_b_sel_24_port, s3_b_sel_23_port, s3_b_sel_22_port, 
      s3_b_sel_21_port, s3_b_sel_20_port, s3_b_sel_19_port, s3_b_sel_18_port, 
      s3_b_sel_17_port, s3_b_sel_16_port, s3_b_sel_15_port, s3_b_sel_14_port, 
      s3_b_sel_13_port, s3_b_sel_12_port, s3_b_sel_11_port, s3_b_sel_10_port, 
      s3_b_sel_9_port, s3_b_sel_8_port, s3_b_sel_7_port, s3_b_sel_6_port, 
      s3_b_sel_5_port, s3_b_sel_4_port, s3_b_sel_3_port, s3_b_sel_2_port, 
      s3_b_sel_1_port, s3_b_sel_0_port, s3_alu_out_31_port, s3_alu_out_30_port,
      s3_alu_out_29_port, s3_alu_out_28_port, s3_alu_out_27_port, 
      s3_alu_out_26_port, s3_alu_out_25_port, s3_alu_out_24_port, 
      s3_alu_out_23_port, s3_alu_out_22_port, s3_alu_out_21_port, 
      s3_alu_out_20_port, s3_alu_out_19_port, s3_alu_out_18_port, 
      s3_alu_out_17_port, s3_alu_out_16_port, s3_alu_out_15_port, 
      s3_alu_out_14_port, s3_alu_out_13_port, s3_alu_out_12_port, 
      s3_alu_out_11_port, s3_alu_out_10_port, s3_alu_out_9_port, 
      s3_alu_out_8_port, s3_alu_out_7_port, s3_alu_out_6_port, 
      s3_alu_out_5_port, s3_alu_out_4_port, s3_alu_out_3_port, 
      s3_alu_out_2_port, s3_alu_out_1_port, s3_alu_out_0_port, s3_mul_sign, 
      s3_mul_out_31_port, s3_mul_out_30_port, s3_mul_out_29_port, 
      s3_mul_out_28_port, s3_mul_out_27_port, s3_mul_out_26_port, 
      s3_mul_out_25_port, s3_mul_out_24_port, s3_mul_out_23_port, 
      s3_mul_out_22_port, s3_mul_out_21_port, s3_mul_out_20_port, 
      s3_mul_out_19_port, s3_mul_out_18_port, s3_mul_out_17_port, 
      s3_mul_out_16_port, s3_mul_out_15_port, s3_mul_out_14_port, 
      s3_mul_out_13_port, s3_mul_out_12_port, s3_mul_out_11_port, 
      s3_mul_out_10_port, s3_mul_out_9_port, s3_mul_out_8_port, 
      s3_mul_out_7_port, s3_mul_out_6_port, s3_mul_out_5_port, 
      s3_mul_out_4_port, s3_mul_out_3_port, s3_mul_out_2_port, 
      s3_mul_out_1_port, s3_mul_out_0_port, s3_div_sign, s3_div_out_31_port, 
      s3_div_out_30_port, s3_div_out_29_port, s3_div_out_28_port, 
      s3_div_out_27_port, s3_div_out_26_port, s3_div_out_25_port, 
      s3_div_out_24_port, s3_div_out_23_port, s3_div_out_22_port, 
      s3_div_out_21_port, s3_div_out_20_port, s3_div_out_19_port, 
      s3_div_out_18_port, s3_div_out_17_port, s3_div_out_16_port, 
      s3_div_out_15_port, s3_div_out_14_port, s3_div_out_13_port, 
      s3_div_out_12_port, s3_div_out_11_port, s3_div_out_10_port, 
      s3_div_out_9_port, s3_div_out_8_port, s3_div_out_7_port, 
      s3_div_out_6_port, s3_div_out_5_port, s3_div_out_4_port, 
      s3_div_out_3_port, s3_div_out_2_port, s3_div_out_1_port, 
      s3_div_out_0_port, s3_exe_sel_1_port, s4_b_fwd_31_port, s4_b_fwd_30_port,
      s4_b_fwd_29_port, s4_b_fwd_28_port, s4_b_fwd_27_port, s4_b_fwd_26_port, 
      s4_b_fwd_25_port, s4_b_fwd_24_port, s4_b_fwd_23_port, s4_b_fwd_22_port, 
      s4_b_fwd_21_port, s4_b_fwd_20_port, s4_b_fwd_19_port, s4_b_fwd_18_port, 
      s4_b_fwd_17_port, s4_b_fwd_16_port, s4_b_fwd_15_port, s4_b_fwd_14_port, 
      s4_b_fwd_13_port, s4_b_fwd_12_port, s4_b_fwd_11_port, s4_b_fwd_10_port, 
      s4_b_fwd_9_port, s4_b_fwd_8_port, s4_b_fwd_7_port, s4_b_fwd_6_port, 
      s4_b_fwd_5_port, s4_b_fwd_4_port, s4_b_fwd_3_port, s4_b_fwd_2_port, 
      s4_b_fwd_1_port, s4_b_fwd_0_port, s4_rd2_addr_4_port, s4_rd2_addr_3_port,
      s4_rd2_addr_2_port, s4_rd2_addr_1_port, s4_rd2_addr_0_port, 
      s6_result_31_port, s6_result_30_port, s6_result_29_port, 
      s6_result_28_port, s6_result_27_port, s6_result_26_port, 
      s6_result_25_port, s6_result_24_port, s6_result_23_port, 
      s6_result_22_port, s6_result_21_port, s6_result_20_port, 
      s6_result_19_port, s6_result_18_port, s6_result_17_port, 
      s6_result_16_port, s6_result_15_port, s6_result_14_port, 
      s6_result_13_port, s6_result_12_port, s6_result_11_port, 
      s6_result_10_port, s6_result_9_port, s6_result_8_port, s6_result_7_port, 
      s6_result_6_port, s6_result_5_port, s6_result_4_port, s6_result_3_port, 
      s6_result_2_port, s6_result_1_port, s6_result_0_port, s6_wr_addr_4_port, 
      s6_wr_addr_3_port, s6_wr_addr_2_port, s6_wr_addr_1_port, 
      s6_wr_addr_0_port, s6_en_wb, net1283, net1284, net1287, net1288, net1290,
      net1291, net1292, net1293, net1294, n45, n48, net107975, net107976, 
      net107977, net107978, net107979, net107980, net107981, net107982, 
      net107983, net107984, net107985, net107986, net107987, net107988, 
      net107989, n43, n46, n49, n50, n51, n54, n55, n56, n57, n58, n59, n60, 
      n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75
      , n76, n77, n78, n79, n47, n52, n53, n80, n81, n82, n83, istr_addr_2_port
      , istr_addr_28_port, n86, n87, n88, n89, n90, n91, sig_sqrt_port, n93, 
      istr_addr_1_port, n95, n96, n97, n98, n99, ir_out_27_port, ir_out_28_port
      , n102, n103, n104, n105, istr_addr_0_port, n107, n108, n109, n110, n111,
      n112, n113, n114, n115, n116, n117, n118, sig_mul_port, net163711, 
      net163712 : std_logic;

begin
   istr_addr <= ( istr_addr_31_port, istr_addr_30_port, istr_addr_29_port, 
      istr_addr_28_port, istr_addr_27_port, istr_addr_26_port, 
      istr_addr_25_port, istr_addr_24_port, istr_addr_23_port, 
      istr_addr_22_port, istr_addr_21_port, istr_addr_20_port, 
      istr_addr_19_port, istr_addr_18_port, istr_addr_17_port, 
      istr_addr_16_port, istr_addr_15_port, istr_addr_14_port, 
      istr_addr_13_port, istr_addr_12_port, istr_addr_11_port, 
      istr_addr_10_port, istr_addr_9_port, istr_addr_8_port, istr_addr_7_port, 
      istr_addr_6_port, istr_addr_5_port, istr_addr_4_port, istr_addr_3_port, 
      istr_addr_2_port, istr_addr_1_port, istr_addr_0_port );
   ir_out <= ( istr_val(31), istr_val(30), istr_val(29), ir_out_28_port, 
      ir_out_27_port, istr_val(26), istr_val(25), istr_val(24), istr_val(23), 
      istr_val(22), istr_val(21), istr_val(20), istr_val(19), istr_val(18), 
      istr_val(17), istr_val(16), istr_val(15), istr_val(14), istr_val(13), 
      istr_val(12), istr_val(11), istr_val(10), istr_val(9), istr_val(8), 
      istr_val(7), istr_val(6), istr_val(5), istr_val(4), istr_val(3), 
      istr_val(2), istr_val(1), istr_val(0) );
   ld_a_out <= ( data_i_val(31), data_i_val(30), data_i_val(29), data_i_val(28)
      , data_i_val(27), data_i_val(26), data_i_val(25), data_i_val(24), 
      data_i_val(23), data_i_val(22), data_i_val(21), data_i_val(20), 
      data_i_val(19), data_i_val(18), data_i_val(17), data_i_val(16), 
      data_i_val(15), data_i_val(14), data_i_val(13), data_i_val(12), 
      data_i_val(11), data_i_val(10), data_i_val(9), data_i_val(8), 
      data_i_val(7), data_i_val(6), data_i_val(5), data_i_val(4), data_i_val(3)
      , data_i_val(2), data_i_val(1), data_i_val(0) );
   data_addr <= ( data_addr_31_port, data_addr_30_port, data_addr_29_port, 
      data_addr_28_port, data_addr_27_port, data_addr_26_port, 
      data_addr_25_port, data_addr_24_port, data_addr_23_port, 
      data_addr_22_port, data_addr_21_port, data_addr_20_port, 
      data_addr_19_port, data_addr_18_port, data_addr_17_port, 
      data_addr_16_port, data_addr_15_port, data_addr_14_port, 
      data_addr_13_port, data_addr_12_port, data_addr_11_port, 
      data_addr_10_port, data_addr_9_port, data_addr_8_port, data_addr_7_port, 
      data_addr_6_port, data_addr_5_port, data_addr_4_port, data_addr_3_port, 
      data_addr_2_port, data_addr_1_port, data_addr_0_port );
   dr_cw <= ( cw(14), cw(13), cw(12), cw(11) );
   sig_ral <= sig_ral_port;
   sig_mul <= sig_mul_port;
   sig_div <= sig_div_port;
   sig_sqrt <= sig_sqrt_port;
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   s3_jump_flag_reg : DFF_X1 port map( D => n48, CK => clk, Q => net163712, QN 
                           => n53);
   s6_en_wb_reg : DFFR_X1 port map( D => n45, CK => clk, RN => n111, Q => 
                           s6_en_wb, QN => net163711);
   U94 : NAND3_X1 port map( A1 => n49, A2 => n79, A3 => cw(6), ZN => n78);
   U95 : NAND3_X1 port map( A1 => n50, A2 => n88, A3 => ir_out_28_port, ZN => 
                           n75);
   ADD_4 : Adder_DATA_SIZE32_0 port map( cin => X_Logic0_port, a(31) => 
                           istr_addr_31_port, a(30) => istr_addr_30_port, a(29)
                           => istr_addr_29_port, a(28) => n120, a(27) => 
                           istr_addr_27_port, a(26) => istr_addr_26_port, a(25)
                           => istr_addr_25_port, a(24) => istr_addr_24_port, 
                           a(23) => istr_addr_23_port, a(22) => 
                           istr_addr_22_port, a(21) => istr_addr_21_port, a(20)
                           => istr_addr_20_port, a(19) => istr_addr_19_port, 
                           a(18) => istr_addr_18_port, a(17) => 
                           istr_addr_17_port, a(16) => istr_addr_16_port, a(15)
                           => istr_addr_15_port, a(14) => istr_addr_14_port, 
                           a(13) => istr_addr_13_port, a(12) => 
                           istr_addr_12_port, a(11) => istr_addr_11_port, a(10)
                           => istr_addr_10_port, a(9) => istr_addr_9_port, a(8)
                           => istr_addr_8_port, a(7) => istr_addr_7_port, a(6) 
                           => istr_addr_6_port, a(5) => istr_addr_5_port, a(4) 
                           => istr_addr_4_port, a(3) => istr_addr_3_port, a(2) 
                           => n121, a(1) => n122, a(0) => n123, b(31) => 
                           X_Logic0_port, b(30) => X_Logic0_port, b(29) => 
                           X_Logic0_port, b(28) => X_Logic0_port, b(27) => 
                           X_Logic0_port, b(26) => X_Logic0_port, b(25) => 
                           X_Logic0_port, b(24) => X_Logic0_port, b(23) => 
                           X_Logic0_port, b(22) => X_Logic0_port, b(21) => 
                           X_Logic0_port, b(20) => X_Logic0_port, b(19) => 
                           X_Logic0_port, b(18) => X_Logic0_port, b(17) => 
                           X_Logic0_port, b(16) => X_Logic0_port, b(15) => 
                           X_Logic0_port, b(14) => X_Logic0_port, b(13) => 
                           X_Logic0_port, b(12) => X_Logic0_port, b(11) => 
                           X_Logic0_port, b(10) => X_Logic0_port, b(9) => 
                           X_Logic0_port, b(8) => X_Logic0_port, b(7) => 
                           X_Logic0_port, b(6) => X_Logic0_port, b(5) => 
                           X_Logic0_port, b(4) => X_Logic0_port, b(3) => 
                           X_Logic0_port, b(2) => X_Logic0_port, b(1) => 
                           X_Logic0_port, b(0) => X_Logic0_port, s(31) => 
                           s1_npc_31_port, s(30) => s1_npc_30_port, s(29) => 
                           s1_npc_29_port, s(28) => s1_npc_28_port, s(27) => 
                           s1_npc_27_port, s(26) => s1_npc_26_port, s(25) => 
                           s1_npc_25_port, s(24) => s1_npc_24_port, s(23) => 
                           s1_npc_23_port, s(22) => s1_npc_22_port, s(21) => 
                           s1_npc_21_port, s(20) => s1_npc_20_port, s(19) => 
                           s1_npc_19_port, s(18) => s1_npc_18_port, s(17) => 
                           s1_npc_17_port, s(16) => s1_npc_16_port, s(15) => 
                           s1_npc_15_port, s(14) => s1_npc_14_port, s(13) => 
                           s1_npc_13_port, s(12) => s1_npc_12_port, s(11) => 
                           s1_npc_11_port, s(10) => s1_npc_10_port, s(9) => 
                           s1_npc_9_port, s(8) => s1_npc_8_port, s(7) => 
                           s1_npc_7_port, s(6) => s1_npc_6_port, s(5) => 
                           s1_npc_5_port, s(4) => s1_npc_4_port, s(3) => 
                           s1_npc_3_port, s(2) => s1_npc_2_port, s(1) => 
                           s1_npc_1_port, s(0) => s1_npc_0_port, cout => 
                           net1294);
   MUX_bpw : Mux_DATA_SIZE32_0 port map( sel => sig_bpw, din0(31) => 
                           s2_pc_sel_31_port, din0(30) => s2_pc_sel_30_port, 
                           din0(29) => s2_pc_sel_29_port, din0(28) => 
                           s2_pc_sel_28_port, din0(27) => s2_pc_sel_27_port, 
                           din0(26) => s2_pc_sel_26_port, din0(25) => 
                           s2_pc_sel_25_port, din0(24) => s2_pc_sel_24_port, 
                           din0(23) => s2_pc_sel_23_port, din0(22) => 
                           s2_pc_sel_22_port, din0(21) => s2_pc_sel_21_port, 
                           din0(20) => s2_pc_sel_20_port, din0(19) => 
                           s2_pc_sel_19_port, din0(18) => s2_pc_sel_18_port, 
                           din0(17) => s2_pc_sel_17_port, din0(16) => 
                           s2_pc_sel_16_port, din0(15) => s2_pc_sel_15_port, 
                           din0(14) => s2_pc_sel_14_port, din0(13) => 
                           s2_pc_sel_13_port, din0(12) => s2_pc_sel_12_port, 
                           din0(11) => s2_pc_sel_11_port, din0(10) => 
                           s2_pc_sel_10_port, din0(9) => s2_pc_sel_9_port, 
                           din0(8) => s2_pc_sel_8_port, din0(7) => 
                           s2_pc_sel_7_port, din0(6) => s2_pc_sel_6_port, 
                           din0(5) => s2_pc_sel_5_port, din0(4) => 
                           s2_pc_sel_4_port, din0(3) => s2_pc_sel_3_port, 
                           din0(2) => s2_pc_sel_2_port, din0(1) => 
                           s2_pc_sel_1_port, din0(0) => s2_pc_sel_0_port, 
                           din1(31) => s3_pc_notsel_31_port, din1(30) => 
                           s3_pc_notsel_30_port, din1(29) => 
                           s3_pc_notsel_29_port, din1(28) => 
                           s3_pc_notsel_28_port, din1(27) => 
                           s3_pc_notsel_27_port, din1(26) => 
                           s3_pc_notsel_26_port, din1(25) => 
                           s3_pc_notsel_25_port, din1(24) => 
                           s3_pc_notsel_24_port, din1(23) => 
                           s3_pc_notsel_23_port, din1(22) => 
                           s3_pc_notsel_22_port, din1(21) => 
                           s3_pc_notsel_21_port, din1(20) => 
                           s3_pc_notsel_20_port, din1(19) => 
                           s3_pc_notsel_19_port, din1(18) => 
                           s3_pc_notsel_18_port, din1(17) => 
                           s3_pc_notsel_17_port, din1(16) => 
                           s3_pc_notsel_16_port, din1(15) => 
                           s3_pc_notsel_15_port, din1(14) => 
                           s3_pc_notsel_14_port, din1(13) => 
                           s3_pc_notsel_13_port, din1(12) => 
                           s3_pc_notsel_12_port, din1(11) => 
                           s3_pc_notsel_11_port, din1(10) => 
                           s3_pc_notsel_10_port, din1(9) => s3_pc_notsel_9_port
                           , din1(8) => s3_pc_notsel_8_port, din1(7) => 
                           s3_pc_notsel_7_port, din1(6) => s3_pc_notsel_6_port,
                           din1(5) => s3_pc_notsel_5_port, din1(4) => 
                           s3_pc_notsel_4_port, din1(3) => s3_pc_notsel_3_port,
                           din1(2) => s3_pc_notsel_2_port, din1(1) => 
                           s3_pc_notsel_1_port, din1(0) => s3_pc_notsel_0_port,
                           dout(31) => istr_addr_31_port, dout(30) => 
                           istr_addr_30_port, dout(29) => istr_addr_29_port, 
                           dout(28) => n120, dout(27) => istr_addr_27_port, 
                           dout(26) => istr_addr_26_port, dout(25) => 
                           istr_addr_25_port, dout(24) => istr_addr_24_port, 
                           dout(23) => istr_addr_23_port, dout(22) => 
                           istr_addr_22_port, dout(21) => istr_addr_21_port, 
                           dout(20) => istr_addr_20_port, dout(19) => 
                           istr_addr_19_port, dout(18) => istr_addr_18_port, 
                           dout(17) => istr_addr_17_port, dout(16) => 
                           istr_addr_16_port, dout(15) => istr_addr_15_port, 
                           dout(14) => istr_addr_14_port, dout(13) => 
                           istr_addr_13_port, dout(12) => istr_addr_12_port, 
                           dout(11) => istr_addr_11_port, dout(10) => 
                           istr_addr_10_port, dout(9) => istr_addr_9_port, 
                           dout(8) => istr_addr_8_port, dout(7) => 
                           istr_addr_7_port, dout(6) => istr_addr_6_port, 
                           dout(5) => istr_addr_5_port, dout(4) => 
                           istr_addr_4_port, dout(3) => istr_addr_3_port, 
                           dout(2) => n121, dout(1) => n122, dout(0) => n123);
   REG_PC : Reg_DATA_SIZE32_0 port map( rst => n111, en => cw(0), clk => clk, 
                           din(31) => istr_addr_31_port, din(30) => 
                           istr_addr_30_port, din(29) => istr_addr_29_port, 
                           din(28) => istr_addr_28_port, din(27) => 
                           istr_addr_27_port, din(26) => istr_addr_26_port, 
                           din(25) => istr_addr_25_port, din(24) => 
                           istr_addr_24_port, din(23) => istr_addr_23_port, 
                           din(22) => istr_addr_22_port, din(21) => 
                           istr_addr_21_port, din(20) => istr_addr_20_port, 
                           din(19) => istr_addr_19_port, din(18) => 
                           istr_addr_18_port, din(17) => istr_addr_17_port, 
                           din(16) => istr_addr_16_port, din(15) => 
                           istr_addr_15_port, din(14) => istr_addr_14_port, 
                           din(13) => istr_addr_13_port, din(12) => 
                           istr_addr_12_port, din(11) => istr_addr_11_port, 
                           din(10) => istr_addr_10_port, din(9) => 
                           istr_addr_9_port, din(8) => istr_addr_8_port, din(7)
                           => istr_addr_7_port, din(6) => istr_addr_6_port, 
                           din(5) => istr_addr_5_port, din(4) => 
                           istr_addr_4_port, din(3) => istr_addr_3_port, din(2)
                           => istr_addr_2_port, din(1) => istr_addr_1_port, 
                           din(0) => istr_addr_0_port, dout(31) => pc_out(31), 
                           dout(30) => pc_out(30), dout(29) => pc_out(29), 
                           dout(28) => pc_out(28), dout(27) => pc_out(27), 
                           dout(26) => pc_out(26), dout(25) => pc_out(25), 
                           dout(24) => pc_out(24), dout(23) => pc_out(23), 
                           dout(22) => pc_out(22), dout(21) => pc_out(21), 
                           dout(20) => pc_out(20), dout(19) => pc_out(19), 
                           dout(18) => pc_out(18), dout(17) => pc_out(17), 
                           dout(16) => pc_out(16), dout(15) => pc_out(15), 
                           dout(14) => pc_out(14), dout(13) => pc_out(13), 
                           dout(12) => pc_out(12), dout(11) => pc_out(11), 
                           dout(10) => pc_out(10), dout(9) => pc_out(9), 
                           dout(8) => pc_out(8), dout(7) => pc_out(7), dout(6) 
                           => pc_out(6), dout(5) => pc_out(5), dout(4) => 
                           pc_out(4), dout(3) => pc_out(3), dout(2) => 
                           pc_out(2), dout(1) => pc_out(1), dout(0) => 
                           pc_out(0));
   REG_NPC : Reg_DATA_SIZE32_12 port map( rst => n111, en => cw(0), clk => clk,
                           din(31) => s1_npc_31_port, din(30) => s1_npc_30_port
                           , din(29) => s1_npc_29_port, din(28) => 
                           s1_npc_28_port, din(27) => s1_npc_27_port, din(26) 
                           => s1_npc_26_port, din(25) => s1_npc_25_port, 
                           din(24) => s1_npc_24_port, din(23) => s1_npc_23_port
                           , din(22) => s1_npc_22_port, din(21) => 
                           s1_npc_21_port, din(20) => s1_npc_20_port, din(19) 
                           => s1_npc_19_port, din(18) => s1_npc_18_port, 
                           din(17) => s1_npc_17_port, din(16) => s1_npc_16_port
                           , din(15) => s1_npc_15_port, din(14) => 
                           s1_npc_14_port, din(13) => s1_npc_13_port, din(12) 
                           => s1_npc_12_port, din(11) => s1_npc_11_port, 
                           din(10) => s1_npc_10_port, din(9) => s1_npc_9_port, 
                           din(8) => s1_npc_8_port, din(7) => s1_npc_7_port, 
                           din(6) => s1_npc_6_port, din(5) => s1_npc_5_port, 
                           din(4) => s1_npc_4_port, din(3) => s1_npc_3_port, 
                           din(2) => s1_npc_2_port, din(1) => s1_npc_1_port, 
                           din(0) => s1_npc_0_port, dout(31) => s2_npc_31_port,
                           dout(30) => s2_npc_30_port, dout(29) => 
                           s2_npc_29_port, dout(28) => s2_npc_28_port, dout(27)
                           => s2_npc_27_port, dout(26) => s2_npc_26_port, 
                           dout(25) => s2_npc_25_port, dout(24) => 
                           s2_npc_24_port, dout(23) => s2_npc_23_port, dout(22)
                           => s2_npc_22_port, dout(21) => s2_npc_21_port, 
                           dout(20) => s2_npc_20_port, dout(19) => 
                           s2_npc_19_port, dout(18) => s2_npc_18_port, dout(17)
                           => s2_npc_17_port, dout(16) => s2_npc_16_port, 
                           dout(15) => s2_npc_15_port, dout(14) => 
                           s2_npc_14_port, dout(13) => s2_npc_13_port, dout(12)
                           => s2_npc_12_port, dout(11) => s2_npc_11_port, 
                           dout(10) => s2_npc_10_port, dout(9) => s2_npc_9_port
                           , dout(8) => s2_npc_8_port, dout(7) => s2_npc_7_port
                           , dout(6) => s2_npc_6_port, dout(5) => s2_npc_5_port
                           , dout(4) => s2_npc_4_port, dout(3) => s2_npc_3_port
                           , dout(2) => s2_npc_2_port, dout(1) => s2_npc_1_port
                           , dout(0) => s2_npc_0_port);
   MUX_PC : Mux_DATA_SIZE32_9 port map( sel => cw(1), din0(31) => 
                           s2_npc_31_port, din0(30) => s2_npc_30_port, din0(29)
                           => s2_npc_29_port, din0(28) => s2_npc_28_port, 
                           din0(27) => s2_npc_27_port, din0(26) => 
                           s2_npc_26_port, din0(25) => s2_npc_25_port, din0(24)
                           => s2_npc_24_port, din0(23) => s2_npc_23_port, 
                           din0(22) => s2_npc_22_port, din0(21) => 
                           s2_npc_21_port, din0(20) => s2_npc_20_port, din0(19)
                           => s2_npc_19_port, din0(18) => s2_npc_18_port, 
                           din0(17) => s2_npc_17_port, din0(16) => 
                           s2_npc_16_port, din0(15) => s2_npc_15_port, din0(14)
                           => s2_npc_14_port, din0(13) => s2_npc_13_port, 
                           din0(12) => s2_npc_12_port, din0(11) => 
                           s2_npc_11_port, din0(10) => s2_npc_10_port, din0(9) 
                           => s2_npc_9_port, din0(8) => s2_npc_8_port, din0(7) 
                           => s2_npc_7_port, din0(6) => s2_npc_6_port, din0(5) 
                           => s2_npc_5_port, din0(4) => s2_npc_4_port, din0(3) 
                           => s2_npc_3_port, din0(2) => s2_npc_2_port, din0(1) 
                           => s2_npc_1_port, din0(0) => s2_npc_0_port, din1(31)
                           => X_Logic0_port, din1(30) => s2_jpc_30_port, 
                           din1(29) => s2_jpc_29_port, din1(28) => 
                           s2_jpc_28_port, din1(27) => s2_jpc_27_port, din1(26)
                           => s2_jpc_26_port, din1(25) => s2_jpc_25_port, 
                           din1(24) => s2_jpc_24_port, din1(23) => 
                           s2_jpc_23_port, din1(22) => s2_jpc_22_port, din1(21)
                           => s2_jpc_21_port, din1(20) => s2_jpc_20_port, 
                           din1(19) => s2_jpc_19_port, din1(18) => 
                           s2_jpc_18_port, din1(17) => s2_jpc_17_port, din1(16)
                           => s2_jpc_16_port, din1(15) => s2_jpc_15_port, 
                           din1(14) => s2_jpc_14_port, din1(13) => 
                           s2_jpc_13_port, din1(12) => s2_jpc_12_port, din1(11)
                           => s2_jpc_11_port, din1(10) => s2_jpc_10_port, 
                           din1(9) => s2_jpc_9_port, din1(8) => s2_jpc_8_port, 
                           din1(7) => s2_jpc_7_port, din1(6) => s2_jpc_6_port, 
                           din1(5) => s2_jpc_5_port, din1(4) => s2_jpc_4_port, 
                           din1(3) => s2_jpc_3_port, din1(2) => s2_jpc_2_port, 
                           din1(1) => s2_jpc_1_port, din1(0) => s2_jpc_0_port, 
                           dout(31) => s2_pc_sel_31_port, dout(30) => 
                           s2_pc_sel_30_port, dout(29) => s2_pc_sel_29_port, 
                           dout(28) => s2_pc_sel_28_port, dout(27) => 
                           s2_pc_sel_27_port, dout(26) => s2_pc_sel_26_port, 
                           dout(25) => s2_pc_sel_25_port, dout(24) => 
                           s2_pc_sel_24_port, dout(23) => s2_pc_sel_23_port, 
                           dout(22) => s2_pc_sel_22_port, dout(21) => 
                           s2_pc_sel_21_port, dout(20) => s2_pc_sel_20_port, 
                           dout(19) => s2_pc_sel_19_port, dout(18) => 
                           s2_pc_sel_18_port, dout(17) => s2_pc_sel_17_port, 
                           dout(16) => s2_pc_sel_16_port, dout(15) => 
                           s2_pc_sel_15_port, dout(14) => s2_pc_sel_14_port, 
                           dout(13) => s2_pc_sel_13_port, dout(12) => 
                           s2_pc_sel_12_port, dout(11) => s2_pc_sel_11_port, 
                           dout(10) => s2_pc_sel_10_port, dout(9) => 
                           s2_pc_sel_9_port, dout(8) => s2_pc_sel_8_port, 
                           dout(7) => s2_pc_sel_7_port, dout(6) => 
                           s2_pc_sel_6_port, dout(5) => s2_pc_sel_5_port, 
                           dout(4) => s2_pc_sel_4_port, dout(3) => 
                           s2_pc_sel_3_port, dout(2) => s2_pc_sel_2_port, 
                           dout(1) => s2_pc_sel_1_port, dout(0) => 
                           s2_pc_sel_0_port);
   MUX_NOTPC : Mux_DATA_SIZE32_8 port map( sel => n107, din0(31) => 
                           X_Logic0_port, din0(30) => s2_jpc_30_port, din0(29) 
                           => s2_jpc_29_port, din0(28) => n52, din0(27) => 
                           s2_jpc_27_port, din0(26) => s2_jpc_26_port, din0(25)
                           => s2_jpc_25_port, din0(24) => s2_jpc_24_port, 
                           din0(23) => s2_jpc_23_port, din0(22) => 
                           s2_jpc_22_port, din0(21) => s2_jpc_21_port, din0(20)
                           => s2_jpc_20_port, din0(19) => s2_jpc_19_port, 
                           din0(18) => s2_jpc_18_port, din0(17) => 
                           s2_jpc_17_port, din0(16) => s2_jpc_16_port, din0(15)
                           => s2_jpc_15_port, din0(14) => s2_jpc_14_port, 
                           din0(13) => s2_jpc_13_port, din0(12) => 
                           s2_jpc_12_port, din0(11) => s2_jpc_11_port, din0(10)
                           => s2_jpc_10_port, din0(9) => s2_jpc_9_port, din0(8)
                           => s2_jpc_8_port, din0(7) => s2_jpc_7_port, din0(6) 
                           => s2_jpc_6_port, din0(5) => s2_jpc_5_port, din0(4) 
                           => s2_jpc_4_port, din0(3) => s2_jpc_3_port, din0(2) 
                           => s2_jpc_2_port, din0(1) => s2_jpc_1_port, din0(0) 
                           => s2_jpc_0_port, din1(31) => s2_npc_31_port, 
                           din1(30) => s2_npc_30_port, din1(29) => 
                           s2_npc_29_port, din1(28) => s2_npc_28_port, din1(27)
                           => s2_npc_27_port, din1(26) => s2_npc_26_port, 
                           din1(25) => s2_npc_25_port, din1(24) => 
                           s2_npc_24_port, din1(23) => s2_npc_23_port, din1(22)
                           => s2_npc_22_port, din1(21) => s2_npc_21_port, 
                           din1(20) => s2_npc_20_port, din1(19) => 
                           s2_npc_19_port, din1(18) => s2_npc_18_port, din1(17)
                           => s2_npc_17_port, din1(16) => s2_npc_16_port, 
                           din1(15) => s2_npc_15_port, din1(14) => 
                           s2_npc_14_port, din1(13) => s2_npc_13_port, din1(12)
                           => s2_npc_12_port, din1(11) => s2_npc_11_port, 
                           din1(10) => s2_npc_10_port, din1(9) => s2_npc_9_port
                           , din1(8) => s2_npc_8_port, din1(7) => s2_npc_7_port
                           , din1(6) => s2_npc_6_port, din1(5) => s2_npc_5_port
                           , din1(4) => s2_npc_4_port, din1(3) => s2_npc_3_port
                           , din1(2) => s2_npc_2_port, din1(1) => s2_npc_1_port
                           , din1(0) => s2_npc_0_port, dout(31) => 
                           s2_pc_notsel_31_port, dout(30) => 
                           s2_pc_notsel_30_port, dout(29) => 
                           s2_pc_notsel_29_port, dout(28) => 
                           s2_pc_notsel_28_port, dout(27) => 
                           s2_pc_notsel_27_port, dout(26) => 
                           s2_pc_notsel_26_port, dout(25) => 
                           s2_pc_notsel_25_port, dout(24) => 
                           s2_pc_notsel_24_port, dout(23) => 
                           s2_pc_notsel_23_port, dout(22) => 
                           s2_pc_notsel_22_port, dout(21) => 
                           s2_pc_notsel_21_port, dout(20) => 
                           s2_pc_notsel_20_port, dout(19) => 
                           s2_pc_notsel_19_port, dout(18) => 
                           s2_pc_notsel_18_port, dout(17) => 
                           s2_pc_notsel_17_port, dout(16) => 
                           s2_pc_notsel_16_port, dout(15) => 
                           s2_pc_notsel_15_port, dout(14) => 
                           s2_pc_notsel_14_port, dout(13) => 
                           s2_pc_notsel_13_port, dout(12) => 
                           s2_pc_notsel_12_port, dout(11) => 
                           s2_pc_notsel_11_port, dout(10) => 
                           s2_pc_notsel_10_port, dout(9) => s2_pc_notsel_9_port
                           , dout(8) => s2_pc_notsel_8_port, dout(7) => 
                           s2_pc_notsel_7_port, dout(6) => s2_pc_notsel_6_port,
                           dout(5) => s2_pc_notsel_5_port, dout(4) => 
                           s2_pc_notsel_4_port, dout(3) => s2_pc_notsel_3_port,
                           dout(2) => s2_pc_notsel_2_port, dout(1) => 
                           s2_pc_notsel_1_port, dout(0) => s2_pc_notsel_0_port)
                           ;
   MUX_WB_ADDR : Mux_DATA_SIZE5 port map( sel => s2_wr_addr_sel, din0(4) => 
                           istr_val(15), din0(3) => istr_val(14), din0(2) => 
                           istr_val(13), din0(1) => istr_val(12), din0(0) => 
                           istr_val(11), din1(4) => istr_val(20), din1(3) => 
                           istr_val(19), din1(2) => istr_val(18), din1(1) => 
                           istr_val(17), din1(0) => istr_val(16), dout(4) => 
                           s2_wr_addr_4_port, dout(3) => s2_wr_addr_3_port, 
                           dout(2) => s2_wr_addr_2_port, dout(1) => 
                           s2_wr_addr_1_port, dout(0) => s2_wr_addr_0_port);
   EXT_L : Extender_SRC_SIZE16_DEST_SIZE32 port map( s => cw(5), i(15) => 
                           istr_val(15), i(14) => istr_val(14), i(13) => 
                           istr_val(13), i(12) => istr_val(12), i(11) => 
                           istr_val(11), i(10) => istr_val(10), i(9) => 
                           istr_val(9), i(8) => istr_val(8), i(7) => 
                           istr_val(7), i(6) => istr_val(6), i(5) => 
                           istr_val(5), i(4) => istr_val(4), i(3) => 
                           istr_val(3), i(2) => istr_val(2), i(1) => 
                           istr_val(1), i(0) => istr_val(0), o(31) => 
                           s2_imm_l_ext_31_port, o(30) => net107975, o(29) => 
                           net107976, o(28) => net107977, o(27) => net107978, 
                           o(26) => net107979, o(25) => net107980, o(24) => 
                           net107981, o(23) => net107982, o(22) => net107983, 
                           o(21) => net107984, o(20) => net107985, o(19) => 
                           net107986, o(18) => net107987, o(17) => net107988, 
                           o(16) => net107989, o(15) => s2_imm_l_ext_15_port, 
                           o(14) => s2_imm_l_ext_14_port, o(13) => 
                           s2_imm_l_ext_13_port, o(12) => s2_imm_l_ext_12_port,
                           o(11) => s2_imm_l_ext_11_port, o(10) => 
                           s2_imm_l_ext_10_port, o(9) => s2_imm_l_ext_9_port, 
                           o(8) => s2_imm_l_ext_8_port, o(7) => 
                           s2_imm_l_ext_7_port, o(6) => s2_imm_l_ext_6_port, 
                           o(5) => s2_imm_l_ext_5_port, o(4) => 
                           s2_imm_l_ext_4_port, o(3) => s2_imm_l_ext_3_port, 
                           o(2) => s2_imm_l_ext_2_port, o(1) => 
                           s2_imm_l_ext_1_port, o(0) => s2_imm_l_ext_0_port);
   EXT_J : Extender_SRC_SIZE26_DEST_SIZE32 port map( s => X_Logic1_port, i(25) 
                           => istr_val(25), i(24) => istr_val(24), i(23) => 
                           istr_val(23), i(22) => istr_val(22), i(21) => 
                           istr_val(21), i(20) => istr_val(20), i(19) => 
                           istr_val(19), i(18) => istr_val(18), i(17) => 
                           istr_val(17), i(16) => istr_val(16), i(15) => 
                           istr_val(15), i(14) => istr_val(14), i(13) => 
                           istr_val(13), i(12) => istr_val(12), i(11) => 
                           istr_val(11), i(10) => istr_val(10), i(9) => 
                           istr_val(9), i(8) => istr_val(8), i(7) => 
                           istr_val(7), i(6) => istr_val(6), i(5) => 
                           istr_val(5), i(4) => istr_val(4), i(3) => 
                           istr_val(3), i(2) => istr_val(2), i(1) => 
                           istr_val(1), i(0) => istr_val(0), o(31) => 
                           s2_imm_j_ext_31_port, o(30) => s2_imm_j_ext_30_port,
                           o(29) => s2_imm_j_ext_29_port, o(28) => 
                           s2_imm_j_ext_28_port, o(27) => s2_imm_j_ext_27_port,
                           o(26) => s2_imm_j_ext_26_port, o(25) => 
                           s2_imm_j_ext_25_port, o(24) => s2_imm_j_ext_24_port,
                           o(23) => s2_imm_j_ext_23_port, o(22) => 
                           s2_imm_j_ext_22_port, o(21) => s2_imm_j_ext_21_port,
                           o(20) => s2_imm_j_ext_20_port, o(19) => 
                           s2_imm_j_ext_19_port, o(18) => s2_imm_j_ext_18_port,
                           o(17) => s2_imm_j_ext_17_port, o(16) => 
                           s2_imm_j_ext_16_port, o(15) => s2_imm_j_ext_15_port,
                           o(14) => s2_imm_j_ext_14_port, o(13) => 
                           s2_imm_j_ext_13_port, o(12) => s2_imm_j_ext_12_port,
                           o(11) => s2_imm_j_ext_11_port, o(10) => 
                           s2_imm_j_ext_10_port, o(9) => s2_imm_j_ext_9_port, 
                           o(8) => s2_imm_j_ext_8_port, o(7) => 
                           s2_imm_j_ext_7_port, o(6) => s2_imm_j_ext_6_port, 
                           o(5) => s2_imm_j_ext_5_port, o(4) => 
                           s2_imm_j_ext_4_port, o(3) => s2_imm_j_ext_3_port, 
                           o(2) => s2_imm_j_ext_2_port, o(1) => 
                           s2_imm_j_ext_1_port, o(0) => s2_imm_j_ext_0_port);
   RF0 : RegisterFile_DATA_SIZE32_REG_NUM32 port map( clk => clk, rst => n110, 
                           en => s2_rf_en, rd1_en => cw(6), rd2_en => cw(6), 
                           wr_en => cw(19), link_en => cw(4), rd1_addr(4) => 
                           istr_val(25), rd1_addr(3) => istr_val(24), 
                           rd1_addr(2) => istr_val(23), rd1_addr(1) => 
                           istr_val(22), rd1_addr(0) => istr_val(21), 
                           rd2_addr(4) => istr_val(20), rd2_addr(3) => 
                           istr_val(19), rd2_addr(2) => istr_val(18), 
                           rd2_addr(1) => istr_val(17), rd2_addr(0) => 
                           istr_val(16), wr_addr(4) => s5_wr_addr_4_port, 
                           wr_addr(3) => s5_wr_addr_3_port, wr_addr(2) => 
                           s5_wr_addr_2_port, wr_addr(1) => s5_wr_addr_1_port, 
                           wr_addr(0) => s5_wr_addr_0_port, d_out1(31) => 
                           s2_a_31_port, d_out1(30) => s2_a_30_port, d_out1(29)
                           => s2_a_29_port, d_out1(28) => s2_a_28_port, 
                           d_out1(27) => s2_a_27_port, d_out1(26) => 
                           s2_a_26_port, d_out1(25) => s2_a_25_port, d_out1(24)
                           => s2_a_24_port, d_out1(23) => s2_a_23_port, 
                           d_out1(22) => s2_a_22_port, d_out1(21) => 
                           s2_a_21_port, d_out1(20) => s2_a_20_port, d_out1(19)
                           => s2_a_19_port, d_out1(18) => s2_a_18_port, 
                           d_out1(17) => s2_a_17_port, d_out1(16) => 
                           s2_a_16_port, d_out1(15) => s2_a_15_port, d_out1(14)
                           => s2_a_14_port, d_out1(13) => s2_a_13_port, 
                           d_out1(12) => s2_a_12_port, d_out1(11) => 
                           s2_a_11_port, d_out1(10) => s2_a_10_port, d_out1(9) 
                           => s2_a_9_port, d_out1(8) => s2_a_8_port, d_out1(7) 
                           => s2_a_7_port, d_out1(6) => s2_a_6_port, d_out1(5) 
                           => s2_a_5_port, d_out1(4) => s2_a_4_port, d_out1(3) 
                           => s2_a_3_port, d_out1(2) => s2_a_2_port, d_out1(1) 
                           => s2_a_1_port, d_out1(0) => s2_a_0_port, d_out2(31)
                           => s2_b_31_port, d_out2(30) => s2_b_30_port, 
                           d_out2(29) => s2_b_29_port, d_out2(28) => 
                           s2_b_28_port, d_out2(27) => s2_b_27_port, d_out2(26)
                           => s2_b_26_port, d_out2(25) => s2_b_25_port, 
                           d_out2(24) => s2_b_24_port, d_out2(23) => 
                           s2_b_23_port, d_out2(22) => s2_b_22_port, d_out2(21)
                           => s2_b_21_port, d_out2(20) => s2_b_20_port, 
                           d_out2(19) => s2_b_19_port, d_out2(18) => 
                           s2_b_18_port, d_out2(17) => s2_b_17_port, d_out2(16)
                           => s2_b_16_port, d_out2(15) => s2_b_15_port, 
                           d_out2(14) => s2_b_14_port, d_out2(13) => 
                           s2_b_13_port, d_out2(12) => s2_b_12_port, d_out2(11)
                           => s2_b_11_port, d_out2(10) => s2_b_10_port, 
                           d_out2(9) => s2_b_9_port, d_out2(8) => s2_b_8_port, 
                           d_out2(7) => s2_b_7_port, d_out2(6) => s2_b_6_port, 
                           d_out2(5) => s2_b_5_port, d_out2(4) => s2_b_4_port, 
                           d_out2(3) => s2_b_3_port, d_out2(2) => s2_b_2_port, 
                           d_out2(1) => s2_b_1_port, d_out2(0) => s2_b_0_port, 
                           d_in(31) => s5_result_31_port, d_in(30) => 
                           s5_result_30_port, d_in(29) => s5_result_29_port, 
                           d_in(28) => s5_result_28_port, d_in(27) => 
                           s5_result_27_port, d_in(26) => s5_result_26_port, 
                           d_in(25) => s5_result_25_port, d_in(24) => 
                           s5_result_24_port, d_in(23) => s5_result_23_port, 
                           d_in(22) => s5_result_22_port, d_in(21) => 
                           s5_result_21_port, d_in(20) => s5_result_20_port, 
                           d_in(19) => s5_result_19_port, d_in(18) => 
                           s5_result_18_port, d_in(17) => s5_result_17_port, 
                           d_in(16) => s5_result_16_port, d_in(15) => 
                           s5_result_15_port, d_in(14) => s5_result_14_port, 
                           d_in(13) => s5_result_13_port, d_in(12) => 
                           s5_result_12_port, d_in(11) => s5_result_11_port, 
                           d_in(10) => s5_result_10_port, d_in(9) => 
                           s5_result_9_port, d_in(8) => s5_result_8_port, 
                           d_in(7) => s5_result_7_port, d_in(6) => 
                           s5_result_6_port, d_in(5) => s5_result_5_port, 
                           d_in(4) => s5_result_4_port, d_in(3) => 
                           s5_result_3_port, d_in(2) => s5_result_2_port, 
                           d_in(1) => s5_result_1_port, d_in(0) => 
                           s5_result_0_port, d_link(31) => s2_npc_31_port, 
                           d_link(30) => s2_npc_30_port, d_link(29) => 
                           s2_npc_29_port, d_link(28) => s2_npc_28_port, 
                           d_link(27) => s2_npc_27_port, d_link(26) => 
                           s2_npc_26_port, d_link(25) => s2_npc_25_port, 
                           d_link(24) => s2_npc_24_port, d_link(23) => 
                           s2_npc_23_port, d_link(22) => s2_npc_22_port, 
                           d_link(21) => s2_npc_21_port, d_link(20) => 
                           s2_npc_20_port, d_link(19) => s2_npc_19_port, 
                           d_link(18) => s2_npc_18_port, d_link(17) => 
                           s2_npc_17_port, d_link(16) => s2_npc_16_port, 
                           d_link(15) => s2_npc_15_port, d_link(14) => 
                           s2_npc_14_port, d_link(13) => s2_npc_13_port, 
                           d_link(12) => s2_npc_12_port, d_link(11) => 
                           s2_npc_11_port, d_link(10) => s2_npc_10_port, 
                           d_link(9) => s2_npc_9_port, d_link(8) => 
                           s2_npc_8_port, d_link(7) => s2_npc_7_port, d_link(6)
                           => s2_npc_6_port, d_link(5) => s2_npc_5_port, 
                           d_link(4) => s2_npc_4_port, d_link(3) => 
                           s2_npc_3_port, d_link(2) => s2_npc_2_port, d_link(1)
                           => s2_npc_1_port, d_link(0) => s2_npc_0_port);
   MUX_JPC0 : Mux_DATA_SIZE32_7 port map( sel => cw(2), din0(31) => 
                           s2_imm_i_ext_31_port, din0(30) => 
                           s2_imm_i_ext_30_port, din0(29) => 
                           s2_imm_i_ext_29_port, din0(28) => 
                           s2_imm_i_ext_28_port, din0(27) => 
                           s2_imm_i_ext_27_port, din0(26) => 
                           s2_imm_i_ext_26_port, din0(25) => 
                           s2_imm_i_ext_25_port, din0(24) => 
                           s2_imm_i_ext_24_port, din0(23) => 
                           s2_imm_i_ext_23_port, din0(22) => 
                           s2_imm_i_ext_22_port, din0(21) => 
                           s2_imm_i_ext_21_port, din0(20) => 
                           s2_imm_i_ext_20_port, din0(19) => 
                           s2_imm_i_ext_19_port, din0(18) => 
                           s2_imm_i_ext_18_port, din0(17) => 
                           s2_imm_i_ext_17_port, din0(16) => 
                           s2_imm_i_ext_16_port, din0(15) => 
                           s2_imm_i_ext_15_port, din0(14) => 
                           s2_imm_i_ext_14_port, din0(13) => 
                           s2_imm_i_ext_13_port, din0(12) => 
                           s2_imm_i_ext_12_port, din0(11) => 
                           s2_imm_i_ext_11_port, din0(10) => 
                           s2_imm_i_ext_10_port, din0(9) => s2_imm_i_ext_9_port
                           , din0(8) => s2_imm_i_ext_8_port, din0(7) => 
                           s2_imm_i_ext_7_port, din0(6) => s2_imm_i_ext_6_port,
                           din0(5) => s2_imm_i_ext_5_port, din0(4) => 
                           s2_imm_i_ext_4_port, din0(3) => s2_imm_i_ext_3_port,
                           din0(2) => s2_imm_i_ext_2_port, din0(1) => 
                           s2_imm_i_ext_1_port, din0(0) => s2_imm_i_ext_0_port,
                           din1(31) => s2_imm_j_ext_31_port, din1(30) => 
                           s2_imm_j_ext_30_port, din1(29) => 
                           s2_imm_j_ext_29_port, din1(28) => 
                           s2_imm_j_ext_28_port, din1(27) => 
                           s2_imm_j_ext_27_port, din1(26) => 
                           s2_imm_j_ext_26_port, din1(25) => 
                           s2_imm_j_ext_25_port, din1(24) => 
                           s2_imm_j_ext_24_port, din1(23) => 
                           s2_imm_j_ext_23_port, din1(22) => 
                           s2_imm_j_ext_22_port, din1(21) => 
                           s2_imm_j_ext_21_port, din1(20) => 
                           s2_imm_j_ext_20_port, din1(19) => 
                           s2_imm_j_ext_19_port, din1(18) => 
                           s2_imm_j_ext_18_port, din1(17) => 
                           s2_imm_j_ext_17_port, din1(16) => 
                           s2_imm_j_ext_16_port, din1(15) => 
                           s2_imm_j_ext_15_port, din1(14) => 
                           s2_imm_j_ext_14_port, din1(13) => 
                           s2_imm_j_ext_13_port, din1(12) => 
                           s2_imm_j_ext_12_port, din1(11) => 
                           s2_imm_j_ext_11_port, din1(10) => 
                           s2_imm_j_ext_10_port, din1(9) => s2_imm_j_ext_9_port
                           , din1(8) => s2_imm_j_ext_8_port, din1(7) => 
                           s2_imm_j_ext_7_port, din1(6) => s2_imm_j_ext_6_port,
                           din1(5) => s2_imm_j_ext_5_port, din1(4) => 
                           s2_imm_j_ext_4_port, din1(3) => s2_imm_j_ext_3_port,
                           din1(2) => s2_imm_j_ext_2_port, din1(1) => 
                           s2_imm_j_ext_1_port, din1(0) => s2_imm_j_ext_0_port,
                           dout(31) => s2_jump_addr_imm_31_port, dout(30) => 
                           s2_jump_addr_imm_30_port, dout(29) => 
                           s2_jump_addr_imm_29_port, dout(28) => 
                           s2_jump_addr_imm_28_port, dout(27) => 
                           s2_jump_addr_imm_27_port, dout(26) => 
                           s2_jump_addr_imm_26_port, dout(25) => 
                           s2_jump_addr_imm_25_port, dout(24) => 
                           s2_jump_addr_imm_24_port, dout(23) => 
                           s2_jump_addr_imm_23_port, dout(22) => 
                           s2_jump_addr_imm_22_port, dout(21) => 
                           s2_jump_addr_imm_21_port, dout(20) => 
                           s2_jump_addr_imm_20_port, dout(19) => 
                           s2_jump_addr_imm_19_port, dout(18) => 
                           s2_jump_addr_imm_18_port, dout(17) => 
                           s2_jump_addr_imm_17_port, dout(16) => 
                           s2_jump_addr_imm_16_port, dout(15) => 
                           s2_jump_addr_imm_15_port, dout(14) => 
                           s2_jump_addr_imm_14_port, dout(13) => 
                           s2_jump_addr_imm_13_port, dout(12) => 
                           s2_jump_addr_imm_12_port, dout(11) => 
                           s2_jump_addr_imm_11_port, dout(10) => 
                           s2_jump_addr_imm_10_port, dout(9) => 
                           s2_jump_addr_imm_9_port, dout(8) => 
                           s2_jump_addr_imm_8_port, dout(7) => 
                           s2_jump_addr_imm_7_port, dout(6) => 
                           s2_jump_addr_imm_6_port, dout(5) => 
                           s2_jump_addr_imm_5_port, dout(4) => 
                           s2_jump_addr_imm_4_port, dout(3) => 
                           s2_jump_addr_imm_3_port, dout(2) => 
                           s2_jump_addr_imm_2_port, dout(1) => 
                           s2_jump_addr_imm_1_port, dout(0) => 
                           s2_jump_addr_imm_0_port);
   ADDER_ADDR : Adder_DATA_SIZE32_7 port map( cin => X_Logic0_port, a(31) => 
                           s2_npc_31_port, a(30) => s2_npc_30_port, a(29) => 
                           s2_npc_29_port, a(28) => s2_npc_28_port, a(27) => 
                           s2_npc_27_port, a(26) => s2_npc_26_port, a(25) => 
                           s2_npc_25_port, a(24) => s2_npc_24_port, a(23) => 
                           s2_npc_23_port, a(22) => s2_npc_22_port, a(21) => 
                           s2_npc_21_port, a(20) => s2_npc_20_port, a(19) => 
                           s2_npc_19_port, a(18) => s2_npc_18_port, a(17) => 
                           s2_npc_17_port, a(16) => s2_npc_16_port, a(15) => 
                           s2_npc_15_port, a(14) => s2_npc_14_port, a(13) => 
                           s2_npc_13_port, a(12) => s2_npc_12_port, a(11) => 
                           s2_npc_11_port, a(10) => s2_npc_10_port, a(9) => 
                           s2_npc_9_port, a(8) => s2_npc_8_port, a(7) => 
                           s2_npc_7_port, a(6) => s2_npc_6_port, a(5) => 
                           s2_npc_5_port, a(4) => s2_npc_4_port, a(3) => 
                           s2_npc_3_port, a(2) => s2_npc_2_port, a(1) => 
                           s2_npc_1_port, a(0) => s2_npc_0_port, b(31) => 
                           s2_jump_addr_imm_31_port, b(30) => 
                           s2_jump_addr_imm_30_port, b(29) => 
                           s2_jump_addr_imm_29_port, b(28) => 
                           s2_jump_addr_imm_28_port, b(27) => 
                           s2_jump_addr_imm_27_port, b(26) => 
                           s2_jump_addr_imm_26_port, b(25) => 
                           s2_jump_addr_imm_25_port, b(24) => 
                           s2_jump_addr_imm_24_port, b(23) => 
                           s2_jump_addr_imm_23_port, b(22) => 
                           s2_jump_addr_imm_22_port, b(21) => 
                           s2_jump_addr_imm_21_port, b(20) => 
                           s2_jump_addr_imm_20_port, b(19) => 
                           s2_jump_addr_imm_19_port, b(18) => 
                           s2_jump_addr_imm_18_port, b(17) => 
                           s2_jump_addr_imm_17_port, b(16) => 
                           s2_jump_addr_imm_16_port, b(15) => 
                           s2_jump_addr_imm_15_port, b(14) => 
                           s2_jump_addr_imm_14_port, b(13) => 
                           s2_jump_addr_imm_13_port, b(12) => 
                           s2_jump_addr_imm_12_port, b(11) => 
                           s2_jump_addr_imm_11_port, b(10) => 
                           s2_jump_addr_imm_10_port, b(9) => 
                           s2_jump_addr_imm_9_port, b(8) => 
                           s2_jump_addr_imm_8_port, b(7) => 
                           s2_jump_addr_imm_7_port, b(6) => 
                           s2_jump_addr_imm_6_port, b(5) => 
                           s2_jump_addr_imm_5_port, b(4) => 
                           s2_jump_addr_imm_4_port, b(3) => 
                           s2_jump_addr_imm_3_port, b(2) => 
                           s2_jump_addr_imm_2_port, b(1) => 
                           s2_jump_addr_imm_1_port, b(0) => 
                           s2_jump_addr_imm_0_port, s(31) => 
                           s2_jump_addr_rel_31_port, s(30) => 
                           s2_jump_addr_rel_30_port, s(29) => 
                           s2_jump_addr_rel_29_port, s(28) => 
                           s2_jump_addr_rel_28_port, s(27) => 
                           s2_jump_addr_rel_27_port, s(26) => 
                           s2_jump_addr_rel_26_port, s(25) => 
                           s2_jump_addr_rel_25_port, s(24) => 
                           s2_jump_addr_rel_24_port, s(23) => 
                           s2_jump_addr_rel_23_port, s(22) => 
                           s2_jump_addr_rel_22_port, s(21) => 
                           s2_jump_addr_rel_21_port, s(20) => 
                           s2_jump_addr_rel_20_port, s(19) => 
                           s2_jump_addr_rel_19_port, s(18) => 
                           s2_jump_addr_rel_18_port, s(17) => 
                           s2_jump_addr_rel_17_port, s(16) => 
                           s2_jump_addr_rel_16_port, s(15) => 
                           s2_jump_addr_rel_15_port, s(14) => 
                           s2_jump_addr_rel_14_port, s(13) => 
                           s2_jump_addr_rel_13_port, s(12) => 
                           s2_jump_addr_rel_12_port, s(11) => 
                           s2_jump_addr_rel_11_port, s(10) => 
                           s2_jump_addr_rel_10_port, s(9) => 
                           s2_jump_addr_rel_9_port, s(8) => 
                           s2_jump_addr_rel_8_port, s(7) => 
                           s2_jump_addr_rel_7_port, s(6) => 
                           s2_jump_addr_rel_6_port, s(5) => 
                           s2_jump_addr_rel_5_port, s(4) => 
                           s2_jump_addr_rel_4_port, s(3) => 
                           s2_jump_addr_rel_3_port, s(2) => 
                           s2_jump_addr_rel_2_port, s(1) => 
                           s2_jump_addr_rel_1_port, s(0) => 
                           s2_jump_addr_rel_0_port, cout => net1293);
   MUX_JPC1 : Mux_DATA_SIZE32_6 port map( sel => cw(3), din0(31) => 
                           s2_jump_addr_rel_31_port, din0(30) => 
                           s2_jump_addr_rel_30_port, din0(29) => 
                           s2_jump_addr_rel_29_port, din0(28) => 
                           s2_jump_addr_rel_28_port, din0(27) => 
                           s2_jump_addr_rel_27_port, din0(26) => 
                           s2_jump_addr_rel_26_port, din0(25) => 
                           s2_jump_addr_rel_25_port, din0(24) => 
                           s2_jump_addr_rel_24_port, din0(23) => 
                           s2_jump_addr_rel_23_port, din0(22) => 
                           s2_jump_addr_rel_22_port, din0(21) => 
                           s2_jump_addr_rel_21_port, din0(20) => 
                           s2_jump_addr_rel_20_port, din0(19) => 
                           s2_jump_addr_rel_19_port, din0(18) => 
                           s2_jump_addr_rel_18_port, din0(17) => 
                           s2_jump_addr_rel_17_port, din0(16) => 
                           s2_jump_addr_rel_16_port, din0(15) => 
                           s2_jump_addr_rel_15_port, din0(14) => 
                           s2_jump_addr_rel_14_port, din0(13) => 
                           s2_jump_addr_rel_13_port, din0(12) => 
                           s2_jump_addr_rel_12_port, din0(11) => 
                           s2_jump_addr_rel_11_port, din0(10) => 
                           s2_jump_addr_rel_10_port, din0(9) => 
                           s2_jump_addr_rel_9_port, din0(8) => 
                           s2_jump_addr_rel_8_port, din0(7) => 
                           s2_jump_addr_rel_7_port, din0(6) => 
                           s2_jump_addr_rel_6_port, din0(5) => 
                           s2_jump_addr_rel_5_port, din0(4) => 
                           s2_jump_addr_rel_4_port, din0(3) => 
                           s2_jump_addr_rel_3_port, din0(2) => 
                           s2_jump_addr_rel_2_port, din0(1) => 
                           s2_jump_addr_rel_1_port, din0(0) => 
                           s2_jump_addr_rel_0_port, din1(31) => 
                           s2_jump_addr_reg_31_port, din1(30) => 
                           s2_jump_addr_reg_30_port, din1(29) => 
                           s2_jump_addr_reg_29_port, din1(28) => 
                           s2_jump_addr_reg_28_port, din1(27) => 
                           s2_jump_addr_reg_27_port, din1(26) => 
                           s2_jump_addr_reg_26_port, din1(25) => 
                           s2_jump_addr_reg_25_port, din1(24) => 
                           s2_jump_addr_reg_24_port, din1(23) => 
                           s2_jump_addr_reg_23_port, din1(22) => 
                           s2_jump_addr_reg_22_port, din1(21) => 
                           s2_jump_addr_reg_21_port, din1(20) => 
                           s2_jump_addr_reg_20_port, din1(19) => 
                           s2_jump_addr_reg_19_port, din1(18) => 
                           s2_jump_addr_reg_18_port, din1(17) => 
                           s2_jump_addr_reg_17_port, din1(16) => 
                           s2_jump_addr_reg_16_port, din1(15) => 
                           s2_jump_addr_reg_15_port, din1(14) => 
                           s2_jump_addr_reg_14_port, din1(13) => 
                           s2_jump_addr_reg_13_port, din1(12) => 
                           s2_jump_addr_reg_12_port, din1(11) => 
                           s2_jump_addr_reg_11_port, din1(10) => 
                           s2_jump_addr_reg_10_port, din1(9) => 
                           s2_jump_addr_reg_9_port, din1(8) => 
                           s2_jump_addr_reg_8_port, din1(7) => 
                           s2_jump_addr_reg_7_port, din1(6) => 
                           s2_jump_addr_reg_6_port, din1(5) => 
                           s2_jump_addr_reg_5_port, din1(4) => 
                           s2_jump_addr_reg_4_port, din1(3) => 
                           s2_jump_addr_reg_3_port, din1(2) => 
                           s2_jump_addr_reg_2_port, din1(1) => 
                           s2_jump_addr_reg_1_port, din1(0) => 
                           s2_jump_addr_reg_0_port, dout(31) => net1292, 
                           dout(30) => s2_jpc_30_port, dout(29) => 
                           s2_jpc_29_port, dout(28) => s2_jpc_28_port, dout(27)
                           => s2_jpc_27_port, dout(26) => s2_jpc_26_port, 
                           dout(25) => s2_jpc_25_port, dout(24) => 
                           s2_jpc_24_port, dout(23) => s2_jpc_23_port, dout(22)
                           => s2_jpc_22_port, dout(21) => s2_jpc_21_port, 
                           dout(20) => s2_jpc_20_port, dout(19) => 
                           s2_jpc_19_port, dout(18) => s2_jpc_18_port, dout(17)
                           => s2_jpc_17_port, dout(16) => s2_jpc_16_port, 
                           dout(15) => s2_jpc_15_port, dout(14) => 
                           s2_jpc_14_port, dout(13) => s2_jpc_13_port, dout(12)
                           => s2_jpc_12_port, dout(11) => s2_jpc_11_port, 
                           dout(10) => s2_jpc_10_port, dout(9) => s2_jpc_9_port
                           , dout(8) => s2_jpc_8_port, dout(7) => s2_jpc_7_port
                           , dout(6) => s2_jpc_6_port, dout(5) => s2_jpc_5_port
                           , dout(4) => s2_jpc_4_port, dout(3) => s2_jpc_3_port
                           , dout(2) => s2_jpc_2_port, dout(1) => s2_jpc_1_port
                           , dout(0) => s2_jpc_0_port);
   FWDMUX_2AB : FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_0 port map( reg_c(31) => 
                           s2_a_31_port, reg_c(30) => s2_a_30_port, reg_c(29) 
                           => s2_a_29_port, reg_c(28) => s2_a_28_port, 
                           reg_c(27) => s2_a_27_port, reg_c(26) => s2_a_26_port
                           , reg_c(25) => s2_a_25_port, reg_c(24) => 
                           s2_a_24_port, reg_c(23) => s2_a_23_port, reg_c(22) 
                           => s2_a_22_port, reg_c(21) => s2_a_21_port, 
                           reg_c(20) => s2_a_20_port, reg_c(19) => s2_a_19_port
                           , reg_c(18) => s2_a_18_port, reg_c(17) => 
                           s2_a_17_port, reg_c(16) => s2_a_16_port, reg_c(15) 
                           => s2_a_15_port, reg_c(14) => s2_a_14_port, 
                           reg_c(13) => s2_a_13_port, reg_c(12) => s2_a_12_port
                           , reg_c(11) => s2_a_11_port, reg_c(10) => 
                           s2_a_10_port, reg_c(9) => s2_a_9_port, reg_c(8) => 
                           s2_a_8_port, reg_c(7) => s2_a_7_port, reg_c(6) => 
                           s2_a_6_port, reg_c(5) => s2_a_5_port, reg_c(4) => 
                           s2_a_4_port, reg_c(3) => s2_a_3_port, reg_c(2) => 
                           s2_a_2_port, reg_c(1) => s2_a_1_port, reg_c(0) => 
                           s2_a_0_port, reg_f(31) => n83, reg_f(30) => n80, 
                           reg_f(29) => n81, reg_f(28) => n82, reg_f(27) => 
                           s3_exe_out_27_port, reg_f(26) => s3_exe_out_26_port,
                           reg_f(25) => s3_exe_out_25_port, reg_f(24) => 
                           s3_exe_out_24_port, reg_f(23) => s3_exe_out_23_port,
                           reg_f(22) => s3_exe_out_22_port, reg_f(21) => 
                           s3_exe_out_21_port, reg_f(20) => s3_exe_out_20_port,
                           reg_f(19) => s3_exe_out_19_port, reg_f(18) => 
                           s3_exe_out_18_port, reg_f(17) => s3_exe_out_17_port,
                           reg_f(16) => s3_exe_out_16_port, reg_f(15) => 
                           s3_exe_out_15_port, reg_f(14) => s3_exe_out_14_port,
                           reg_f(13) => s3_exe_out_13_port, reg_f(12) => 
                           s3_exe_out_12_port, reg_f(11) => s3_exe_out_11_port,
                           reg_f(10) => s3_exe_out_10_port, reg_f(9) => 
                           s3_exe_out_9_port, reg_f(8) => s3_exe_out_8_port, 
                           reg_f(7) => s3_exe_out_7_port, reg_f(6) => 
                           s3_exe_out_6_port, reg_f(5) => s3_exe_out_5_port, 
                           reg_f(4) => s3_exe_out_4_port, reg_f(3) => 
                           s3_exe_out_3_port, reg_f(2) => s3_exe_out_2_port, 
                           reg_f(1) => s3_exe_out_1_port, reg_f(0) => n105, 
                           reg_ff(31) => s4_result_31_port, reg_ff(30) => 
                           s4_result_30_port, reg_ff(29) => s4_result_29_port, 
                           reg_ff(28) => s4_result_28_port, reg_ff(27) => 
                           s4_result_27_port, reg_ff(26) => s4_result_26_port, 
                           reg_ff(25) => s4_result_25_port, reg_ff(24) => 
                           s4_result_24_port, reg_ff(23) => s4_result_23_port, 
                           reg_ff(22) => s4_result_22_port, reg_ff(21) => 
                           s4_result_21_port, reg_ff(20) => s4_result_20_port, 
                           reg_ff(19) => s4_result_19_port, reg_ff(18) => 
                           s4_result_18_port, reg_ff(17) => s4_result_17_port, 
                           reg_ff(16) => s4_result_16_port, reg_ff(15) => 
                           s4_result_15_port, reg_ff(14) => s4_result_14_port, 
                           reg_ff(13) => s4_result_13_port, reg_ff(12) => 
                           s4_result_12_port, reg_ff(11) => s4_result_11_port, 
                           reg_ff(10) => s4_result_10_port, reg_ff(9) => 
                           s4_result_9_port, reg_ff(8) => s4_result_8_port, 
                           reg_ff(7) => s4_result_7_port, reg_ff(6) => 
                           s4_result_6_port, reg_ff(5) => s4_result_5_port, 
                           reg_ff(4) => s4_result_4_port, reg_ff(3) => 
                           s4_result_3_port, reg_ff(2) => s4_result_2_port, 
                           reg_ff(1) => s4_result_1_port, reg_ff(0) => 
                           s4_result_0_port, addr_c(4) => istr_val(25), 
                           addr_c(3) => istr_val(24), addr_c(2) => istr_val(23)
                           , addr_c(1) => istr_val(22), addr_c(0) => 
                           istr_val(21), addr_f(4) => s3_wr_addr_4_port, 
                           addr_f(3) => s3_wr_addr_3_port, addr_f(2) => 
                           s3_wr_addr_2_port, addr_f(1) => s3_wr_addr_1_port, 
                           addr_f(0) => s3_wr_addr_0_port, addr_ff(4) => 
                           s4_wr_addr_4_port, addr_ff(3) => s4_wr_addr_3_port, 
                           addr_ff(2) => s4_wr_addr_2_port, addr_ff(1) => 
                           s4_wr_addr_1_port, addr_ff(0) => s4_wr_addr_0_port, 
                           valid_f => s2_a_f_b_en, valid_ff => s2_a_ff_b_en, 
                           dirty_f => cw(8), dirty_ff => X_Logic0_port, en => 
                           X_Logic1_port, output(31) => reg_a_out(31), 
                           output(30) => reg_a_out(30), output(29) => 
                           reg_a_out(29), output(28) => reg_a_out(28), 
                           output(27) => reg_a_out(27), output(26) => 
                           reg_a_out(26), output(25) => reg_a_out(25), 
                           output(24) => reg_a_out(24), output(23) => 
                           reg_a_out(23), output(22) => reg_a_out(22), 
                           output(21) => reg_a_out(21), output(20) => 
                           reg_a_out(20), output(19) => reg_a_out(19), 
                           output(18) => reg_a_out(18), output(17) => 
                           reg_a_out(17), output(16) => reg_a_out(16), 
                           output(15) => reg_a_out(15), output(14) => 
                           reg_a_out(14), output(13) => reg_a_out(13), 
                           output(12) => reg_a_out(12), output(11) => 
                           reg_a_out(11), output(10) => reg_a_out(10), 
                           output(9) => reg_a_out(9), output(8) => reg_a_out(8)
                           , output(7) => reg_a_out(7), output(6) => 
                           reg_a_out(6), output(5) => reg_a_out(5), output(4) 
                           => reg_a_out(4), output(3) => reg_a_out(3), 
                           output(2) => reg_a_out(2), output(1) => reg_a_out(1)
                           , output(0) => reg_a_out(0), match_dirty_f => 
                           sig_bal, match_dirty_ff => net1291);
   FWDMUX_2AJ : FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_4 port map( reg_c(31) => 
                           s2_a_31_port, reg_c(30) => s2_a_30_port, reg_c(29) 
                           => s2_a_29_port, reg_c(28) => s2_a_28_port, 
                           reg_c(27) => s2_a_27_port, reg_c(26) => s2_a_26_port
                           , reg_c(25) => s2_a_25_port, reg_c(24) => 
                           s2_a_24_port, reg_c(23) => s2_a_23_port, reg_c(22) 
                           => s2_a_22_port, reg_c(21) => s2_a_21_port, 
                           reg_c(20) => s2_a_20_port, reg_c(19) => s2_a_19_port
                           , reg_c(18) => s2_a_18_port, reg_c(17) => 
                           s2_a_17_port, reg_c(16) => s2_a_16_port, reg_c(15) 
                           => s2_a_15_port, reg_c(14) => s2_a_14_port, 
                           reg_c(13) => s2_a_13_port, reg_c(12) => s2_a_12_port
                           , reg_c(11) => s2_a_11_port, reg_c(10) => 
                           s2_a_10_port, reg_c(9) => s2_a_9_port, reg_c(8) => 
                           s2_a_8_port, reg_c(7) => s2_a_7_port, reg_c(6) => 
                           s2_a_6_port, reg_c(5) => s2_a_5_port, reg_c(4) => 
                           s2_a_4_port, reg_c(3) => s2_a_3_port, reg_c(2) => 
                           s2_a_2_port, reg_c(1) => s2_a_1_port, reg_c(0) => 
                           s2_a_0_port, reg_f(31) => n83, reg_f(30) => n80, 
                           reg_f(29) => n81, reg_f(28) => n82, reg_f(27) => 
                           s3_exe_out_27_port, reg_f(26) => s3_exe_out_26_port,
                           reg_f(25) => s3_exe_out_25_port, reg_f(24) => 
                           s3_exe_out_24_port, reg_f(23) => s3_exe_out_23_port,
                           reg_f(22) => s3_exe_out_22_port, reg_f(21) => 
                           s3_exe_out_21_port, reg_f(20) => s3_exe_out_20_port,
                           reg_f(19) => s3_exe_out_19_port, reg_f(18) => 
                           s3_exe_out_18_port, reg_f(17) => s3_exe_out_17_port,
                           reg_f(16) => s3_exe_out_16_port, reg_f(15) => 
                           s3_exe_out_15_port, reg_f(14) => s3_exe_out_14_port,
                           reg_f(13) => s3_exe_out_13_port, reg_f(12) => 
                           s3_exe_out_12_port, reg_f(11) => s3_exe_out_11_port,
                           reg_f(10) => s3_exe_out_10_port, reg_f(9) => 
                           s3_exe_out_9_port, reg_f(8) => s3_exe_out_8_port, 
                           reg_f(7) => s3_exe_out_7_port, reg_f(6) => 
                           s3_exe_out_6_port, reg_f(5) => s3_exe_out_5_port, 
                           reg_f(4) => s3_exe_out_4_port, reg_f(3) => 
                           s3_exe_out_3_port, reg_f(2) => s3_exe_out_2_port, 
                           reg_f(1) => s3_exe_out_1_port, reg_f(0) => n105, 
                           reg_ff(31) => s4_result_31_port, reg_ff(30) => 
                           s4_result_30_port, reg_ff(29) => s4_result_29_port, 
                           reg_ff(28) => s4_result_28_port, reg_ff(27) => 
                           s4_result_27_port, reg_ff(26) => s4_result_26_port, 
                           reg_ff(25) => s4_result_25_port, reg_ff(24) => 
                           s4_result_24_port, reg_ff(23) => s4_result_23_port, 
                           reg_ff(22) => s4_result_22_port, reg_ff(21) => 
                           s4_result_21_port, reg_ff(20) => s4_result_20_port, 
                           reg_ff(19) => s4_result_19_port, reg_ff(18) => 
                           s4_result_18_port, reg_ff(17) => s4_result_17_port, 
                           reg_ff(16) => s4_result_16_port, reg_ff(15) => 
                           s4_result_15_port, reg_ff(14) => s4_result_14_port, 
                           reg_ff(13) => s4_result_13_port, reg_ff(12) => 
                           s4_result_12_port, reg_ff(11) => s4_result_11_port, 
                           reg_ff(10) => s4_result_10_port, reg_ff(9) => 
                           s4_result_9_port, reg_ff(8) => s4_result_8_port, 
                           reg_ff(7) => s4_result_7_port, reg_ff(6) => 
                           s4_result_6_port, reg_ff(5) => s4_result_5_port, 
                           reg_ff(4) => s4_result_4_port, reg_ff(3) => 
                           s4_result_3_port, reg_ff(2) => s4_result_2_port, 
                           reg_ff(1) => s4_result_1_port, reg_ff(0) => 
                           s4_result_0_port, addr_c(4) => istr_val(25), 
                           addr_c(3) => istr_val(24), addr_c(2) => istr_val(23)
                           , addr_c(1) => istr_val(22), addr_c(0) => 
                           istr_val(21), addr_f(4) => s3_wr_addr_4_port, 
                           addr_f(3) => s3_wr_addr_3_port, addr_f(2) => 
                           s3_wr_addr_2_port, addr_f(1) => s3_wr_addr_1_port, 
                           addr_f(0) => s3_wr_addr_0_port, addr_ff(4) => 
                           s4_wr_addr_4_port, addr_ff(3) => s4_wr_addr_3_port, 
                           addr_ff(2) => s4_wr_addr_2_port, addr_ff(1) => 
                           s4_wr_addr_1_port, addr_ff(0) => s4_wr_addr_0_port, 
                           valid_f => s2_a_f_j_en, valid_ff => s2_a_ff_j_en, 
                           dirty_f => cw(8), dirty_ff => X_Logic0_port, en => 
                           X_Logic1_port, output(31) => 
                           s2_jump_addr_reg_31_port, output(30) => 
                           s2_jump_addr_reg_30_port, output(29) => 
                           s2_jump_addr_reg_29_port, output(28) => 
                           s2_jump_addr_reg_28_port, output(27) => 
                           s2_jump_addr_reg_27_port, output(26) => 
                           s2_jump_addr_reg_26_port, output(25) => 
                           s2_jump_addr_reg_25_port, output(24) => 
                           s2_jump_addr_reg_24_port, output(23) => 
                           s2_jump_addr_reg_23_port, output(22) => 
                           s2_jump_addr_reg_22_port, output(21) => 
                           s2_jump_addr_reg_21_port, output(20) => 
                           s2_jump_addr_reg_20_port, output(19) => 
                           s2_jump_addr_reg_19_port, output(18) => 
                           s2_jump_addr_reg_18_port, output(17) => 
                           s2_jump_addr_reg_17_port, output(16) => 
                           s2_jump_addr_reg_16_port, output(15) => 
                           s2_jump_addr_reg_15_port, output(14) => 
                           s2_jump_addr_reg_14_port, output(13) => 
                           s2_jump_addr_reg_13_port, output(12) => 
                           s2_jump_addr_reg_12_port, output(11) => 
                           s2_jump_addr_reg_11_port, output(10) => 
                           s2_jump_addr_reg_10_port, output(9) => 
                           s2_jump_addr_reg_9_port, output(8) => 
                           s2_jump_addr_reg_8_port, output(7) => 
                           s2_jump_addr_reg_7_port, output(6) => 
                           s2_jump_addr_reg_6_port, output(5) => 
                           s2_jump_addr_reg_5_port, output(4) => 
                           s2_jump_addr_reg_4_port, output(3) => 
                           s2_jump_addr_reg_3_port, output(2) => 
                           s2_jump_addr_reg_2_port, output(1) => 
                           s2_jump_addr_reg_1_port, output(0) => 
                           s2_jump_addr_reg_0_port, match_dirty_f => sig_jral, 
                           match_dirty_ff => net1290);
   REG_A : Reg_DATA_SIZE32_11 port map( rst => n110, en => cw(6), clk => clk, 
                           din(31) => s2_a_31_port, din(30) => s2_a_30_port, 
                           din(29) => s2_a_29_port, din(28) => s2_a_28_port, 
                           din(27) => s2_a_27_port, din(26) => s2_a_26_port, 
                           din(25) => s2_a_25_port, din(24) => s2_a_24_port, 
                           din(23) => s2_a_23_port, din(22) => s2_a_22_port, 
                           din(21) => s2_a_21_port, din(20) => s2_a_20_port, 
                           din(19) => s2_a_19_port, din(18) => s2_a_18_port, 
                           din(17) => s2_a_17_port, din(16) => s2_a_16_port, 
                           din(15) => s2_a_15_port, din(14) => s2_a_14_port, 
                           din(13) => s2_a_13_port, din(12) => s2_a_12_port, 
                           din(11) => s2_a_11_port, din(10) => s2_a_10_port, 
                           din(9) => s2_a_9_port, din(8) => s2_a_8_port, din(7)
                           => s2_a_7_port, din(6) => s2_a_6_port, din(5) => 
                           s2_a_5_port, din(4) => s2_a_4_port, din(3) => 
                           s2_a_3_port, din(2) => s2_a_2_port, din(1) => 
                           s2_a_1_port, din(0) => s2_a_0_port, dout(31) => 
                           s3_a_31_port, dout(30) => s3_a_30_port, dout(29) => 
                           s3_a_29_port, dout(28) => s3_a_28_port, dout(27) => 
                           s3_a_27_port, dout(26) => s3_a_26_port, dout(25) => 
                           s3_a_25_port, dout(24) => s3_a_24_port, dout(23) => 
                           s3_a_23_port, dout(22) => s3_a_22_port, dout(21) => 
                           s3_a_21_port, dout(20) => s3_a_20_port, dout(19) => 
                           s3_a_19_port, dout(18) => s3_a_18_port, dout(17) => 
                           s3_a_17_port, dout(16) => s3_a_16_port, dout(15) => 
                           s3_a_15_port, dout(14) => s3_a_14_port, dout(13) => 
                           s3_a_13_port, dout(12) => s3_a_12_port, dout(11) => 
                           s3_a_11_port, dout(10) => s3_a_10_port, dout(9) => 
                           s3_a_9_port, dout(8) => s3_a_8_port, dout(7) => 
                           s3_a_7_port, dout(6) => s3_a_6_port, dout(5) => 
                           s3_a_5_port, dout(4) => s3_a_4_port, dout(3) => 
                           s3_a_3_port, dout(2) => s3_a_2_port, dout(1) => 
                           s3_a_1_port, dout(0) => s3_a_0_port);
   REG_B : Reg_DATA_SIZE32_10 port map( rst => n111, en => cw(6), clk => clk, 
                           din(31) => s2_b_31_port, din(30) => s2_b_30_port, 
                           din(29) => s2_b_29_port, din(28) => s2_b_28_port, 
                           din(27) => s2_b_27_port, din(26) => s2_b_26_port, 
                           din(25) => s2_b_25_port, din(24) => s2_b_24_port, 
                           din(23) => s2_b_23_port, din(22) => s2_b_22_port, 
                           din(21) => s2_b_21_port, din(20) => s2_b_20_port, 
                           din(19) => s2_b_19_port, din(18) => s2_b_18_port, 
                           din(17) => s2_b_17_port, din(16) => s2_b_16_port, 
                           din(15) => s2_b_15_port, din(14) => s2_b_14_port, 
                           din(13) => s2_b_13_port, din(12) => s2_b_12_port, 
                           din(11) => s2_b_11_port, din(10) => s2_b_10_port, 
                           din(9) => s2_b_9_port, din(8) => s2_b_8_port, din(7)
                           => s2_b_7_port, din(6) => s2_b_6_port, din(5) => 
                           s2_b_5_port, din(4) => s2_b_4_port, din(3) => 
                           s2_b_3_port, din(2) => s2_b_2_port, din(1) => 
                           s2_b_1_port, din(0) => s2_b_0_port, dout(31) => 
                           s3_b_31_port, dout(30) => s3_b_30_port, dout(29) => 
                           s3_b_29_port, dout(28) => s3_b_28_port, dout(27) => 
                           s3_b_27_port, dout(26) => s3_b_26_port, dout(25) => 
                           s3_b_25_port, dout(24) => s3_b_24_port, dout(23) => 
                           s3_b_23_port, dout(22) => s3_b_22_port, dout(21) => 
                           s3_b_21_port, dout(20) => s3_b_20_port, dout(19) => 
                           s3_b_19_port, dout(18) => s3_b_18_port, dout(17) => 
                           s3_b_17_port, dout(16) => s3_b_16_port, dout(15) => 
                           s3_b_15_port, dout(14) => s3_b_14_port, dout(13) => 
                           s3_b_13_port, dout(12) => s3_b_12_port, dout(11) => 
                           s3_b_11_port, dout(10) => s3_b_10_port, dout(9) => 
                           s3_b_9_port, dout(8) => s3_b_8_port, dout(7) => 
                           s3_b_7_port, dout(6) => s3_b_6_port, dout(5) => 
                           s3_b_5_port, dout(4) => s3_b_4_port, dout(3) => 
                           s3_b_3_port, dout(2) => s3_b_2_port, dout(1) => 
                           s3_b_1_port, dout(0) => s3_b_0_port);
   REG_I : Reg_DATA_SIZE32_9 port map( rst => n111, en => cw(6), clk => clk, 
                           din(31) => s2_imm_i_ext_31_port, din(30) => 
                           s2_imm_i_ext_30_port, din(29) => 
                           s2_imm_i_ext_29_port, din(28) => 
                           s2_imm_i_ext_28_port, din(27) => 
                           s2_imm_i_ext_27_port, din(26) => 
                           s2_imm_i_ext_26_port, din(25) => 
                           s2_imm_i_ext_25_port, din(24) => 
                           s2_imm_i_ext_24_port, din(23) => 
                           s2_imm_i_ext_23_port, din(22) => 
                           s2_imm_i_ext_22_port, din(21) => 
                           s2_imm_i_ext_21_port, din(20) => 
                           s2_imm_i_ext_20_port, din(19) => 
                           s2_imm_i_ext_19_port, din(18) => 
                           s2_imm_i_ext_18_port, din(17) => 
                           s2_imm_i_ext_17_port, din(16) => 
                           s2_imm_i_ext_16_port, din(15) => 
                           s2_imm_i_ext_15_port, din(14) => 
                           s2_imm_i_ext_14_port, din(13) => 
                           s2_imm_i_ext_13_port, din(12) => 
                           s2_imm_i_ext_12_port, din(11) => 
                           s2_imm_i_ext_11_port, din(10) => 
                           s2_imm_i_ext_10_port, din(9) => s2_imm_i_ext_9_port,
                           din(8) => s2_imm_i_ext_8_port, din(7) => 
                           s2_imm_i_ext_7_port, din(6) => s2_imm_i_ext_6_port, 
                           din(5) => s2_imm_i_ext_5_port, din(4) => 
                           s2_imm_i_ext_4_port, din(3) => s2_imm_i_ext_3_port, 
                           din(2) => s2_imm_i_ext_2_port, din(1) => 
                           s2_imm_i_ext_1_port, din(0) => s2_imm_i_ext_0_port, 
                           dout(31) => s3_imm_i_ext_31_port, dout(30) => 
                           s3_imm_i_ext_30_port, dout(29) => 
                           s3_imm_i_ext_29_port, dout(28) => 
                           s3_imm_i_ext_28_port, dout(27) => 
                           s3_imm_i_ext_27_port, dout(26) => 
                           s3_imm_i_ext_26_port, dout(25) => 
                           s3_imm_i_ext_25_port, dout(24) => 
                           s3_imm_i_ext_24_port, dout(23) => 
                           s3_imm_i_ext_23_port, dout(22) => 
                           s3_imm_i_ext_22_port, dout(21) => 
                           s3_imm_i_ext_21_port, dout(20) => 
                           s3_imm_i_ext_20_port, dout(19) => 
                           s3_imm_i_ext_19_port, dout(18) => 
                           s3_imm_i_ext_18_port, dout(17) => 
                           s3_imm_i_ext_17_port, dout(16) => 
                           s3_imm_i_ext_16_port, dout(15) => 
                           s3_imm_i_ext_15_port, dout(14) => 
                           s3_imm_i_ext_14_port, dout(13) => 
                           s3_imm_i_ext_13_port, dout(12) => 
                           s3_imm_i_ext_12_port, dout(11) => 
                           s3_imm_i_ext_11_port, dout(10) => 
                           s3_imm_i_ext_10_port, dout(9) => s3_imm_i_ext_9_port
                           , dout(8) => s3_imm_i_ext_8_port, dout(7) => 
                           s3_imm_i_ext_7_port, dout(6) => s3_imm_i_ext_6_port,
                           dout(5) => s3_imm_i_ext_5_port, dout(4) => 
                           s3_imm_i_ext_4_port, dout(3) => s3_imm_i_ext_3_port,
                           dout(2) => s3_imm_i_ext_2_port, dout(1) => 
                           s3_imm_i_ext_1_port, dout(0) => s3_imm_i_ext_0_port)
                           ;
   REG_WR2 : Reg_DATA_SIZE5_0 port map( rst => n110, en => cw(6), clk => clk, 
                           din(4) => s2_wr_addr_4_port, din(3) => 
                           s2_wr_addr_3_port, din(2) => s2_wr_addr_2_port, 
                           din(1) => s2_wr_addr_1_port, din(0) => 
                           s2_wr_addr_0_port, dout(4) => s3_wr_addr_4_port, 
                           dout(3) => s3_wr_addr_3_port, dout(2) => 
                           s3_wr_addr_2_port, dout(1) => s3_wr_addr_1_port, 
                           dout(0) => s3_wr_addr_0_port);
   REG_A_ADDR_2 : Reg_DATA_SIZE5_6 port map( rst => n110, en => cw(6), clk => 
                           clk, din(4) => istr_val(25), din(3) => istr_val(24),
                           din(2) => istr_val(23), din(1) => istr_val(22), 
                           din(0) => istr_val(21), dout(4) => 
                           s3_rd1_addr_4_port, dout(3) => s3_rd1_addr_3_port, 
                           dout(2) => s3_rd1_addr_2_port, dout(1) => 
                           s3_rd1_addr_1_port, dout(0) => s3_rd1_addr_0_port);
   REG_B_ADDR_2 : Reg_DATA_SIZE5_5 port map( rst => n110, en => cw(6), clk => 
                           clk, din(4) => istr_val(20), din(3) => istr_val(19),
                           din(2) => istr_val(18), din(1) => istr_val(17), 
                           din(0) => istr_val(16), dout(4) => 
                           s3_rd2_addr_4_port, dout(3) => s3_rd2_addr_3_port, 
                           dout(2) => s3_rd2_addr_2_port, dout(1) => 
                           s3_rd2_addr_1_port, dout(0) => s3_rd2_addr_0_port);
   REG_PC_NOT_SEL : Reg_DATA_SIZE32_8 port map( rst => n111, en => cw(6), clk 
                           => clk, din(31) => s2_pc_notsel_31_port, din(30) => 
                           s2_pc_notsel_30_port, din(29) => 
                           s2_pc_notsel_29_port, din(28) => 
                           s2_pc_notsel_28_port, din(27) => 
                           s2_pc_notsel_27_port, din(26) => 
                           s2_pc_notsel_26_port, din(25) => 
                           s2_pc_notsel_25_port, din(24) => 
                           s2_pc_notsel_24_port, din(23) => 
                           s2_pc_notsel_23_port, din(22) => 
                           s2_pc_notsel_22_port, din(21) => 
                           s2_pc_notsel_21_port, din(20) => 
                           s2_pc_notsel_20_port, din(19) => 
                           s2_pc_notsel_19_port, din(18) => 
                           s2_pc_notsel_18_port, din(17) => 
                           s2_pc_notsel_17_port, din(16) => 
                           s2_pc_notsel_16_port, din(15) => 
                           s2_pc_notsel_15_port, din(14) => 
                           s2_pc_notsel_14_port, din(13) => 
                           s2_pc_notsel_13_port, din(12) => 
                           s2_pc_notsel_12_port, din(11) => 
                           s2_pc_notsel_11_port, din(10) => 
                           s2_pc_notsel_10_port, din(9) => s2_pc_notsel_9_port,
                           din(8) => s2_pc_notsel_8_port, din(7) => 
                           s2_pc_notsel_7_port, din(6) => s2_pc_notsel_6_port, 
                           din(5) => s2_pc_notsel_5_port, din(4) => 
                           s2_pc_notsel_4_port, din(3) => s2_pc_notsel_3_port, 
                           din(2) => s2_pc_notsel_2_port, din(1) => 
                           s2_pc_notsel_1_port, din(0) => s2_pc_notsel_0_port, 
                           dout(31) => s3_pc_notsel_31_port, dout(30) => 
                           s3_pc_notsel_30_port, dout(29) => 
                           s3_pc_notsel_29_port, dout(28) => 
                           s3_pc_notsel_28_port, dout(27) => 
                           s3_pc_notsel_27_port, dout(26) => 
                           s3_pc_notsel_26_port, dout(25) => 
                           s3_pc_notsel_25_port, dout(24) => 
                           s3_pc_notsel_24_port, dout(23) => 
                           s3_pc_notsel_23_port, dout(22) => 
                           s3_pc_notsel_22_port, dout(21) => 
                           s3_pc_notsel_21_port, dout(20) => 
                           s3_pc_notsel_20_port, dout(19) => 
                           s3_pc_notsel_19_port, dout(18) => 
                           s3_pc_notsel_18_port, dout(17) => 
                           s3_pc_notsel_17_port, dout(16) => 
                           s3_pc_notsel_16_port, dout(15) => 
                           s3_pc_notsel_15_port, dout(14) => 
                           s3_pc_notsel_14_port, dout(13) => 
                           s3_pc_notsel_13_port, dout(12) => 
                           s3_pc_notsel_12_port, dout(11) => 
                           s3_pc_notsel_11_port, dout(10) => 
                           s3_pc_notsel_10_port, dout(9) => s3_pc_notsel_9_port
                           , dout(8) => s3_pc_notsel_8_port, dout(7) => 
                           s3_pc_notsel_7_port, dout(6) => s3_pc_notsel_6_port,
                           dout(5) => s3_pc_notsel_5_port, dout(4) => 
                           s3_pc_notsel_4_port, dout(3) => s3_pc_notsel_3_port,
                           dout(2) => s3_pc_notsel_2_port, dout(1) => 
                           s3_pc_notsel_1_port, dout(0) => s3_pc_notsel_0_port)
                           ;
   MUX_KEEP_A : Mux_DATA_SIZE32_5 port map( sel => s4_reg_b_wait, din0(31) => 
                           s3_a_31_port, din0(30) => s3_a_30_port, din0(29) => 
                           s3_a_29_port, din0(28) => s3_a_28_port, din0(27) => 
                           s3_a_27_port, din0(26) => s3_a_26_port, din0(25) => 
                           s3_a_25_port, din0(24) => s3_a_24_port, din0(23) => 
                           s3_a_23_port, din0(22) => s3_a_22_port, din0(21) => 
                           s3_a_21_port, din0(20) => s3_a_20_port, din0(19) => 
                           s3_a_19_port, din0(18) => s3_a_18_port, din0(17) => 
                           s3_a_17_port, din0(16) => s3_a_16_port, din0(15) => 
                           s3_a_15_port, din0(14) => s3_a_14_port, din0(13) => 
                           s3_a_13_port, din0(12) => s3_a_12_port, din0(11) => 
                           s3_a_11_port, din0(10) => s3_a_10_port, din0(9) => 
                           s3_a_9_port, din0(8) => s3_a_8_port, din0(7) => 
                           s3_a_7_port, din0(6) => s3_a_6_port, din0(5) => 
                           s3_a_5_port, din0(4) => s3_a_4_port, din0(3) => 
                           s3_a_3_port, din0(2) => s3_a_2_port, din0(1) => 
                           s3_a_1_port, din0(0) => s3_a_0_port, din1(31) => 
                           s4_a_31_port, din1(30) => s4_a_30_port, din1(29) => 
                           s4_a_29_port, din1(28) => s4_a_28_port, din1(27) => 
                           s4_a_27_port, din1(26) => s4_a_26_port, din1(25) => 
                           s4_a_25_port, din1(24) => s4_a_24_port, din1(23) => 
                           s4_a_23_port, din1(22) => s4_a_22_port, din1(21) => 
                           s4_a_21_port, din1(20) => s4_a_20_port, din1(19) => 
                           s4_a_19_port, din1(18) => s4_a_18_port, din1(17) => 
                           s4_a_17_port, din1(16) => s4_a_16_port, din1(15) => 
                           s4_a_15_port, din1(14) => s4_a_14_port, din1(13) => 
                           s4_a_13_port, din1(12) => s4_a_12_port, din1(11) => 
                           s4_a_11_port, din1(10) => s4_a_10_port, din1(9) => 
                           s4_a_9_port, din1(8) => s4_a_8_port, din1(7) => 
                           s4_a_7_port, din1(6) => s4_a_6_port, din1(5) => 
                           s4_a_5_port, din1(4) => s4_a_4_port, din1(3) => 
                           s4_a_3_port, din1(2) => s4_a_2_port, din1(1) => 
                           s4_a_1_port, din1(0) => s4_a_0_port, dout(31) => 
                           s3_a_keep_31_port, dout(30) => s3_a_keep_30_port, 
                           dout(29) => s3_a_keep_29_port, dout(28) => 
                           s3_a_keep_28_port, dout(27) => s3_a_keep_27_port, 
                           dout(26) => s3_a_keep_26_port, dout(25) => 
                           s3_a_keep_25_port, dout(24) => s3_a_keep_24_port, 
                           dout(23) => s3_a_keep_23_port, dout(22) => 
                           s3_a_keep_22_port, dout(21) => s3_a_keep_21_port, 
                           dout(20) => s3_a_keep_20_port, dout(19) => 
                           s3_a_keep_19_port, dout(18) => s3_a_keep_18_port, 
                           dout(17) => s3_a_keep_17_port, dout(16) => 
                           s3_a_keep_16_port, dout(15) => s3_a_keep_15_port, 
                           dout(14) => s3_a_keep_14_port, dout(13) => 
                           s3_a_keep_13_port, dout(12) => s3_a_keep_12_port, 
                           dout(11) => s3_a_keep_11_port, dout(10) => 
                           s3_a_keep_10_port, dout(9) => s3_a_keep_9_port, 
                           dout(8) => s3_a_keep_8_port, dout(7) => 
                           s3_a_keep_7_port, dout(6) => s3_a_keep_6_port, 
                           dout(5) => s3_a_keep_5_port, dout(4) => 
                           s3_a_keep_4_port, dout(3) => s3_a_keep_3_port, 
                           dout(2) => s3_a_keep_2_port, dout(1) => 
                           s3_a_keep_1_port, dout(0) => s3_a_keep_0_port);
   MUX_KEEP_B : Mux_DATA_SIZE32_4 port map( sel => s4_reg_a_wait, din0(31) => 
                           s3_b_31_port, din0(30) => s3_b_30_port, din0(29) => 
                           s3_b_29_port, din0(28) => s3_b_28_port, din0(27) => 
                           s3_b_27_port, din0(26) => s3_b_26_port, din0(25) => 
                           s3_b_25_port, din0(24) => s3_b_24_port, din0(23) => 
                           s3_b_23_port, din0(22) => s3_b_22_port, din0(21) => 
                           s3_b_21_port, din0(20) => s3_b_20_port, din0(19) => 
                           s3_b_19_port, din0(18) => s3_b_18_port, din0(17) => 
                           s3_b_17_port, din0(16) => s3_b_16_port, din0(15) => 
                           s3_b_15_port, din0(14) => s3_b_14_port, din0(13) => 
                           s3_b_13_port, din0(12) => s3_b_12_port, din0(11) => 
                           s3_b_11_port, din0(10) => s3_b_10_port, din0(9) => 
                           s3_b_9_port, din0(8) => s3_b_8_port, din0(7) => 
                           s3_b_7_port, din0(6) => s3_b_6_port, din0(5) => 
                           s3_b_5_port, din0(4) => s3_b_4_port, din0(3) => 
                           s3_b_3_port, din0(2) => s3_b_2_port, din0(1) => 
                           s3_b_1_port, din0(0) => s3_b_0_port, din1(31) => 
                           s4_b_31_port, din1(30) => s4_b_30_port, din1(29) => 
                           s4_b_29_port, din1(28) => s4_b_28_port, din1(27) => 
                           s4_b_27_port, din1(26) => s4_b_26_port, din1(25) => 
                           s4_b_25_port, din1(24) => s4_b_24_port, din1(23) => 
                           s4_b_23_port, din1(22) => s4_b_22_port, din1(21) => 
                           s4_b_21_port, din1(20) => s4_b_20_port, din1(19) => 
                           s4_b_19_port, din1(18) => s4_b_18_port, din1(17) => 
                           s4_b_17_port, din1(16) => s4_b_16_port, din1(15) => 
                           s4_b_15_port, din1(14) => s4_b_14_port, din1(13) => 
                           s4_b_13_port, din1(12) => s4_b_12_port, din1(11) => 
                           s4_b_11_port, din1(10) => s4_b_10_port, din1(9) => 
                           s4_b_9_port, din1(8) => s4_b_8_port, din1(7) => 
                           s4_b_7_port, din1(6) => s4_b_6_port, din1(5) => 
                           s4_b_5_port, din1(4) => s4_b_4_port, din1(3) => 
                           s4_b_3_port, din1(2) => s4_b_2_port, din1(1) => 
                           s4_b_1_port, din1(0) => s4_b_0_port, dout(31) => 
                           s3_b_keep_31_port, dout(30) => s3_b_keep_30_port, 
                           dout(29) => s3_b_keep_29_port, dout(28) => 
                           s3_b_keep_28_port, dout(27) => s3_b_keep_27_port, 
                           dout(26) => s3_b_keep_26_port, dout(25) => 
                           s3_b_keep_25_port, dout(24) => s3_b_keep_24_port, 
                           dout(23) => s3_b_keep_23_port, dout(22) => 
                           s3_b_keep_22_port, dout(21) => s3_b_keep_21_port, 
                           dout(20) => s3_b_keep_20_port, dout(19) => 
                           s3_b_keep_19_port, dout(18) => s3_b_keep_18_port, 
                           dout(17) => s3_b_keep_17_port, dout(16) => 
                           s3_b_keep_16_port, dout(15) => s3_b_keep_15_port, 
                           dout(14) => s3_b_keep_14_port, dout(13) => 
                           s3_b_keep_13_port, dout(12) => s3_b_keep_12_port, 
                           dout(11) => s3_b_keep_11_port, dout(10) => 
                           s3_b_keep_10_port, dout(9) => s3_b_keep_9_port, 
                           dout(8) => s3_b_keep_8_port, dout(7) => 
                           s3_b_keep_7_port, dout(6) => s3_b_keep_6_port, 
                           dout(5) => s3_b_keep_5_port, dout(4) => 
                           s3_b_keep_4_port, dout(3) => s3_b_keep_3_port, 
                           dout(2) => s3_b_keep_2_port, dout(1) => 
                           s3_b_keep_1_port, dout(0) => s3_b_keep_0_port);
   FWDMUX_A : FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_3 port map( reg_c(31) => 
                           s3_a_keep_31_port, reg_c(30) => s3_a_keep_30_port, 
                           reg_c(29) => s3_a_keep_29_port, reg_c(28) => 
                           s3_a_keep_28_port, reg_c(27) => s3_a_keep_27_port, 
                           reg_c(26) => s3_a_keep_26_port, reg_c(25) => 
                           s3_a_keep_25_port, reg_c(24) => s3_a_keep_24_port, 
                           reg_c(23) => s3_a_keep_23_port, reg_c(22) => 
                           s3_a_keep_22_port, reg_c(21) => s3_a_keep_21_port, 
                           reg_c(20) => s3_a_keep_20_port, reg_c(19) => 
                           s3_a_keep_19_port, reg_c(18) => s3_a_keep_18_port, 
                           reg_c(17) => s3_a_keep_17_port, reg_c(16) => 
                           s3_a_keep_16_port, reg_c(15) => s3_a_keep_15_port, 
                           reg_c(14) => s3_a_keep_14_port, reg_c(13) => 
                           s3_a_keep_13_port, reg_c(12) => s3_a_keep_12_port, 
                           reg_c(11) => s3_a_keep_11_port, reg_c(10) => 
                           s3_a_keep_10_port, reg_c(9) => s3_a_keep_9_port, 
                           reg_c(8) => s3_a_keep_8_port, reg_c(7) => 
                           s3_a_keep_7_port, reg_c(6) => s3_a_keep_6_port, 
                           reg_c(5) => s3_a_keep_5_port, reg_c(4) => 
                           s3_a_keep_4_port, reg_c(3) => s3_a_keep_3_port, 
                           reg_c(2) => s3_a_keep_2_port, reg_c(1) => 
                           s3_a_keep_1_port, reg_c(0) => s3_a_keep_0_port, 
                           reg_f(31) => data_addr_31_port, reg_f(30) => 
                           data_addr_30_port, reg_f(29) => data_addr_29_port, 
                           reg_f(28) => data_addr_28_port, reg_f(27) => 
                           data_addr_27_port, reg_f(26) => data_addr_26_port, 
                           reg_f(25) => data_addr_25_port, reg_f(24) => 
                           data_addr_24_port, reg_f(23) => data_addr_23_port, 
                           reg_f(22) => data_addr_22_port, reg_f(21) => 
                           data_addr_21_port, reg_f(20) => data_addr_20_port, 
                           reg_f(19) => data_addr_19_port, reg_f(18) => 
                           data_addr_18_port, reg_f(17) => data_addr_17_port, 
                           reg_f(16) => data_addr_16_port, reg_f(15) => 
                           data_addr_15_port, reg_f(14) => data_addr_14_port, 
                           reg_f(13) => data_addr_13_port, reg_f(12) => 
                           data_addr_12_port, reg_f(11) => data_addr_11_port, 
                           reg_f(10) => data_addr_10_port, reg_f(9) => 
                           data_addr_9_port, reg_f(8) => data_addr_8_port, 
                           reg_f(7) => data_addr_7_port, reg_f(6) => 
                           data_addr_6_port, reg_f(5) => data_addr_5_port, 
                           reg_f(4) => data_addr_4_port, reg_f(3) => 
                           data_addr_3_port, reg_f(2) => data_addr_2_port, 
                           reg_f(1) => data_addr_1_port, reg_f(0) => 
                           data_addr_0_port, reg_ff(31) => s5_result_31_port, 
                           reg_ff(30) => s5_result_30_port, reg_ff(29) => 
                           s5_result_29_port, reg_ff(28) => s5_result_28_port, 
                           reg_ff(27) => s5_result_27_port, reg_ff(26) => 
                           s5_result_26_port, reg_ff(25) => s5_result_25_port, 
                           reg_ff(24) => s5_result_24_port, reg_ff(23) => 
                           s5_result_23_port, reg_ff(22) => s5_result_22_port, 
                           reg_ff(21) => s5_result_21_port, reg_ff(20) => 
                           s5_result_20_port, reg_ff(19) => s5_result_19_port, 
                           reg_ff(18) => s5_result_18_port, reg_ff(17) => 
                           s5_result_17_port, reg_ff(16) => s5_result_16_port, 
                           reg_ff(15) => s5_result_15_port, reg_ff(14) => 
                           s5_result_14_port, reg_ff(13) => s5_result_13_port, 
                           reg_ff(12) => s5_result_12_port, reg_ff(11) => 
                           s5_result_11_port, reg_ff(10) => s5_result_10_port, 
                           reg_ff(9) => s5_result_9_port, reg_ff(8) => 
                           s5_result_8_port, reg_ff(7) => s5_result_7_port, 
                           reg_ff(6) => s5_result_6_port, reg_ff(5) => 
                           s5_result_5_port, reg_ff(4) => s5_result_4_port, 
                           reg_ff(3) => s5_result_3_port, reg_ff(2) => 
                           s5_result_2_port, reg_ff(1) => s5_result_1_port, 
                           reg_ff(0) => s5_result_0_port, addr_c(4) => 
                           s3_rd1_addr_4_port, addr_c(3) => s3_rd1_addr_3_port,
                           addr_c(2) => s3_rd1_addr_2_port, addr_c(1) => 
                           s3_rd1_addr_1_port, addr_c(0) => s3_rd1_addr_0_port,
                           addr_f(4) => s4_wr_addr_4_port, addr_f(3) => 
                           s4_wr_addr_3_port, addr_f(2) => s4_wr_addr_2_port, 
                           addr_f(1) => s4_wr_addr_1_port, addr_f(0) => 
                           s4_wr_addr_0_port, addr_ff(4) => s5_wr_addr_4_port, 
                           addr_ff(3) => s5_wr_addr_3_port, addr_ff(2) => 
                           s5_wr_addr_2_port, addr_ff(1) => s5_wr_addr_1_port, 
                           addr_ff(0) => s5_wr_addr_0_port, valid_f => 
                           s3_a_sel_f_en, valid_ff => s3_a_sel_ff_en, dirty_f 
                           => cw(16), dirty_ff => X_Logic0_port, en => 
                           X_Logic1_port, output(31) => s3_a_sel_31_port, 
                           output(30) => s3_a_sel_30_port, output(29) => 
                           s3_a_sel_29_port, output(28) => s3_a_sel_28_port, 
                           output(27) => s3_a_sel_27_port, output(26) => 
                           s3_a_sel_26_port, output(25) => s3_a_sel_25_port, 
                           output(24) => s3_a_sel_24_port, output(23) => 
                           s3_a_sel_23_port, output(22) => s3_a_sel_22_port, 
                           output(21) => s3_a_sel_21_port, output(20) => 
                           s3_a_sel_20_port, output(19) => s3_a_sel_19_port, 
                           output(18) => s3_a_sel_18_port, output(17) => 
                           s3_a_sel_17_port, output(16) => s3_a_sel_16_port, 
                           output(15) => s3_a_sel_15_port, output(14) => 
                           s3_a_sel_14_port, output(13) => s3_a_sel_13_port, 
                           output(12) => s3_a_sel_12_port, output(11) => 
                           s3_a_sel_11_port, output(10) => s3_a_sel_10_port, 
                           output(9) => s3_a_sel_9_port, output(8) => 
                           s3_a_sel_8_port, output(7) => s3_a_sel_7_port, 
                           output(6) => s3_a_sel_6_port, output(5) => 
                           s3_a_sel_5_port, output(4) => s3_a_sel_4_port, 
                           output(3) => s3_a_sel_3_port, output(2) => 
                           s3_a_sel_2_port, output(1) => s3_a_sel_1_port, 
                           output(0) => s3_a_sel_0_port, match_dirty_f => 
                           s3_reg_a_wait, match_dirty_ff => net1288);
   FWDMUX_B : FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_2 port map( reg_c(31) => 
                           s3_b_keep_31_port, reg_c(30) => s3_b_keep_30_port, 
                           reg_c(29) => s3_b_keep_29_port, reg_c(28) => 
                           s3_b_keep_28_port, reg_c(27) => s3_b_keep_27_port, 
                           reg_c(26) => s3_b_keep_26_port, reg_c(25) => 
                           s3_b_keep_25_port, reg_c(24) => s3_b_keep_24_port, 
                           reg_c(23) => s3_b_keep_23_port, reg_c(22) => 
                           s3_b_keep_22_port, reg_c(21) => s3_b_keep_21_port, 
                           reg_c(20) => s3_b_keep_20_port, reg_c(19) => 
                           s3_b_keep_19_port, reg_c(18) => s3_b_keep_18_port, 
                           reg_c(17) => s3_b_keep_17_port, reg_c(16) => 
                           s3_b_keep_16_port, reg_c(15) => s3_b_keep_15_port, 
                           reg_c(14) => s3_b_keep_14_port, reg_c(13) => 
                           s3_b_keep_13_port, reg_c(12) => s3_b_keep_12_port, 
                           reg_c(11) => s3_b_keep_11_port, reg_c(10) => 
                           s3_b_keep_10_port, reg_c(9) => s3_b_keep_9_port, 
                           reg_c(8) => s3_b_keep_8_port, reg_c(7) => 
                           s3_b_keep_7_port, reg_c(6) => s3_b_keep_6_port, 
                           reg_c(5) => s3_b_keep_5_port, reg_c(4) => 
                           s3_b_keep_4_port, reg_c(3) => s3_b_keep_3_port, 
                           reg_c(2) => s3_b_keep_2_port, reg_c(1) => 
                           s3_b_keep_1_port, reg_c(0) => s3_b_keep_0_port, 
                           reg_f(31) => data_addr_31_port, reg_f(30) => 
                           data_addr_30_port, reg_f(29) => data_addr_29_port, 
                           reg_f(28) => data_addr_28_port, reg_f(27) => 
                           data_addr_27_port, reg_f(26) => data_addr_26_port, 
                           reg_f(25) => data_addr_25_port, reg_f(24) => 
                           data_addr_24_port, reg_f(23) => data_addr_23_port, 
                           reg_f(22) => data_addr_22_port, reg_f(21) => 
                           data_addr_21_port, reg_f(20) => data_addr_20_port, 
                           reg_f(19) => data_addr_19_port, reg_f(18) => 
                           data_addr_18_port, reg_f(17) => data_addr_17_port, 
                           reg_f(16) => data_addr_16_port, reg_f(15) => 
                           data_addr_15_port, reg_f(14) => data_addr_14_port, 
                           reg_f(13) => data_addr_13_port, reg_f(12) => 
                           data_addr_12_port, reg_f(11) => data_addr_11_port, 
                           reg_f(10) => data_addr_10_port, reg_f(9) => 
                           data_addr_9_port, reg_f(8) => data_addr_8_port, 
                           reg_f(7) => data_addr_7_port, reg_f(6) => 
                           data_addr_6_port, reg_f(5) => data_addr_5_port, 
                           reg_f(4) => data_addr_4_port, reg_f(3) => 
                           data_addr_3_port, reg_f(2) => data_addr_2_port, 
                           reg_f(1) => data_addr_1_port, reg_f(0) => 
                           data_addr_0_port, reg_ff(31) => s5_result_31_port, 
                           reg_ff(30) => s5_result_30_port, reg_ff(29) => 
                           s5_result_29_port, reg_ff(28) => s5_result_28_port, 
                           reg_ff(27) => s5_result_27_port, reg_ff(26) => 
                           s5_result_26_port, reg_ff(25) => s5_result_25_port, 
                           reg_ff(24) => s5_result_24_port, reg_ff(23) => 
                           s5_result_23_port, reg_ff(22) => s5_result_22_port, 
                           reg_ff(21) => s5_result_21_port, reg_ff(20) => 
                           s5_result_20_port, reg_ff(19) => s5_result_19_port, 
                           reg_ff(18) => s5_result_18_port, reg_ff(17) => 
                           s5_result_17_port, reg_ff(16) => s5_result_16_port, 
                           reg_ff(15) => s5_result_15_port, reg_ff(14) => 
                           s5_result_14_port, reg_ff(13) => s5_result_13_port, 
                           reg_ff(12) => s5_result_12_port, reg_ff(11) => 
                           s5_result_11_port, reg_ff(10) => s5_result_10_port, 
                           reg_ff(9) => s5_result_9_port, reg_ff(8) => 
                           s5_result_8_port, reg_ff(7) => s5_result_7_port, 
                           reg_ff(6) => s5_result_6_port, reg_ff(5) => 
                           s5_result_5_port, reg_ff(4) => s5_result_4_port, 
                           reg_ff(3) => s5_result_3_port, reg_ff(2) => 
                           s5_result_2_port, reg_ff(1) => s5_result_1_port, 
                           reg_ff(0) => s5_result_0_port, addr_c(4) => 
                           s3_rd2_addr_4_port, addr_c(3) => s3_rd2_addr_3_port,
                           addr_c(2) => s3_rd2_addr_2_port, addr_c(1) => 
                           s3_rd2_addr_1_port, addr_c(0) => s3_rd2_addr_0_port,
                           addr_f(4) => s4_wr_addr_4_port, addr_f(3) => 
                           s4_wr_addr_3_port, addr_f(2) => s4_wr_addr_2_port, 
                           addr_f(1) => s4_wr_addr_1_port, addr_f(0) => 
                           s4_wr_addr_0_port, addr_ff(4) => s5_wr_addr_4_port, 
                           addr_ff(3) => s5_wr_addr_3_port, addr_ff(2) => 
                           s5_wr_addr_2_port, addr_ff(1) => s5_wr_addr_1_port, 
                           addr_ff(0) => s5_wr_addr_0_port, valid_f => 
                           s3_b_sel_f_en, valid_ff => s3_b_sel_ff_en, dirty_f 
                           => cw(16), dirty_ff => X_Logic0_port, en => 
                           X_Logic1_port, output(31) => s3_b_fwd_31_port, 
                           output(30) => s3_b_fwd_30_port, output(29) => 
                           s3_b_fwd_29_port, output(28) => s3_b_fwd_28_port, 
                           output(27) => s3_b_fwd_27_port, output(26) => 
                           s3_b_fwd_26_port, output(25) => s3_b_fwd_25_port, 
                           output(24) => s3_b_fwd_24_port, output(23) => 
                           s3_b_fwd_23_port, output(22) => s3_b_fwd_22_port, 
                           output(21) => s3_b_fwd_21_port, output(20) => 
                           s3_b_fwd_20_port, output(19) => s3_b_fwd_19_port, 
                           output(18) => s3_b_fwd_18_port, output(17) => 
                           s3_b_fwd_17_port, output(16) => s3_b_fwd_16_port, 
                           output(15) => s3_b_fwd_15_port, output(14) => 
                           s3_b_fwd_14_port, output(13) => s3_b_fwd_13_port, 
                           output(12) => s3_b_fwd_12_port, output(11) => 
                           s3_b_fwd_11_port, output(10) => s3_b_fwd_10_port, 
                           output(9) => s3_b_fwd_9_port, output(8) => 
                           s3_b_fwd_8_port, output(7) => s3_b_fwd_7_port, 
                           output(6) => s3_b_fwd_6_port, output(5) => 
                           s3_b_fwd_5_port, output(4) => s3_b_fwd_4_port, 
                           output(3) => s3_b_fwd_3_port, output(2) => 
                           s3_b_fwd_2_port, output(1) => s3_b_fwd_1_port, 
                           output(0) => s3_b_fwd_0_port, match_dirty_f => 
                           s3_reg_b_wait, match_dirty_ff => net1287);
   MUXB : Mux_DATA_SIZE32_3 port map( sel => cw(7), din0(31) => 
                           s3_b_fwd_31_port, din0(30) => s3_b_fwd_30_port, 
                           din0(29) => s3_b_fwd_29_port, din0(28) => 
                           s3_b_fwd_28_port, din0(27) => s3_b_fwd_27_port, 
                           din0(26) => s3_b_fwd_26_port, din0(25) => 
                           s3_b_fwd_25_port, din0(24) => s3_b_fwd_24_port, 
                           din0(23) => s3_b_fwd_23_port, din0(22) => 
                           s3_b_fwd_22_port, din0(21) => s3_b_fwd_21_port, 
                           din0(20) => s3_b_fwd_20_port, din0(19) => 
                           s3_b_fwd_19_port, din0(18) => s3_b_fwd_18_port, 
                           din0(17) => s3_b_fwd_17_port, din0(16) => 
                           s3_b_fwd_16_port, din0(15) => s3_b_fwd_15_port, 
                           din0(14) => s3_b_fwd_14_port, din0(13) => 
                           s3_b_fwd_13_port, din0(12) => s3_b_fwd_12_port, 
                           din0(11) => s3_b_fwd_11_port, din0(10) => 
                           s3_b_fwd_10_port, din0(9) => s3_b_fwd_9_port, 
                           din0(8) => s3_b_fwd_8_port, din0(7) => 
                           s3_b_fwd_7_port, din0(6) => s3_b_fwd_6_port, din0(5)
                           => s3_b_fwd_5_port, din0(4) => s3_b_fwd_4_port, 
                           din0(3) => s3_b_fwd_3_port, din0(2) => 
                           s3_b_fwd_2_port, din0(1) => s3_b_fwd_1_port, din0(0)
                           => s3_b_fwd_0_port, din1(31) => s3_imm_i_ext_31_port
                           , din1(30) => s3_imm_i_ext_30_port, din1(29) => 
                           s3_imm_i_ext_29_port, din1(28) => 
                           s3_imm_i_ext_28_port, din1(27) => 
                           s3_imm_i_ext_27_port, din1(26) => 
                           s3_imm_i_ext_26_port, din1(25) => 
                           s3_imm_i_ext_25_port, din1(24) => 
                           s3_imm_i_ext_24_port, din1(23) => 
                           s3_imm_i_ext_23_port, din1(22) => 
                           s3_imm_i_ext_22_port, din1(21) => 
                           s3_imm_i_ext_21_port, din1(20) => 
                           s3_imm_i_ext_20_port, din1(19) => 
                           s3_imm_i_ext_19_port, din1(18) => 
                           s3_imm_i_ext_18_port, din1(17) => 
                           s3_imm_i_ext_17_port, din1(16) => 
                           s3_imm_i_ext_16_port, din1(15) => 
                           s3_imm_i_ext_15_port, din1(14) => 
                           s3_imm_i_ext_14_port, din1(13) => 
                           s3_imm_i_ext_13_port, din1(12) => 
                           s3_imm_i_ext_12_port, din1(11) => 
                           s3_imm_i_ext_11_port, din1(10) => 
                           s3_imm_i_ext_10_port, din1(9) => s3_imm_i_ext_9_port
                           , din1(8) => s3_imm_i_ext_8_port, din1(7) => 
                           s3_imm_i_ext_7_port, din1(6) => s3_imm_i_ext_6_port,
                           din1(5) => s3_imm_i_ext_5_port, din1(4) => 
                           s3_imm_i_ext_4_port, din1(3) => s3_imm_i_ext_3_port,
                           din1(2) => s3_imm_i_ext_2_port, din1(1) => 
                           s3_imm_i_ext_1_port, din1(0) => s3_imm_i_ext_0_port,
                           dout(31) => s3_b_sel_31_port, dout(30) => 
                           s3_b_sel_30_port, dout(29) => s3_b_sel_29_port, 
                           dout(28) => s3_b_sel_28_port, dout(27) => 
                           s3_b_sel_27_port, dout(26) => s3_b_sel_26_port, 
                           dout(25) => s3_b_sel_25_port, dout(24) => 
                           s3_b_sel_24_port, dout(23) => s3_b_sel_23_port, 
                           dout(22) => s3_b_sel_22_port, dout(21) => 
                           s3_b_sel_21_port, dout(20) => s3_b_sel_20_port, 
                           dout(19) => s3_b_sel_19_port, dout(18) => 
                           s3_b_sel_18_port, dout(17) => s3_b_sel_17_port, 
                           dout(16) => s3_b_sel_16_port, dout(15) => 
                           s3_b_sel_15_port, dout(14) => s3_b_sel_14_port, 
                           dout(13) => s3_b_sel_13_port, dout(12) => 
                           s3_b_sel_12_port, dout(11) => s3_b_sel_11_port, 
                           dout(10) => s3_b_sel_10_port, dout(9) => 
                           s3_b_sel_9_port, dout(8) => s3_b_sel_8_port, dout(7)
                           => s3_b_sel_7_port, dout(6) => s3_b_sel_6_port, 
                           dout(5) => s3_b_sel_5_port, dout(4) => 
                           s3_b_sel_4_port, dout(3) => s3_b_sel_3_port, dout(2)
                           => s3_b_sel_2_port, dout(1) => s3_b_sel_1_port, 
                           dout(0) => s3_b_sel_0_port);
   ALU0 : Alu_DATA_SIZE32 port map( f(4) => calu(4), f(3) => calu(3), f(2) => 
                           calu(2), f(1) => n93, f(0) => calu(0), a(31) => 
                           s3_a_sel_31_port, a(30) => s3_a_sel_30_port, a(29) 
                           => s3_a_sel_29_port, a(28) => s3_a_sel_28_port, 
                           a(27) => s3_a_sel_27_port, a(26) => s3_a_sel_26_port
                           , a(25) => s3_a_sel_25_port, a(24) => 
                           s3_a_sel_24_port, a(23) => s3_a_sel_23_port, a(22) 
                           => s3_a_sel_22_port, a(21) => s3_a_sel_21_port, 
                           a(20) => s3_a_sel_20_port, a(19) => s3_a_sel_19_port
                           , a(18) => s3_a_sel_18_port, a(17) => 
                           s3_a_sel_17_port, a(16) => s3_a_sel_16_port, a(15) 
                           => s3_a_sel_15_port, a(14) => s3_a_sel_14_port, 
                           a(13) => s3_a_sel_13_port, a(12) => s3_a_sel_12_port
                           , a(11) => s3_a_sel_11_port, a(10) => 
                           s3_a_sel_10_port, a(9) => s3_a_sel_9_port, a(8) => 
                           s3_a_sel_8_port, a(7) => s3_a_sel_7_port, a(6) => 
                           s3_a_sel_6_port, a(5) => s3_a_sel_5_port, a(4) => 
                           s3_a_sel_4_port, a(3) => s3_a_sel_3_port, a(2) => 
                           s3_a_sel_2_port, a(1) => s3_a_sel_1_port, a(0) => 
                           s3_a_sel_0_port, b(31) => s3_b_sel_31_port, b(30) =>
                           s3_b_sel_30_port, b(29) => s3_b_sel_29_port, b(28) 
                           => s3_b_sel_28_port, b(27) => s3_b_sel_27_port, 
                           b(26) => s3_b_sel_26_port, b(25) => s3_b_sel_25_port
                           , b(24) => s3_b_sel_24_port, b(23) => 
                           s3_b_sel_23_port, b(22) => s3_b_sel_22_port, b(21) 
                           => s3_b_sel_21_port, b(20) => s3_b_sel_20_port, 
                           b(19) => s3_b_sel_19_port, b(18) => s3_b_sel_18_port
                           , b(17) => s3_b_sel_17_port, b(16) => 
                           s3_b_sel_16_port, b(15) => s3_b_sel_15_port, b(14) 
                           => s3_b_sel_14_port, b(13) => s3_b_sel_13_port, 
                           b(12) => s3_b_sel_12_port, b(11) => s3_b_sel_11_port
                           , b(10) => s3_b_sel_10_port, b(9) => s3_b_sel_9_port
                           , b(8) => s3_b_sel_8_port, b(7) => s3_b_sel_7_port, 
                           b(6) => s3_b_sel_6_port, b(5) => s3_b_sel_5_port, 
                           b(4) => s3_b_sel_4_port, b(3) => s3_b_sel_3_port, 
                           b(2) => s3_b_sel_2_port, b(1) => s3_b_sel_1_port, 
                           b(0) => s3_b_sel_0_port, o(31) => s3_alu_out_31_port
                           , o(30) => s3_alu_out_30_port, o(29) => 
                           s3_alu_out_29_port, o(28) => s3_alu_out_28_port, 
                           o(27) => s3_alu_out_27_port, o(26) => 
                           s3_alu_out_26_port, o(25) => s3_alu_out_25_port, 
                           o(24) => s3_alu_out_24_port, o(23) => 
                           s3_alu_out_23_port, o(22) => s3_alu_out_22_port, 
                           o(21) => s3_alu_out_21_port, o(20) => 
                           s3_alu_out_20_port, o(19) => s3_alu_out_19_port, 
                           o(18) => s3_alu_out_18_port, o(17) => 
                           s3_alu_out_17_port, o(16) => s3_alu_out_16_port, 
                           o(15) => s3_alu_out_15_port, o(14) => 
                           s3_alu_out_14_port, o(13) => s3_alu_out_13_port, 
                           o(12) => s3_alu_out_12_port, o(11) => 
                           s3_alu_out_11_port, o(10) => s3_alu_out_10_port, 
                           o(9) => s3_alu_out_9_port, o(8) => s3_alu_out_8_port
                           , o(7) => s3_alu_out_7_port, o(6) => 
                           s3_alu_out_6_port, o(5) => s3_alu_out_5_port, o(4) 
                           => s3_alu_out_4_port, o(3) => s3_alu_out_3_port, 
                           o(2) => s3_alu_out_2_port, o(1) => s3_alu_out_1_port
                           , o(0) => s3_alu_out_0_port);
   MUL0 : Mul_DATA_SIZE16_STAGE10 port map( rst => n111, clk => clk, en => 
                           sig_mul_port, lock => sig_ral_port, sign => 
                           s3_mul_sign, a(15) => s3_a_sel_15_port, a(14) => 
                           s3_a_sel_14_port, a(13) => s3_a_sel_13_port, a(12) 
                           => s3_a_sel_12_port, a(11) => s3_a_sel_11_port, 
                           a(10) => s3_a_sel_10_port, a(9) => s3_a_sel_9_port, 
                           a(8) => s3_a_sel_8_port, a(7) => s3_a_sel_7_port, 
                           a(6) => s3_a_sel_6_port, a(5) => s3_a_sel_5_port, 
                           a(4) => s3_a_sel_4_port, a(3) => s3_a_sel_3_port, 
                           a(2) => s3_a_sel_2_port, a(1) => s3_a_sel_1_port, 
                           a(0) => s3_a_sel_0_port, b(15) => s3_b_sel_15_port, 
                           b(14) => s3_b_sel_14_port, b(13) => s3_b_sel_13_port
                           , b(12) => s3_b_sel_12_port, b(11) => 
                           s3_b_sel_11_port, b(10) => s3_b_sel_10_port, b(9) =>
                           s3_b_sel_9_port, b(8) => s3_b_sel_8_port, b(7) => 
                           s3_b_sel_7_port, b(6) => s3_b_sel_6_port, b(5) => 
                           s3_b_sel_5_port, b(4) => s3_b_sel_4_port, b(3) => 
                           s3_b_sel_3_port, b(2) => s3_b_sel_2_port, b(1) => 
                           s3_b_sel_1_port, b(0) => n90, o(31) => 
                           s3_mul_out_31_port, o(30) => s3_mul_out_30_port, 
                           o(29) => s3_mul_out_29_port, o(28) => 
                           s3_mul_out_28_port, o(27) => s3_mul_out_27_port, 
                           o(26) => s3_mul_out_26_port, o(25) => 
                           s3_mul_out_25_port, o(24) => s3_mul_out_24_port, 
                           o(23) => s3_mul_out_23_port, o(22) => 
                           s3_mul_out_22_port, o(21) => s3_mul_out_21_port, 
                           o(20) => s3_mul_out_20_port, o(19) => 
                           s3_mul_out_19_port, o(18) => s3_mul_out_18_port, 
                           o(17) => s3_mul_out_17_port, o(16) => 
                           s3_mul_out_16_port, o(15) => s3_mul_out_15_port, 
                           o(14) => s3_mul_out_14_port, o(13) => 
                           s3_mul_out_13_port, o(12) => s3_mul_out_12_port, 
                           o(11) => s3_mul_out_11_port, o(10) => 
                           s3_mul_out_10_port, o(9) => s3_mul_out_9_port, o(8) 
                           => s3_mul_out_8_port, o(7) => s3_mul_out_7_port, 
                           o(6) => s3_mul_out_6_port, o(5) => s3_mul_out_5_port
                           , o(4) => s3_mul_out_4_port, o(3) => 
                           s3_mul_out_3_port, o(2) => s3_mul_out_2_port, o(1) 
                           => s3_mul_out_1_port, o(0) => s3_mul_out_0_port);
   DIV0 : Div_DATA_SIZE32_DIV_STAGE34_SQRT_STAGE18 port map( rst => n111, clk 
                           => clk, en => s3_exe_sel_1_port, lock => 
                           sig_ral_port, sign => s3_div_sign, func => n104, 
                           a(31) => s3_a_sel_31_port, a(30) => s3_a_sel_30_port
                           , a(29) => s3_a_sel_29_port, a(28) => 
                           s3_a_sel_28_port, a(27) => s3_a_sel_27_port, a(26) 
                           => s3_a_sel_26_port, a(25) => s3_a_sel_25_port, 
                           a(24) => s3_a_sel_24_port, a(23) => s3_a_sel_23_port
                           , a(22) => s3_a_sel_22_port, a(21) => 
                           s3_a_sel_21_port, a(20) => s3_a_sel_20_port, a(19) 
                           => s3_a_sel_19_port, a(18) => s3_a_sel_18_port, 
                           a(17) => s3_a_sel_17_port, a(16) => s3_a_sel_16_port
                           , a(15) => s3_a_sel_15_port, a(14) => 
                           s3_a_sel_14_port, a(13) => s3_a_sel_13_port, a(12) 
                           => s3_a_sel_12_port, a(11) => s3_a_sel_11_port, 
                           a(10) => s3_a_sel_10_port, a(9) => s3_a_sel_9_port, 
                           a(8) => s3_a_sel_8_port, a(7) => s3_a_sel_7_port, 
                           a(6) => s3_a_sel_6_port, a(5) => s3_a_sel_5_port, 
                           a(4) => s3_a_sel_4_port, a(3) => s3_a_sel_3_port, 
                           a(2) => s3_a_sel_2_port, a(1) => s3_a_sel_1_port, 
                           a(0) => s3_a_sel_0_port, b(31) => s3_b_sel_31_port, 
                           b(30) => s3_b_sel_30_port, b(29) => s3_b_sel_29_port
                           , b(28) => s3_b_sel_28_port, b(27) => 
                           s3_b_sel_27_port, b(26) => s3_b_sel_26_port, b(25) 
                           => s3_b_sel_25_port, b(24) => s3_b_sel_24_port, 
                           b(23) => s3_b_sel_23_port, b(22) => s3_b_sel_22_port
                           , b(21) => s3_b_sel_21_port, b(20) => 
                           s3_b_sel_20_port, b(19) => s3_b_sel_19_port, b(18) 
                           => s3_b_sel_18_port, b(17) => s3_b_sel_17_port, 
                           b(16) => s3_b_sel_16_port, b(15) => s3_b_sel_15_port
                           , b(14) => s3_b_sel_14_port, b(13) => 
                           s3_b_sel_13_port, b(12) => s3_b_sel_12_port, b(11) 
                           => s3_b_sel_11_port, b(10) => s3_b_sel_10_port, b(9)
                           => s3_b_sel_9_port, b(8) => s3_b_sel_8_port, b(7) =>
                           s3_b_sel_7_port, b(6) => s3_b_sel_6_port, b(5) => 
                           s3_b_sel_5_port, b(4) => s3_b_sel_4_port, b(3) => 
                           s3_b_sel_3_port, b(2) => s3_b_sel_2_port, b(1) => 
                           s3_b_sel_1_port, b(0) => n87, o(31) => 
                           s3_div_out_31_port, o(30) => s3_div_out_30_port, 
                           o(29) => s3_div_out_29_port, o(28) => 
                           s3_div_out_28_port, o(27) => s3_div_out_27_port, 
                           o(26) => s3_div_out_26_port, o(25) => 
                           s3_div_out_25_port, o(24) => s3_div_out_24_port, 
                           o(23) => s3_div_out_23_port, o(22) => 
                           s3_div_out_22_port, o(21) => s3_div_out_21_port, 
                           o(20) => s3_div_out_20_port, o(19) => 
                           s3_div_out_19_port, o(18) => s3_div_out_18_port, 
                           o(17) => s3_div_out_17_port, o(16) => 
                           s3_div_out_16_port, o(15) => s3_div_out_15_port, 
                           o(14) => s3_div_out_14_port, o(13) => 
                           s3_div_out_13_port, o(12) => s3_div_out_12_port, 
                           o(11) => s3_div_out_11_port, o(10) => 
                           s3_div_out_10_port, o(9) => s3_div_out_9_port, o(8) 
                           => s3_div_out_8_port, o(7) => s3_div_out_7_port, 
                           o(6) => s3_div_out_6_port, o(5) => s3_div_out_5_port
                           , o(4) => s3_div_out_4_port, o(3) => 
                           s3_div_out_3_port, o(2) => s3_div_out_2_port, o(1) 
                           => s3_div_out_1_port, o(0) => s3_div_out_0_port);
   MUXEXE : Mux4_DATA_SIZE32 port map( sel(1) => s3_exe_sel_1_port, sel(0) => 
                           sig_mul_port, din0(31) => s3_alu_out_31_port, 
                           din0(30) => s3_alu_out_30_port, din0(29) => 
                           s3_alu_out_29_port, din0(28) => s3_alu_out_28_port, 
                           din0(27) => s3_alu_out_27_port, din0(26) => 
                           s3_alu_out_26_port, din0(25) => s3_alu_out_25_port, 
                           din0(24) => s3_alu_out_24_port, din0(23) => 
                           s3_alu_out_23_port, din0(22) => s3_alu_out_22_port, 
                           din0(21) => s3_alu_out_21_port, din0(20) => 
                           s3_alu_out_20_port, din0(19) => s3_alu_out_19_port, 
                           din0(18) => s3_alu_out_18_port, din0(17) => 
                           s3_alu_out_17_port, din0(16) => s3_alu_out_16_port, 
                           din0(15) => s3_alu_out_15_port, din0(14) => 
                           s3_alu_out_14_port, din0(13) => s3_alu_out_13_port, 
                           din0(12) => s3_alu_out_12_port, din0(11) => 
                           s3_alu_out_11_port, din0(10) => s3_alu_out_10_port, 
                           din0(9) => s3_alu_out_9_port, din0(8) => 
                           s3_alu_out_8_port, din0(7) => s3_alu_out_7_port, 
                           din0(6) => s3_alu_out_6_port, din0(5) => 
                           s3_alu_out_5_port, din0(4) => s3_alu_out_4_port, 
                           din0(3) => s3_alu_out_3_port, din0(2) => 
                           s3_alu_out_2_port, din0(1) => s3_alu_out_1_port, 
                           din0(0) => s3_alu_out_0_port, din1(31) => 
                           s3_mul_out_31_port, din1(30) => s3_mul_out_30_port, 
                           din1(29) => s3_mul_out_29_port, din1(28) => 
                           s3_mul_out_28_port, din1(27) => s3_mul_out_27_port, 
                           din1(26) => s3_mul_out_26_port, din1(25) => 
                           s3_mul_out_25_port, din1(24) => s3_mul_out_24_port, 
                           din1(23) => s3_mul_out_23_port, din1(22) => 
                           s3_mul_out_22_port, din1(21) => s3_mul_out_21_port, 
                           din1(20) => s3_mul_out_20_port, din1(19) => 
                           s3_mul_out_19_port, din1(18) => s3_mul_out_18_port, 
                           din1(17) => s3_mul_out_17_port, din1(16) => 
                           s3_mul_out_16_port, din1(15) => s3_mul_out_15_port, 
                           din1(14) => s3_mul_out_14_port, din1(13) => 
                           s3_mul_out_13_port, din1(12) => s3_mul_out_12_port, 
                           din1(11) => s3_mul_out_11_port, din1(10) => 
                           s3_mul_out_10_port, din1(9) => s3_mul_out_9_port, 
                           din1(8) => s3_mul_out_8_port, din1(7) => 
                           s3_mul_out_7_port, din1(6) => s3_mul_out_6_port, 
                           din1(5) => s3_mul_out_5_port, din1(4) => 
                           s3_mul_out_4_port, din1(3) => s3_mul_out_3_port, 
                           din1(2) => s3_mul_out_2_port, din1(1) => 
                           s3_mul_out_1_port, din1(0) => s3_mul_out_0_port, 
                           din2(31) => s3_div_out_31_port, din2(30) => 
                           s3_div_out_30_port, din2(29) => s3_div_out_29_port, 
                           din2(28) => s3_div_out_28_port, din2(27) => 
                           s3_div_out_27_port, din2(26) => s3_div_out_26_port, 
                           din2(25) => s3_div_out_25_port, din2(24) => 
                           s3_div_out_24_port, din2(23) => s3_div_out_23_port, 
                           din2(22) => s3_div_out_22_port, din2(21) => 
                           s3_div_out_21_port, din2(20) => s3_div_out_20_port, 
                           din2(19) => s3_div_out_19_port, din2(18) => 
                           s3_div_out_18_port, din2(17) => s3_div_out_17_port, 
                           din2(16) => s3_div_out_16_port, din2(15) => 
                           s3_div_out_15_port, din2(14) => s3_div_out_14_port, 
                           din2(13) => s3_div_out_13_port, din2(12) => 
                           s3_div_out_12_port, din2(11) => s3_div_out_11_port, 
                           din2(10) => s3_div_out_10_port, din2(9) => 
                           s3_div_out_9_port, din2(8) => s3_div_out_8_port, 
                           din2(7) => s3_div_out_7_port, din2(6) => 
                           s3_div_out_6_port, din2(5) => s3_div_out_5_port, 
                           din2(4) => s3_div_out_4_port, din2(3) => 
                           s3_div_out_3_port, din2(2) => s3_div_out_2_port, 
                           din2(1) => s3_div_out_1_port, din2(0) => 
                           s3_div_out_0_port, din3(31) => X_Logic0_port, 
                           din3(30) => X_Logic0_port, din3(29) => X_Logic0_port
                           , din3(28) => X_Logic0_port, din3(27) => 
                           X_Logic0_port, din3(26) => X_Logic0_port, din3(25) 
                           => X_Logic0_port, din3(24) => X_Logic0_port, 
                           din3(23) => X_Logic0_port, din3(22) => X_Logic0_port
                           , din3(21) => X_Logic0_port, din3(20) => 
                           X_Logic0_port, din3(19) => X_Logic0_port, din3(18) 
                           => X_Logic0_port, din3(17) => X_Logic0_port, 
                           din3(16) => X_Logic0_port, din3(15) => X_Logic0_port
                           , din3(14) => X_Logic0_port, din3(13) => 
                           X_Logic0_port, din3(12) => X_Logic0_port, din3(11) 
                           => X_Logic0_port, din3(10) => X_Logic0_port, din3(9)
                           => X_Logic0_port, din3(8) => X_Logic0_port, din3(7) 
                           => X_Logic0_port, din3(6) => X_Logic0_port, din3(5) 
                           => X_Logic0_port, din3(4) => X_Logic0_port, din3(3) 
                           => X_Logic0_port, din3(2) => X_Logic0_port, din3(1) 
                           => X_Logic0_port, din3(0) => X_Logic0_port, dout(31)
                           => s3_exe_out_31_port, dout(30) => 
                           s3_exe_out_30_port, dout(29) => s3_exe_out_29_port, 
                           dout(28) => s3_exe_out_28_port, dout(27) => 
                           s3_exe_out_27_port, dout(26) => s3_exe_out_26_port, 
                           dout(25) => s3_exe_out_25_port, dout(24) => 
                           s3_exe_out_24_port, dout(23) => s3_exe_out_23_port, 
                           dout(22) => s3_exe_out_22_port, dout(21) => 
                           s3_exe_out_21_port, dout(20) => s3_exe_out_20_port, 
                           dout(19) => s3_exe_out_19_port, dout(18) => 
                           s3_exe_out_18_port, dout(17) => s3_exe_out_17_port, 
                           dout(16) => s3_exe_out_16_port, dout(15) => 
                           s3_exe_out_15_port, dout(14) => s3_exe_out_14_port, 
                           dout(13) => s3_exe_out_13_port, dout(12) => 
                           s3_exe_out_12_port, dout(11) => s3_exe_out_11_port, 
                           dout(10) => s3_exe_out_10_port, dout(9) => 
                           s3_exe_out_9_port, dout(8) => s3_exe_out_8_port, 
                           dout(7) => s3_exe_out_7_port, dout(6) => 
                           s3_exe_out_6_port, dout(5) => s3_exe_out_5_port, 
                           dout(4) => s3_exe_out_4_port, dout(3) => 
                           s3_exe_out_3_port, dout(2) => s3_exe_out_2_port, 
                           dout(1) => s3_exe_out_1_port, dout(0) => 
                           s3_exe_out_0_port);
   REG_ALU : Reg_DATA_SIZE32_7 port map( rst => n111, en => cw(10), clk => clk,
                           din(31) => s3_exe_out_31_port, din(30) => 
                           s3_exe_out_30_port, din(29) => s3_exe_out_29_port, 
                           din(28) => s3_exe_out_28_port, din(27) => 
                           s3_exe_out_27_port, din(26) => s3_exe_out_26_port, 
                           din(25) => s3_exe_out_25_port, din(24) => 
                           s3_exe_out_24_port, din(23) => s3_exe_out_23_port, 
                           din(22) => s3_exe_out_22_port, din(21) => 
                           s3_exe_out_21_port, din(20) => s3_exe_out_20_port, 
                           din(19) => s3_exe_out_19_port, din(18) => 
                           s3_exe_out_18_port, din(17) => s3_exe_out_17_port, 
                           din(16) => s3_exe_out_16_port, din(15) => 
                           s3_exe_out_15_port, din(14) => s3_exe_out_14_port, 
                           din(13) => s3_exe_out_13_port, din(12) => 
                           s3_exe_out_12_port, din(11) => s3_exe_out_11_port, 
                           din(10) => s3_exe_out_10_port, din(9) => 
                           s3_exe_out_9_port, din(8) => s3_exe_out_8_port, 
                           din(7) => s3_exe_out_7_port, din(6) => 
                           s3_exe_out_6_port, din(5) => s3_exe_out_5_port, 
                           din(4) => s3_exe_out_4_port, din(3) => 
                           s3_exe_out_3_port, din(2) => s3_exe_out_2_port, 
                           din(1) => s3_exe_out_1_port, din(0) => 
                           s3_exe_out_0_port, dout(31) => data_addr_31_port, 
                           dout(30) => data_addr_30_port, dout(29) => 
                           data_addr_29_port, dout(28) => data_addr_28_port, 
                           dout(27) => data_addr_27_port, dout(26) => 
                           data_addr_26_port, dout(25) => data_addr_25_port, 
                           dout(24) => data_addr_24_port, dout(23) => 
                           data_addr_23_port, dout(22) => data_addr_22_port, 
                           dout(21) => data_addr_21_port, dout(20) => 
                           data_addr_20_port, dout(19) => data_addr_19_port, 
                           dout(18) => data_addr_18_port, dout(17) => 
                           data_addr_17_port, dout(16) => data_addr_16_port, 
                           dout(15) => data_addr_15_port, dout(14) => 
                           data_addr_14_port, dout(13) => data_addr_13_port, 
                           dout(12) => data_addr_12_port, dout(11) => 
                           data_addr_11_port, dout(10) => data_addr_10_port, 
                           dout(9) => data_addr_9_port, dout(8) => 
                           data_addr_8_port, dout(7) => data_addr_7_port, 
                           dout(6) => data_addr_6_port, dout(5) => 
                           data_addr_5_port, dout(4) => data_addr_4_port, 
                           dout(3) => data_addr_3_port, dout(2) => 
                           data_addr_2_port, dout(1) => data_addr_1_port, 
                           dout(0) => data_addr_0_port);
   REG_BB : Reg_DATA_SIZE32_6 port map( rst => n111, en => cw(10), clk => clk, 
                           din(31) => s3_b_fwd_31_port, din(30) => 
                           s3_b_fwd_30_port, din(29) => s3_b_fwd_29_port, 
                           din(28) => s3_b_fwd_28_port, din(27) => 
                           s3_b_fwd_27_port, din(26) => s3_b_fwd_26_port, 
                           din(25) => s3_b_fwd_25_port, din(24) => 
                           s3_b_fwd_24_port, din(23) => s3_b_fwd_23_port, 
                           din(22) => s3_b_fwd_22_port, din(21) => 
                           s3_b_fwd_21_port, din(20) => s3_b_fwd_20_port, 
                           din(19) => s3_b_fwd_19_port, din(18) => 
                           s3_b_fwd_18_port, din(17) => s3_b_fwd_17_port, 
                           din(16) => s3_b_fwd_16_port, din(15) => 
                           s3_b_fwd_15_port, din(14) => s3_b_fwd_14_port, 
                           din(13) => s3_b_fwd_13_port, din(12) => 
                           s3_b_fwd_12_port, din(11) => s3_b_fwd_11_port, 
                           din(10) => s3_b_fwd_10_port, din(9) => 
                           s3_b_fwd_9_port, din(8) => s3_b_fwd_8_port, din(7) 
                           => s3_b_fwd_7_port, din(6) => s3_b_fwd_6_port, 
                           din(5) => s3_b_fwd_5_port, din(4) => s3_b_fwd_4_port
                           , din(3) => s3_b_fwd_3_port, din(2) => 
                           s3_b_fwd_2_port, din(1) => s3_b_fwd_1_port, din(0) 
                           => s3_b_fwd_0_port, dout(31) => s4_b_fwd_31_port, 
                           dout(30) => s4_b_fwd_30_port, dout(29) => 
                           s4_b_fwd_29_port, dout(28) => s4_b_fwd_28_port, 
                           dout(27) => s4_b_fwd_27_port, dout(26) => 
                           s4_b_fwd_26_port, dout(25) => s4_b_fwd_25_port, 
                           dout(24) => s4_b_fwd_24_port, dout(23) => 
                           s4_b_fwd_23_port, dout(22) => s4_b_fwd_22_port, 
                           dout(21) => s4_b_fwd_21_port, dout(20) => 
                           s4_b_fwd_20_port, dout(19) => s4_b_fwd_19_port, 
                           dout(18) => s4_b_fwd_18_port, dout(17) => 
                           s4_b_fwd_17_port, dout(16) => s4_b_fwd_16_port, 
                           dout(15) => s4_b_fwd_15_port, dout(14) => 
                           s4_b_fwd_14_port, dout(13) => s4_b_fwd_13_port, 
                           dout(12) => s4_b_fwd_12_port, dout(11) => 
                           s4_b_fwd_11_port, dout(10) => s4_b_fwd_10_port, 
                           dout(9) => s4_b_fwd_9_port, dout(8) => 
                           s4_b_fwd_8_port, dout(7) => s4_b_fwd_7_port, dout(6)
                           => s4_b_fwd_6_port, dout(5) => s4_b_fwd_5_port, 
                           dout(4) => s4_b_fwd_4_port, dout(3) => 
                           s4_b_fwd_3_port, dout(2) => s4_b_fwd_2_port, dout(1)
                           => s4_b_fwd_1_port, dout(0) => s4_b_fwd_0_port);
   REG_B_ADDR_3 : Reg_DATA_SIZE5_4 port map( rst => n110, en => cw(10), clk => 
                           clk, din(4) => s3_rd2_addr_4_port, din(3) => 
                           s3_rd2_addr_3_port, din(2) => s3_rd2_addr_2_port, 
                           din(1) => s3_rd2_addr_1_port, din(0) => 
                           s3_rd2_addr_0_port, dout(4) => s4_rd2_addr_4_port, 
                           dout(3) => s4_rd2_addr_3_port, dout(2) => 
                           s4_rd2_addr_2_port, dout(1) => s4_rd2_addr_1_port, 
                           dout(0) => s4_rd2_addr_0_port);
   REG_WR3 : Reg_DATA_SIZE5_3 port map( rst => n110, en => cw(10), clk => clk, 
                           din(4) => s3_wr_addr_4_port, din(3) => 
                           s3_wr_addr_3_port, din(2) => s3_wr_addr_2_port, 
                           din(1) => s3_wr_addr_1_port, din(0) => 
                           s3_wr_addr_0_port, dout(4) => s4_wr_addr_4_port, 
                           dout(3) => s4_wr_addr_3_port, dout(2) => 
                           s4_wr_addr_2_port, dout(1) => s4_wr_addr_1_port, 
                           dout(0) => s4_wr_addr_0_port);
   REG_OPRD_A_WAIT : Reg_DATA_SIZE32_5 port map( rst => n111, en => 
                           X_Logic1_port, clk => clk, din(31) => 
                           s3_a_sel_31_port, din(30) => s3_a_sel_30_port, 
                           din(29) => s3_a_sel_29_port, din(28) => 
                           s3_a_sel_28_port, din(27) => s3_a_sel_27_port, 
                           din(26) => s3_a_sel_26_port, din(25) => 
                           s3_a_sel_25_port, din(24) => s3_a_sel_24_port, 
                           din(23) => s3_a_sel_23_port, din(22) => 
                           s3_a_sel_22_port, din(21) => s3_a_sel_21_port, 
                           din(20) => s3_a_sel_20_port, din(19) => 
                           s3_a_sel_19_port, din(18) => s3_a_sel_18_port, 
                           din(17) => s3_a_sel_17_port, din(16) => 
                           s3_a_sel_16_port, din(15) => s3_a_sel_15_port, 
                           din(14) => s3_a_sel_14_port, din(13) => 
                           s3_a_sel_13_port, din(12) => s3_a_sel_12_port, 
                           din(11) => s3_a_sel_11_port, din(10) => 
                           s3_a_sel_10_port, din(9) => s3_a_sel_9_port, din(8) 
                           => s3_a_sel_8_port, din(7) => s3_a_sel_7_port, 
                           din(6) => s3_a_sel_6_port, din(5) => s3_a_sel_5_port
                           , din(4) => s3_a_sel_4_port, din(3) => 
                           s3_a_sel_3_port, din(2) => s3_a_sel_2_port, din(1) 
                           => s3_a_sel_1_port, din(0) => s3_a_sel_0_port, 
                           dout(31) => s4_a_31_port, dout(30) => s4_a_30_port, 
                           dout(29) => s4_a_29_port, dout(28) => s4_a_28_port, 
                           dout(27) => s4_a_27_port, dout(26) => s4_a_26_port, 
                           dout(25) => s4_a_25_port, dout(24) => s4_a_24_port, 
                           dout(23) => s4_a_23_port, dout(22) => s4_a_22_port, 
                           dout(21) => s4_a_21_port, dout(20) => s4_a_20_port, 
                           dout(19) => s4_a_19_port, dout(18) => s4_a_18_port, 
                           dout(17) => s4_a_17_port, dout(16) => s4_a_16_port, 
                           dout(15) => s4_a_15_port, dout(14) => s4_a_14_port, 
                           dout(13) => s4_a_13_port, dout(12) => s4_a_12_port, 
                           dout(11) => s4_a_11_port, dout(10) => s4_a_10_port, 
                           dout(9) => s4_a_9_port, dout(8) => s4_a_8_port, 
                           dout(7) => s4_a_7_port, dout(6) => s4_a_6_port, 
                           dout(5) => s4_a_5_port, dout(4) => s4_a_4_port, 
                           dout(3) => s4_a_3_port, dout(2) => s4_a_2_port, 
                           dout(1) => s4_a_1_port, dout(0) => s4_a_0_port);
   REG_OPRD_B_WAIT : Reg_DATA_SIZE32_4 port map( rst => n111, en => 
                           X_Logic1_port, clk => clk, din(31) => 
                           s3_b_sel_31_port, din(30) => s3_b_sel_30_port, 
                           din(29) => s3_b_sel_29_port, din(28) => 
                           s3_b_sel_28_port, din(27) => s3_b_sel_27_port, 
                           din(26) => s3_b_sel_26_port, din(25) => 
                           s3_b_sel_25_port, din(24) => s3_b_sel_24_port, 
                           din(23) => s3_b_sel_23_port, din(22) => 
                           s3_b_sel_22_port, din(21) => s3_b_sel_21_port, 
                           din(20) => s3_b_sel_20_port, din(19) => 
                           s3_b_sel_19_port, din(18) => s3_b_sel_18_port, 
                           din(17) => s3_b_sel_17_port, din(16) => 
                           s3_b_sel_16_port, din(15) => s3_b_sel_15_port, 
                           din(14) => s3_b_sel_14_port, din(13) => 
                           s3_b_sel_13_port, din(12) => s3_b_sel_12_port, 
                           din(11) => s3_b_sel_11_port, din(10) => 
                           s3_b_sel_10_port, din(9) => s3_b_sel_9_port, din(8) 
                           => s3_b_sel_8_port, din(7) => s3_b_sel_7_port, 
                           din(6) => s3_b_sel_6_port, din(5) => s3_b_sel_5_port
                           , din(4) => s3_b_sel_4_port, din(3) => 
                           s3_b_sel_3_port, din(2) => s3_b_sel_2_port, din(1) 
                           => s3_b_sel_1_port, din(0) => n90, dout(31) => 
                           s4_b_31_port, dout(30) => s4_b_30_port, dout(29) => 
                           s4_b_29_port, dout(28) => s4_b_28_port, dout(27) => 
                           s4_b_27_port, dout(26) => s4_b_26_port, dout(25) => 
                           s4_b_25_port, dout(24) => s4_b_24_port, dout(23) => 
                           s4_b_23_port, dout(22) => s4_b_22_port, dout(21) => 
                           s4_b_21_port, dout(20) => s4_b_20_port, dout(19) => 
                           s4_b_19_port, dout(18) => s4_b_18_port, dout(17) => 
                           s4_b_17_port, dout(16) => s4_b_16_port, dout(15) => 
                           s4_b_15_port, dout(14) => s4_b_14_port, dout(13) => 
                           s4_b_13_port, dout(12) => s4_b_12_port, dout(11) => 
                           s4_b_11_port, dout(10) => s4_b_10_port, dout(9) => 
                           s4_b_9_port, dout(8) => s4_b_8_port, dout(7) => 
                           s4_b_7_port, dout(6) => s4_b_6_port, dout(5) => 
                           s4_b_5_port, dout(4) => s4_b_4_port, dout(3) => 
                           s4_b_3_port, dout(2) => s4_b_2_port, dout(1) => 
                           s4_b_1_port, dout(0) => s4_b_0_port);
   FWDMUX_BB : FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_1 port map( reg_c(31) => 
                           s4_b_fwd_31_port, reg_c(30) => s4_b_fwd_30_port, 
                           reg_c(29) => s4_b_fwd_29_port, reg_c(28) => 
                           s4_b_fwd_28_port, reg_c(27) => s4_b_fwd_27_port, 
                           reg_c(26) => s4_b_fwd_26_port, reg_c(25) => 
                           s4_b_fwd_25_port, reg_c(24) => s4_b_fwd_24_port, 
                           reg_c(23) => s4_b_fwd_23_port, reg_c(22) => 
                           s4_b_fwd_22_port, reg_c(21) => s4_b_fwd_21_port, 
                           reg_c(20) => s4_b_fwd_20_port, reg_c(19) => 
                           s4_b_fwd_19_port, reg_c(18) => s4_b_fwd_18_port, 
                           reg_c(17) => s4_b_fwd_17_port, reg_c(16) => 
                           s4_b_fwd_16_port, reg_c(15) => s4_b_fwd_15_port, 
                           reg_c(14) => s4_b_fwd_14_port, reg_c(13) => 
                           s4_b_fwd_13_port, reg_c(12) => s4_b_fwd_12_port, 
                           reg_c(11) => s4_b_fwd_11_port, reg_c(10) => 
                           s4_b_fwd_10_port, reg_c(9) => s4_b_fwd_9_port, 
                           reg_c(8) => s4_b_fwd_8_port, reg_c(7) => 
                           s4_b_fwd_7_port, reg_c(6) => s4_b_fwd_6_port, 
                           reg_c(5) => s4_b_fwd_5_port, reg_c(4) => 
                           s4_b_fwd_4_port, reg_c(3) => s4_b_fwd_3_port, 
                           reg_c(2) => s4_b_fwd_2_port, reg_c(1) => 
                           s4_b_fwd_1_port, reg_c(0) => s4_b_fwd_0_port, 
                           reg_f(31) => s5_result_31_port, reg_f(30) => 
                           s5_result_30_port, reg_f(29) => s5_result_29_port, 
                           reg_f(28) => s5_result_28_port, reg_f(27) => 
                           s5_result_27_port, reg_f(26) => s5_result_26_port, 
                           reg_f(25) => s5_result_25_port, reg_f(24) => 
                           s5_result_24_port, reg_f(23) => s5_result_23_port, 
                           reg_f(22) => s5_result_22_port, reg_f(21) => 
                           s5_result_21_port, reg_f(20) => s5_result_20_port, 
                           reg_f(19) => s5_result_19_port, reg_f(18) => 
                           s5_result_18_port, reg_f(17) => s5_result_17_port, 
                           reg_f(16) => s5_result_16_port, reg_f(15) => 
                           s5_result_15_port, reg_f(14) => s5_result_14_port, 
                           reg_f(13) => s5_result_13_port, reg_f(12) => 
                           s5_result_12_port, reg_f(11) => s5_result_11_port, 
                           reg_f(10) => s5_result_10_port, reg_f(9) => 
                           s5_result_9_port, reg_f(8) => s5_result_8_port, 
                           reg_f(7) => s5_result_7_port, reg_f(6) => 
                           s5_result_6_port, reg_f(5) => s5_result_5_port, 
                           reg_f(4) => s5_result_4_port, reg_f(3) => 
                           s5_result_3_port, reg_f(2) => s5_result_2_port, 
                           reg_f(1) => s5_result_1_port, reg_f(0) => 
                           s5_result_0_port, reg_ff(31) => s6_result_31_port, 
                           reg_ff(30) => s6_result_30_port, reg_ff(29) => 
                           s6_result_29_port, reg_ff(28) => s6_result_28_port, 
                           reg_ff(27) => s6_result_27_port, reg_ff(26) => 
                           s6_result_26_port, reg_ff(25) => s6_result_25_port, 
                           reg_ff(24) => s6_result_24_port, reg_ff(23) => 
                           s6_result_23_port, reg_ff(22) => s6_result_22_port, 
                           reg_ff(21) => s6_result_21_port, reg_ff(20) => 
                           s6_result_20_port, reg_ff(19) => s6_result_19_port, 
                           reg_ff(18) => s6_result_18_port, reg_ff(17) => 
                           s6_result_17_port, reg_ff(16) => s6_result_16_port, 
                           reg_ff(15) => s6_result_15_port, reg_ff(14) => 
                           s6_result_14_port, reg_ff(13) => s6_result_13_port, 
                           reg_ff(12) => s6_result_12_port, reg_ff(11) => 
                           s6_result_11_port, reg_ff(10) => s6_result_10_port, 
                           reg_ff(9) => s6_result_9_port, reg_ff(8) => 
                           s6_result_8_port, reg_ff(7) => s6_result_7_port, 
                           reg_ff(6) => s6_result_6_port, reg_ff(5) => 
                           s6_result_5_port, reg_ff(4) => s6_result_4_port, 
                           reg_ff(3) => s6_result_3_port, reg_ff(2) => 
                           s6_result_2_port, reg_ff(1) => s6_result_1_port, 
                           reg_ff(0) => s6_result_0_port, addr_c(4) => 
                           s4_rd2_addr_4_port, addr_c(3) => s4_rd2_addr_3_port,
                           addr_c(2) => s4_rd2_addr_2_port, addr_c(1) => 
                           s4_rd2_addr_1_port, addr_c(0) => s4_rd2_addr_0_port,
                           addr_f(4) => s5_wr_addr_4_port, addr_f(3) => 
                           s5_wr_addr_3_port, addr_f(2) => s5_wr_addr_2_port, 
                           addr_f(1) => s5_wr_addr_1_port, addr_f(0) => 
                           s5_wr_addr_0_port, addr_ff(4) => s6_wr_addr_4_port, 
                           addr_ff(3) => s6_wr_addr_3_port, addr_ff(2) => 
                           s6_wr_addr_2_port, addr_ff(1) => s6_wr_addr_1_port, 
                           addr_ff(0) => s6_wr_addr_0_port, valid_f => cw(19), 
                           valid_ff => s6_en_wb, dirty_f => X_Logic0_port, 
                           dirty_ff => X_Logic0_port, en => cw(14), output(31) 
                           => data_o_val(31), output(30) => data_o_val(30), 
                           output(29) => data_o_val(29), output(28) => 
                           data_o_val(28), output(27) => data_o_val(27), 
                           output(26) => data_o_val(26), output(25) => 
                           data_o_val(25), output(24) => data_o_val(24), 
                           output(23) => data_o_val(23), output(22) => 
                           data_o_val(22), output(21) => data_o_val(21), 
                           output(20) => data_o_val(20), output(19) => 
                           data_o_val(19), output(18) => data_o_val(18), 
                           output(17) => data_o_val(17), output(16) => 
                           data_o_val(16), output(15) => data_o_val(15), 
                           output(14) => data_o_val(14), output(13) => 
                           data_o_val(13), output(12) => data_o_val(12), 
                           output(11) => data_o_val(11), output(10) => 
                           data_o_val(10), output(9) => data_o_val(9), 
                           output(8) => data_o_val(8), output(7) => 
                           data_o_val(7), output(6) => data_o_val(6), output(5)
                           => data_o_val(5), output(4) => data_o_val(4), 
                           output(3) => data_o_val(3), output(2) => 
                           data_o_val(2), output(1) => data_o_val(1), output(0)
                           => data_o_val(0), match_dirty_f => net1283, 
                           match_dirty_ff => net1284);
   MUX_RESULT : Mux_DATA_SIZE32_2 port map( sel => cw(15), din0(31) => 
                           data_addr_31_port, din0(30) => data_addr_30_port, 
                           din0(29) => data_addr_29_port, din0(28) => 
                           data_addr_28_port, din0(27) => data_addr_27_port, 
                           din0(26) => data_addr_26_port, din0(25) => 
                           data_addr_25_port, din0(24) => data_addr_24_port, 
                           din0(23) => data_addr_23_port, din0(22) => 
                           data_addr_22_port, din0(21) => data_addr_21_port, 
                           din0(20) => data_addr_20_port, din0(19) => 
                           data_addr_19_port, din0(18) => data_addr_18_port, 
                           din0(17) => data_addr_17_port, din0(16) => 
                           data_addr_16_port, din0(15) => data_addr_15_port, 
                           din0(14) => data_addr_14_port, din0(13) => 
                           data_addr_13_port, din0(12) => data_addr_12_port, 
                           din0(11) => data_addr_11_port, din0(10) => 
                           data_addr_10_port, din0(9) => data_addr_9_port, 
                           din0(8) => data_addr_8_port, din0(7) => 
                           data_addr_7_port, din0(6) => data_addr_6_port, 
                           din0(5) => data_addr_5_port, din0(4) => 
                           data_addr_4_port, din0(3) => data_addr_3_port, 
                           din0(2) => data_addr_2_port, din0(1) => 
                           data_addr_1_port, din0(0) => data_addr_0_port, 
                           din1(31) => data_i_val(31), din1(30) => 
                           data_i_val(30), din1(29) => data_i_val(29), din1(28)
                           => data_i_val(28), din1(27) => data_i_val(27), 
                           din1(26) => data_i_val(26), din1(25) => 
                           data_i_val(25), din1(24) => data_i_val(24), din1(23)
                           => data_i_val(23), din1(22) => data_i_val(22), 
                           din1(21) => data_i_val(21), din1(20) => 
                           data_i_val(20), din1(19) => data_i_val(19), din1(18)
                           => data_i_val(18), din1(17) => data_i_val(17), 
                           din1(16) => data_i_val(16), din1(15) => 
                           data_i_val(15), din1(14) => data_i_val(14), din1(13)
                           => data_i_val(13), din1(12) => data_i_val(12), 
                           din1(11) => data_i_val(11), din1(10) => 
                           data_i_val(10), din1(9) => data_i_val(9), din1(8) =>
                           data_i_val(8), din1(7) => data_i_val(7), din1(6) => 
                           data_i_val(6), din1(5) => data_i_val(5), din1(4) => 
                           data_i_val(4), din1(3) => data_i_val(3), din1(2) => 
                           data_i_val(2), din1(1) => data_i_val(1), din1(0) => 
                           data_i_val(0), dout(31) => s4_result_31_port, 
                           dout(30) => s4_result_30_port, dout(29) => 
                           s4_result_29_port, dout(28) => s4_result_28_port, 
                           dout(27) => s4_result_27_port, dout(26) => 
                           s4_result_26_port, dout(25) => s4_result_25_port, 
                           dout(24) => s4_result_24_port, dout(23) => 
                           s4_result_23_port, dout(22) => s4_result_22_port, 
                           dout(21) => s4_result_21_port, dout(20) => 
                           s4_result_20_port, dout(19) => s4_result_19_port, 
                           dout(18) => s4_result_18_port, dout(17) => 
                           s4_result_17_port, dout(16) => s4_result_16_port, 
                           dout(15) => s4_result_15_port, dout(14) => 
                           s4_result_14_port, dout(13) => s4_result_13_port, 
                           dout(12) => s4_result_12_port, dout(11) => 
                           s4_result_11_port, dout(10) => s4_result_10_port, 
                           dout(9) => s4_result_9_port, dout(8) => 
                           s4_result_8_port, dout(7) => s4_result_7_port, 
                           dout(6) => s4_result_6_port, dout(5) => 
                           s4_result_5_port, dout(4) => s4_result_4_port, 
                           dout(3) => s4_result_3_port, dout(2) => 
                           s4_result_2_port, dout(1) => s4_result_1_port, 
                           dout(0) => s4_result_0_port);
   REG_RESULT : Reg_DATA_SIZE32_3 port map( rst => n111, en => cw(18), clk => 
                           clk, din(31) => s4_result_31_port, din(30) => 
                           s4_result_30_port, din(29) => s4_result_29_port, 
                           din(28) => s4_result_28_port, din(27) => 
                           s4_result_27_port, din(26) => s4_result_26_port, 
                           din(25) => s4_result_25_port, din(24) => 
                           s4_result_24_port, din(23) => s4_result_23_port, 
                           din(22) => s4_result_22_port, din(21) => 
                           s4_result_21_port, din(20) => s4_result_20_port, 
                           din(19) => s4_result_19_port, din(18) => 
                           s4_result_18_port, din(17) => s4_result_17_port, 
                           din(16) => s4_result_16_port, din(15) => 
                           s4_result_15_port, din(14) => s4_result_14_port, 
                           din(13) => s4_result_13_port, din(12) => 
                           s4_result_12_port, din(11) => s4_result_11_port, 
                           din(10) => s4_result_10_port, din(9) => 
                           s4_result_9_port, din(8) => s4_result_8_port, din(7)
                           => s4_result_7_port, din(6) => s4_result_6_port, 
                           din(5) => s4_result_5_port, din(4) => 
                           s4_result_4_port, din(3) => s4_result_3_port, din(2)
                           => s4_result_2_port, din(1) => s4_result_1_port, 
                           din(0) => s4_result_0_port, dout(31) => 
                           s5_result_31_port, dout(30) => s5_result_30_port, 
                           dout(29) => s5_result_29_port, dout(28) => 
                           s5_result_28_port, dout(27) => s5_result_27_port, 
                           dout(26) => s5_result_26_port, dout(25) => 
                           s5_result_25_port, dout(24) => s5_result_24_port, 
                           dout(23) => s5_result_23_port, dout(22) => 
                           s5_result_22_port, dout(21) => s5_result_21_port, 
                           dout(20) => s5_result_20_port, dout(19) => 
                           s5_result_19_port, dout(18) => s5_result_18_port, 
                           dout(17) => s5_result_17_port, dout(16) => 
                           s5_result_16_port, dout(15) => s5_result_15_port, 
                           dout(14) => s5_result_14_port, dout(13) => 
                           s5_result_13_port, dout(12) => s5_result_12_port, 
                           dout(11) => s5_result_11_port, dout(10) => 
                           s5_result_10_port, dout(9) => s5_result_9_port, 
                           dout(8) => s5_result_8_port, dout(7) => 
                           s5_result_7_port, dout(6) => s5_result_6_port, 
                           dout(5) => s5_result_5_port, dout(4) => 
                           s5_result_4_port, dout(3) => s5_result_3_port, 
                           dout(2) => s5_result_2_port, dout(1) => 
                           s5_result_1_port, dout(0) => s5_result_0_port);
   REG_WR4 : Reg_DATA_SIZE5_2 port map( rst => n110, en => cw(18), clk => clk, 
                           din(4) => s4_wr_addr_4_port, din(3) => 
                           s4_wr_addr_3_port, din(2) => s4_wr_addr_2_port, 
                           din(1) => s4_wr_addr_1_port, din(0) => 
                           s4_wr_addr_0_port, dout(4) => s5_wr_addr_4_port, 
                           dout(3) => s5_wr_addr_3_port, dout(2) => 
                           s5_wr_addr_2_port, dout(1) => s5_wr_addr_1_port, 
                           dout(0) => s5_wr_addr_0_port);
   REG_RESULT5 : Reg_DATA_SIZE32_2 port map( rst => n111, en => cw(19), clk => 
                           clk, din(31) => s5_result_31_port, din(30) => 
                           s5_result_30_port, din(29) => s5_result_29_port, 
                           din(28) => s5_result_28_port, din(27) => 
                           s5_result_27_port, din(26) => s5_result_26_port, 
                           din(25) => s5_result_25_port, din(24) => 
                           s5_result_24_port, din(23) => s5_result_23_port, 
                           din(22) => s5_result_22_port, din(21) => 
                           s5_result_21_port, din(20) => s5_result_20_port, 
                           din(19) => s5_result_19_port, din(18) => 
                           s5_result_18_port, din(17) => s5_result_17_port, 
                           din(16) => s5_result_16_port, din(15) => 
                           s5_result_15_port, din(14) => s5_result_14_port, 
                           din(13) => s5_result_13_port, din(12) => 
                           s5_result_12_port, din(11) => s5_result_11_port, 
                           din(10) => s5_result_10_port, din(9) => 
                           s5_result_9_port, din(8) => s5_result_8_port, din(7)
                           => s5_result_7_port, din(6) => s5_result_6_port, 
                           din(5) => s5_result_5_port, din(4) => 
                           s5_result_4_port, din(3) => s5_result_3_port, din(2)
                           => s5_result_2_port, din(1) => s5_result_1_port, 
                           din(0) => s5_result_0_port, dout(31) => 
                           s6_result_31_port, dout(30) => s6_result_30_port, 
                           dout(29) => s6_result_29_port, dout(28) => 
                           s6_result_28_port, dout(27) => s6_result_27_port, 
                           dout(26) => s6_result_26_port, dout(25) => 
                           s6_result_25_port, dout(24) => s6_result_24_port, 
                           dout(23) => s6_result_23_port, dout(22) => 
                           s6_result_22_port, dout(21) => s6_result_21_port, 
                           dout(20) => s6_result_20_port, dout(19) => 
                           s6_result_19_port, dout(18) => s6_result_18_port, 
                           dout(17) => s6_result_17_port, dout(16) => 
                           s6_result_16_port, dout(15) => s6_result_15_port, 
                           dout(14) => s6_result_14_port, dout(13) => 
                           s6_result_13_port, dout(12) => s6_result_12_port, 
                           dout(11) => s6_result_11_port, dout(10) => 
                           s6_result_10_port, dout(9) => s6_result_9_port, 
                           dout(8) => s6_result_8_port, dout(7) => 
                           s6_result_7_port, dout(6) => s6_result_6_port, 
                           dout(5) => s6_result_5_port, dout(4) => 
                           s6_result_4_port, dout(3) => s6_result_3_port, 
                           dout(2) => s6_result_2_port, dout(1) => 
                           s6_result_1_port, dout(0) => s6_result_0_port);
   REG_WR5 : Reg_DATA_SIZE5_1 port map( rst => n110, en => cw(19), clk => clk, 
                           din(4) => s5_wr_addr_4_port, din(3) => 
                           s5_wr_addr_3_port, din(2) => s5_wr_addr_2_port, 
                           din(1) => s5_wr_addr_1_port, din(0) => 
                           s5_wr_addr_0_port, dout(4) => s6_wr_addr_4_port, 
                           dout(3) => s6_wr_addr_3_port, dout(2) => 
                           s6_wr_addr_2_port, dout(1) => s6_wr_addr_1_port, 
                           dout(0) => s6_wr_addr_0_port);
   s4_reg_a_wait_reg : DFF_X1 port map( D => s3_reg_a_wait, CK => clk, Q => 
                           s4_reg_a_wait, QN => n97);
   s4_reg_b_wait_reg : DFF_X1 port map( D => s3_reg_b_wait, CK => clk, Q => 
                           s4_reg_b_wait, QN => n96);
   U3 : BUF_X1 port map( A => n103, Z => n108);
   U4 : AND3_X1 port map( A1 => istr_val(29), A2 => istr_val(27), A3 => 
                           istr_val(28), ZN => n72);
   U5 : INV_X1 port map( A => istr_val(30), ZN => n47);
   U6 : CLKBUF_X1 port map( A => s2_jpc_28_port, Z => n52);
   U7 : CLKBUF_X1 port map( A => s3_exe_out_30_port, Z => n80);
   U8 : AND2_X1 port map( A1 => s2_imm_l_ext_1_port, A2 => n103, ZN => 
                           s2_imm_i_ext_1_port);
   U9 : CLKBUF_X1 port map( A => s3_exe_out_29_port, Z => n81);
   U10 : CLKBUF_X1 port map( A => s3_exe_out_28_port, Z => n82);
   U11 : CLKBUF_X1 port map( A => s3_exe_out_31_port, Z => n83);
   U12 : CLKBUF_X1 port map( A => n121, Z => istr_addr_2_port);
   U13 : CLKBUF_X1 port map( A => n120, Z => istr_addr_28_port);
   U14 : AND2_X2 port map( A1 => calu(3), A2 => n109, ZN => n95);
   U15 : BUF_X1 port map( A => istr_val(28), Z => n86);
   U16 : CLKBUF_X1 port map( A => s3_b_sel_0_port, Z => n87);
   U17 : INV_X1 port map( A => istr_val(30), ZN => n88);
   U18 : AND3_X1 port map( A1 => istr_val(29), A2 => istr_val(27), A3 => n86, 
                           ZN => n89);
   U19 : CLKBUF_X1 port map( A => n87, Z => n90);
   U20 : INV_X1 port map( A => sig_div_port, ZN => n91);
   U21 : CLKBUF_X1 port map( A => n104, Z => sig_sqrt_port);
   U22 : CLKBUF_X1 port map( A => calu(1), Z => n93);
   U23 : CLKBUF_X1 port map( A => n122, Z => istr_addr_1_port);
   U24 : NOR2_X1 port map( A1 => n117, A2 => n116, ZN => s3_mul_sign);
   U25 : INV_X1 port map( A => n49, ZN => n76);
   U26 : NAND2_X1 port map( A1 => s2_imm_l_ext_31_port, A2 => n98, ZN => n55);
   U27 : INV_X1 port map( A => istr_val(4), ZN => n66);
   U28 : INV_X1 port map( A => istr_val(8), ZN => n62);
   U29 : INV_X1 port map( A => istr_val(9), ZN => n61);
   U30 : INV_X1 port map( A => istr_val(10), ZN => n60);
   U31 : INV_X1 port map( A => istr_val(13), ZN => n57);
   U32 : INV_X1 port map( A => istr_val(11), ZN => n59);
   U33 : INV_X1 port map( A => istr_val(2), ZN => n68);
   U34 : INV_X1 port map( A => istr_val(0), ZN => n70);
   U35 : INV_X1 port map( A => istr_val(3), ZN => n67);
   U36 : OAI21_X1 port map( B1 => n98, B2 => n63, A => n55, ZN => 
                           s2_imm_i_ext_23_port);
   U37 : INV_X1 port map( A => istr_val(7), ZN => n63);
   U38 : OAI21_X1 port map( B1 => n98, B2 => n65, A => n55, ZN => 
                           s2_imm_i_ext_21_port);
   U39 : INV_X1 port map( A => istr_val(5), ZN => n65);
   U40 : OAI21_X1 port map( B1 => n98, B2 => n64, A => n55, ZN => 
                           s2_imm_i_ext_22_port);
   U41 : INV_X1 port map( A => istr_val(6), ZN => n64);
   U42 : OAI21_X1 port map( B1 => n98, B2 => n58, A => n55, ZN => 
                           s2_imm_i_ext_28_port);
   U43 : INV_X1 port map( A => istr_val(12), ZN => n58);
   U44 : OAI21_X1 port map( B1 => n98, B2 => n69, A => n55, ZN => 
                           s2_imm_i_ext_17_port);
   U45 : INV_X1 port map( A => istr_val(1), ZN => n69);
   U46 : INV_X1 port map( A => istr_val(27), ZN => n50);
   U47 : AND2_X1 port map( A1 => s2_imm_l_ext_7_port, A2 => n98, ZN => 
                           s2_imm_i_ext_7_port);
   U48 : INV_X1 port map( A => istr_val(31), ZN => n71);
   U49 : BUF_X2 port map( A => rst, Z => n111);
   U50 : INV_X1 port map( A => istr_val(14), ZN => n56);
   U51 : NOR2_X1 port map( A1 => istr_val(29), A2 => istr_val(31), ZN => n49);
   U52 : OAI21_X1 port map( B1 => n99, B2 => n54, A => n55, ZN => 
                           s2_imm_i_ext_31_port);
   U53 : INV_X1 port map( A => istr_val(15), ZN => n54);
   U54 : BUF_X2 port map( A => rst, Z => n110);
   U55 : OAI21_X1 port map( B1 => cw(6), B2 => n53, A => n78, ZN => n48);
   U56 : OAI21_X1 port map( B1 => ir_out_28_port, B2 => n50, A => n75, ZN => 
                           n79);
   U57 : OR2_X1 port map( A1 => s6_en_wb, A2 => cw(19), ZN => n45);
   U58 : NOR3_X1 port map( A1 => n77, A2 => n76, A3 => n75, ZN => s2_a_f_b_en);
   U59 : OR2_X1 port map( A1 => s3_reg_a_wait, A2 => s3_reg_b_wait, ZN => 
                           sig_ral_port);
   U60 : NOR2_X1 port map( A1 => cw(7), A2 => n46, ZN => s3_b_sel_f_en);
   U61 : INV_X1 port map( A => n46, ZN => s3_a_sel_f_en);
   U62 : NOR2_X1 port map( A1 => n74, A2 => n77, ZN => s2_a_f_j_en);
   U63 : NAND2_X1 port map( A1 => cw(17), A2 => n53, ZN => n46);
   U64 : NAND2_X1 port map( A1 => cw(19), A2 => n53, ZN => n43);
   U65 : NOR2_X1 port map( A1 => cw(7), A2 => n43, ZN => s3_b_sel_ff_en);
   U66 : INV_X1 port map( A => n43, ZN => s3_a_sel_ff_en);
   U67 : NOR2_X1 port map( A1 => n73, A2 => n74, ZN => s2_a_ff_j_en);
   U68 : NOR3_X1 port map( A1 => n75, A2 => n73, A3 => n76, ZN => s2_a_ff_b_en)
                           ;
   U69 : OR2_X1 port map( A1 => cw(19), A2 => cw(6), ZN => s2_rf_en);
   U70 : INV_X1 port map( A => cw(17), ZN => n73);
   U71 : INV_X1 port map( A => cw(9), ZN => n77);
   U72 : CLKBUF_X1 port map( A => n108, Z => n99);
   U73 : BUF_X4 port map( A => n108, Z => n98);
   U74 : NAND4_X1 port map( A1 => n49, A2 => n50, A3 => n51, A4 => n88, ZN => 
                           s2_wr_addr_sel);
   U75 : INV_X1 port map( A => n50, ZN => ir_out_27_port);
   U76 : NAND4_X1 port map( A1 => istr_val(30), A2 => ir_out_27_port, A3 => n49
                           , A4 => n51, ZN => n74);
   U77 : INV_X1 port map( A => n51, ZN => ir_out_28_port);
   U78 : INV_X1 port map( A => n86, ZN => n51);
   U79 : NAND4_X1 port map( A1 => n72, A2 => n71, A3 => istr_val(26), A4 => n47
                           , ZN => n102);
   U80 : NAND4_X1 port map( A1 => n89, A2 => n71, A3 => istr_val(26), A4 => n88
                           , ZN => n103);
   U81 : OAI21_X1 port map( B1 => n98, B2 => n56, A => n55, ZN => 
                           s2_imm_i_ext_30_port);
   U82 : OAI21_X1 port map( B1 => n98, B2 => n60, A => n55, ZN => 
                           s2_imm_i_ext_26_port);
   U83 : INV_X1 port map( A => sig_sqrt_port, ZN => n113);
   U84 : AND3_X2 port map( A1 => calu(2), A2 => n95, A3 => n112, ZN => n104);
   U85 : CLKBUF_X1 port map( A => s3_exe_out_0_port, Z => n105);
   U86 : OAI21_X1 port map( B1 => n98, B2 => n57, A => n55, ZN => 
                           s2_imm_i_ext_29_port);
   U87 : OAI21_X1 port map( B1 => n98, B2 => n59, A => n55, ZN => 
                           s2_imm_i_ext_27_port);
   U88 : OAI21_X1 port map( B1 => n98, B2 => n61, A => n55, ZN => 
                           s2_imm_i_ext_25_port);
   U89 : OAI21_X1 port map( B1 => n98, B2 => n62, A => n55, ZN => 
                           s2_imm_i_ext_24_port);
   U90 : AND2_X1 port map( A1 => s2_imm_l_ext_8_port, A2 => n98, ZN => 
                           s2_imm_i_ext_8_port);
   U91 : NAND2_X1 port map( A1 => n113, A2 => n91, ZN => s3_exe_sel_1_port);
   U92 : NOR2_X1 port map( A1 => n118, A2 => n116, ZN => s3_div_sign);
   U93 : AND2_X1 port map( A1 => s2_imm_l_ext_9_port, A2 => n98, ZN => 
                           s2_imm_i_ext_9_port);
   U96 : AND2_X1 port map( A1 => s2_imm_l_ext_6_port, A2 => n98, ZN => 
                           s2_imm_i_ext_6_port);
   U97 : AND2_X1 port map( A1 => s2_imm_l_ext_5_port, A2 => n98, ZN => 
                           s2_imm_i_ext_5_port);
   U98 : AND2_X1 port map( A1 => s2_imm_l_ext_4_port, A2 => n98, ZN => 
                           s2_imm_i_ext_4_port);
   U99 : AND2_X1 port map( A1 => s2_imm_l_ext_3_port, A2 => n99, ZN => 
                           s2_imm_i_ext_3_port);
   U100 : AND2_X1 port map( A1 => s2_imm_l_ext_2_port, A2 => n108, ZN => 
                           s2_imm_i_ext_2_port);
   U101 : AND2_X1 port map( A1 => n102, A2 => s2_imm_l_ext_0_port, ZN => 
                           s2_imm_i_ext_0_port);
   U102 : OAI21_X1 port map( B1 => n98, B2 => n66, A => n55, ZN => 
                           s2_imm_i_ext_20_port);
   U103 : OAI21_X1 port map( B1 => n98, B2 => n67, A => n55, ZN => 
                           s2_imm_i_ext_19_port);
   U104 : AND2_X1 port map( A1 => s2_imm_l_ext_15_port, A2 => n98, ZN => 
                           s2_imm_i_ext_15_port);
   U105 : OAI21_X1 port map( B1 => n98, B2 => n68, A => n55, ZN => 
                           s2_imm_i_ext_18_port);
   U106 : OAI21_X1 port map( B1 => n98, B2 => n70, A => n55, ZN => 
                           s2_imm_i_ext_16_port);
   U107 : AND2_X1 port map( A1 => s2_imm_l_ext_14_port, A2 => n98, ZN => 
                           s2_imm_i_ext_14_port);
   U108 : AND2_X1 port map( A1 => s2_imm_l_ext_13_port, A2 => n98, ZN => 
                           s2_imm_i_ext_13_port);
   U109 : AND2_X1 port map( A1 => s2_imm_l_ext_11_port, A2 => n98, ZN => 
                           s2_imm_i_ext_11_port);
   U110 : AND2_X1 port map( A1 => s2_imm_l_ext_12_port, A2 => n98, ZN => 
                           s2_imm_i_ext_12_port);
   U111 : AND2_X1 port map( A1 => s2_imm_l_ext_10_port, A2 => n98, ZN => 
                           s2_imm_i_ext_10_port);
   U112 : CLKBUF_X1 port map( A => n123, Z => istr_addr_0_port);
   U113 : CLKBUF_X1 port map( A => cw(1), Z => n107);
   U114 : INV_X1 port map( A => calu(4), ZN => n109);
   U115 : NOR2_X1 port map( A1 => calu(1), A2 => calu(0), ZN => n112);
   U116 : INV_X1 port map( A => calu(2), ZN => n114);
   U117 : NAND3_X1 port map( A1 => n114, A2 => n95, A3 => calu(1), ZN => n118);
   U118 : INV_X1 port map( A => calu(0), ZN => n116);
   U119 : INV_X1 port map( A => calu(1), ZN => n115);
   U120 : NAND3_X1 port map( A1 => n115, A2 => n95, A3 => n114, ZN => n117);
   U121 : INV_X1 port map( A => n117, ZN => sig_mul_port);
   U122 : INV_X1 port map( A => n118, ZN => sig_div_port);

end SYN_data_path_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity 
   ControlUnit_ISTR_SIZE32_DATA_SIZE32_OPCD_SIZE6_FUNC_SIZE11_CWRD_SIZE20_CALU_SIZE5_ADDR_SIZE32 
   is

   port( clk, rst : in std_logic;  ir, pc, reg_a, ld_a : in std_logic_vector 
         (31 downto 0);  sig_bal : in std_logic;  sig_bpw : out std_logic;  
         sig_jral, sig_ral, sig_mul, sig_div, sig_sqrt : in std_logic;  cw : 
         out std_logic_vector (19 downto 0);  calu : out std_logic_vector (4 
         downto 0));

end 
   ControlUnit_ISTR_SIZE32_DATA_SIZE32_OPCD_SIZE6_FUNC_SIZE11_CWRD_SIZE20_CALU_SIZE5_ADDR_SIZE32;

architecture SYN_control_unit_arch of 
   ControlUnit_ISTR_SIZE32_DATA_SIZE32_OPCD_SIZE6_FUNC_SIZE11_CWRD_SIZE20_CALU_SIZE5_ADDR_SIZE32 
   is

   component Branch_DATA_SIZE32_OPCD_SIZE6_ADDR_SIZE32
      port( rst, clk : in std_logic;  reg_a, ld_a : in std_logic_vector (31 
            downto 0);  opcd : in std_logic_vector (5 downto 0);  addr : in 
            std_logic_vector (31 downto 0);  sig_bal : in std_logic;  sig_bpw, 
            sig_brt : out std_logic);
   end component;
   
   component StallGenerator_CWRD_SIZE20
      port( rst, clk, sig_ral, sig_bpw, sig_jral, sig_mul, sig_div, sig_sqrt : 
            in std_logic;  stall_flag : out std_logic_vector (4 downto 0));
   end component;
   
   component 
      CwGenerator_DATA_SIZE32_OPCD_SIZE6_FUNC_SIZE11_CWRD_SIZE20_CALU_SIZE5
      port( clk, rst : in std_logic;  opcd : in std_logic_vector (5 downto 0); 
            func : in std_logic_vector (10 downto 0);  stall_flag : in 
            std_logic_vector (4 downto 0);  taken : in std_logic;  cw : out 
            std_logic_vector (19 downto 0);  calu : out std_logic_vector (4 
            downto 0));
   end component;
   
   signal sig_bpw_port, stall_flag_4_port, stall_flag_3_port, stall_flag_2_port
      , stall_flag_1_port, stall_flag_0_port, sig_brt, net163693, net163694, 
      net163695, net163696, net163697, net163698, net163699, net163700, 
      net163701, net163702, net163703, net163704, net163705, net163706, 
      net163707, net163708, net163709, net163710 : std_logic;

begin
   sig_bpw <= sig_bpw_port;
   
   cw(2) <= '0';
   cw(3) <= '0';
   cw(4) <= '0';
   cw(5) <= '0';
   cw(6) <= '0';
   cw(7) <= '0';
   cw(8) <= '0';
   cw(9) <= '0';
   cw(10) <= '0';
   cw(11) <= '0';
   cw(12) <= '0';
   cw(13) <= '0';
   cw(14) <= '0';
   cw(15) <= '0';
   cw(16) <= '0';
   cw(17) <= '0';
   cw(18) <= '0';
   cw(19) <= '0';
   CW_GEN : 
                           CwGenerator_DATA_SIZE32_OPCD_SIZE6_FUNC_SIZE11_CWRD_SIZE20_CALU_SIZE5 
                           port map( clk => clk, rst => rst, opcd(5) => ir(31),
                           opcd(4) => ir(30), opcd(3) => ir(29), opcd(2) => 
                           ir(28), opcd(1) => ir(27), opcd(0) => ir(26), 
                           func(10) => ir(10), func(9) => ir(9), func(8) => 
                           ir(8), func(7) => ir(7), func(6) => ir(6), func(5) 
                           => ir(5), func(4) => ir(4), func(3) => ir(3), 
                           func(2) => ir(2), func(1) => ir(1), func(0) => ir(0)
                           , stall_flag(4) => stall_flag_4_port, stall_flag(3) 
                           => stall_flag_3_port, stall_flag(2) => 
                           stall_flag_2_port, stall_flag(1) => 
                           stall_flag_1_port, stall_flag(0) => 
                           stall_flag_0_port, taken => sig_brt, cw(19) => 
                           net163693, cw(18) => net163694, cw(17) => net163695,
                           cw(16) => net163696, cw(15) => net163697, cw(14) => 
                           net163698, cw(13) => net163699, cw(12) => net163700,
                           cw(11) => net163701, cw(10) => net163702, cw(9) => 
                           net163703, cw(8) => net163704, cw(7) => net163705, 
                           cw(6) => net163706, cw(5) => net163707, cw(4) => 
                           net163708, cw(3) => net163709, cw(2) => net163710, 
                           cw(1) => cw(1), cw(0) => cw(0), calu(4) => calu(4), 
                           calu(3) => calu(3), calu(2) => calu(2), calu(1) => 
                           calu(1), calu(0) => calu(0));
   S_GEN : StallGenerator_CWRD_SIZE20 port map( rst => rst, clk => clk, sig_ral
                           => sig_ral, sig_bpw => sig_bpw_port, sig_jral => 
                           sig_jral, sig_mul => sig_mul, sig_div => sig_div, 
                           sig_sqrt => sig_sqrt, stall_flag(4) => 
                           stall_flag_4_port, stall_flag(3) => 
                           stall_flag_3_port, stall_flag(2) => 
                           stall_flag_2_port, stall_flag(1) => 
                           stall_flag_1_port, stall_flag(0) => 
                           stall_flag_0_port);
   BR : Branch_DATA_SIZE32_OPCD_SIZE6_ADDR_SIZE32 port map( rst => rst, clk => 
                           clk, reg_a(31) => reg_a(31), reg_a(30) => reg_a(30),
                           reg_a(29) => reg_a(29), reg_a(28) => reg_a(28), 
                           reg_a(27) => reg_a(27), reg_a(26) => reg_a(26), 
                           reg_a(25) => reg_a(25), reg_a(24) => reg_a(24), 
                           reg_a(23) => reg_a(23), reg_a(22) => reg_a(22), 
                           reg_a(21) => reg_a(21), reg_a(20) => reg_a(20), 
                           reg_a(19) => reg_a(19), reg_a(18) => reg_a(18), 
                           reg_a(17) => reg_a(17), reg_a(16) => reg_a(16), 
                           reg_a(15) => reg_a(15), reg_a(14) => reg_a(14), 
                           reg_a(13) => reg_a(13), reg_a(12) => reg_a(12), 
                           reg_a(11) => reg_a(11), reg_a(10) => reg_a(10), 
                           reg_a(9) => reg_a(9), reg_a(8) => reg_a(8), reg_a(7)
                           => reg_a(7), reg_a(6) => reg_a(6), reg_a(5) => 
                           reg_a(5), reg_a(4) => reg_a(4), reg_a(3) => reg_a(3)
                           , reg_a(2) => reg_a(2), reg_a(1) => reg_a(1), 
                           reg_a(0) => reg_a(0), ld_a(31) => ld_a(31), ld_a(30)
                           => ld_a(30), ld_a(29) => ld_a(29), ld_a(28) => 
                           ld_a(28), ld_a(27) => ld_a(27), ld_a(26) => ld_a(26)
                           , ld_a(25) => ld_a(25), ld_a(24) => ld_a(24), 
                           ld_a(23) => ld_a(23), ld_a(22) => ld_a(22), ld_a(21)
                           => ld_a(21), ld_a(20) => ld_a(20), ld_a(19) => 
                           ld_a(19), ld_a(18) => ld_a(18), ld_a(17) => ld_a(17)
                           , ld_a(16) => ld_a(16), ld_a(15) => ld_a(15), 
                           ld_a(14) => ld_a(14), ld_a(13) => ld_a(13), ld_a(12)
                           => ld_a(12), ld_a(11) => ld_a(11), ld_a(10) => 
                           ld_a(10), ld_a(9) => ld_a(9), ld_a(8) => ld_a(8), 
                           ld_a(7) => ld_a(7), ld_a(6) => ld_a(6), ld_a(5) => 
                           ld_a(5), ld_a(4) => ld_a(4), ld_a(3) => ld_a(3), 
                           ld_a(2) => ld_a(2), ld_a(1) => ld_a(1), ld_a(0) => 
                           ld_a(0), opcd(5) => ir(31), opcd(4) => ir(30), 
                           opcd(3) => ir(29), opcd(2) => ir(28), opcd(1) => 
                           ir(27), opcd(0) => ir(26), addr(31) => pc(31), 
                           addr(30) => pc(30), addr(29) => pc(29), addr(28) => 
                           pc(28), addr(27) => pc(27), addr(26) => pc(26), 
                           addr(25) => pc(25), addr(24) => pc(24), addr(23) => 
                           pc(23), addr(22) => pc(22), addr(21) => pc(21), 
                           addr(20) => pc(20), addr(19) => pc(19), addr(18) => 
                           pc(18), addr(17) => pc(17), addr(16) => pc(16), 
                           addr(15) => pc(15), addr(14) => pc(14), addr(13) => 
                           pc(13), addr(12) => pc(12), addr(11) => pc(11), 
                           addr(10) => pc(10), addr(9) => pc(9), addr(8) => 
                           pc(8), addr(7) => pc(7), addr(6) => pc(6), addr(5) 
                           => pc(5), addr(4) => pc(4), addr(3) => pc(3), 
                           addr(2) => pc(2), addr(1) => pc(1), addr(0) => pc(0)
                           , sig_bal => sig_bal, sig_bpw => sig_bpw_port, 
                           sig_brt => sig_brt);

end SYN_control_unit_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4 is

   port( clk, rst : in std_logic;  en_iram : out std_logic;  pc_bus : out 
         std_logic_vector (31 downto 0);  ir_bus : in std_logic_vector (31 
         downto 0);  en_dram : out std_logic;  addr_bus, di_bus : out 
         std_logic_vector (31 downto 0);  do_bus : in std_logic_vector (31 
         downto 0);  dr_cw : out std_logic_vector (3 downto 0));

end Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4;

architecture SYN_dlx_arch of Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4
   is

   component 
      DataPath_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_OPCD_SIZE6_IMME_SIZE16_CWRD_SIZE20_CALU_SIZE5_DRCW_SIZE4
      port( clk, rst : in std_logic;  istr_addr : out std_logic_vector (31 
            downto 0);  istr_val : in std_logic_vector (31 downto 0);  ir_out, 
            pc_out, reg_a_out, ld_a_out, data_addr : out std_logic_vector (31 
            downto 0);  data_i_val : in std_logic_vector (31 downto 0);  
            data_o_val : out std_logic_vector (31 downto 0);  cw : in 
            std_logic_vector (19 downto 0);  dr_cw : out std_logic_vector (3 
            downto 0);  calu : in std_logic_vector (4 downto 0);  sig_bal : out
            std_logic;  sig_bpw : in std_logic;  sig_jral, sig_ral, sig_mul, 
            sig_div, sig_sqrt : out std_logic);
   end component;
   
   component 
      ControlUnit_ISTR_SIZE32_DATA_SIZE32_OPCD_SIZE6_FUNC_SIZE11_CWRD_SIZE20_CALU_SIZE5_ADDR_SIZE32
      port( clk, rst : in std_logic;  ir, pc, reg_a, ld_a : in std_logic_vector
            (31 downto 0);  sig_bal : in std_logic;  sig_bpw : out std_logic;  
            sig_jral, sig_ral, sig_mul, sig_div, sig_sqrt : in std_logic;  cw :
            out std_logic_vector (19 downto 0);  calu : out std_logic_vector (4
            downto 0));
   end component;
   
   signal en_iram_port, ir_31_port, ir_30_port, ir_29_port, ir_28_port, 
      ir_27_port, ir_26_port, ir_25_port, ir_24_port, ir_23_port, ir_22_port, 
      ir_21_port, ir_20_port, ir_19_port, ir_18_port, ir_17_port, ir_16_port, 
      ir_15_port, ir_14_port, ir_13_port, ir_12_port, ir_11_port, ir_10_port, 
      ir_9_port, ir_8_port, ir_7_port, ir_6_port, ir_5_port, ir_4_port, 
      ir_3_port, ir_2_port, ir_1_port, ir_0_port, pc_31_port, pc_30_port, 
      pc_29_port, pc_28_port, pc_27_port, pc_26_port, pc_25_port, pc_24_port, 
      pc_23_port, pc_22_port, pc_21_port, pc_20_port, pc_19_port, pc_18_port, 
      pc_17_port, pc_16_port, pc_15_port, pc_14_port, pc_13_port, pc_12_port, 
      pc_11_port, pc_10_port, pc_9_port, pc_8_port, pc_7_port, pc_6_port, 
      pc_5_port, pc_4_port, pc_3_port, pc_2_port, pc_1_port, pc_0_port, 
      reg_a_val_31_port, reg_a_val_30_port, reg_a_val_29_port, 
      reg_a_val_28_port, reg_a_val_27_port, reg_a_val_26_port, 
      reg_a_val_25_port, reg_a_val_24_port, reg_a_val_23_port, 
      reg_a_val_22_port, reg_a_val_21_port, reg_a_val_20_port, 
      reg_a_val_19_port, reg_a_val_18_port, reg_a_val_17_port, 
      reg_a_val_16_port, reg_a_val_15_port, reg_a_val_14_port, 
      reg_a_val_13_port, reg_a_val_12_port, reg_a_val_11_port, 
      reg_a_val_10_port, reg_a_val_9_port, reg_a_val_8_port, reg_a_val_7_port, 
      reg_a_val_6_port, reg_a_val_5_port, reg_a_val_4_port, reg_a_val_3_port, 
      reg_a_val_2_port, reg_a_val_1_port, reg_a_val_0_port, ld_a_val_31_port, 
      ld_a_val_30_port, ld_a_val_29_port, ld_a_val_28_port, ld_a_val_27_port, 
      ld_a_val_26_port, ld_a_val_25_port, ld_a_val_24_port, ld_a_val_23_port, 
      ld_a_val_22_port, ld_a_val_21_port, ld_a_val_20_port, ld_a_val_19_port, 
      ld_a_val_18_port, ld_a_val_17_port, ld_a_val_16_port, ld_a_val_15_port, 
      ld_a_val_14_port, ld_a_val_13_port, ld_a_val_12_port, ld_a_val_11_port, 
      ld_a_val_10_port, ld_a_val_9_port, ld_a_val_8_port, ld_a_val_7_port, 
      ld_a_val_6_port, ld_a_val_5_port, ld_a_val_4_port, ld_a_val_3_port, 
      ld_a_val_2_port, ld_a_val_1_port, ld_a_val_0_port, sig_bal, sig_bpw, 
      sig_jral, sig_ral, sig_mul, sig_div, sig_sqrt, cw_19_port, cw_18_port, 
      cw_17_port, cw_16_port, cw_15_port, cw_14_port, cw_13_port, cw_12_port, 
      cw_11_port, cw_10_port, cw_9_port, cw_8_port, cw_7_port, cw_6_port, 
      cw_5_port, cw_4_port, cw_3_port, cw_2_port, cw_1_port, calu_4_port, 
      calu_3_port, calu_2_port, calu_1_port, calu_0_port, net163675, net163676,
      net163677, net163678, net163679, net163680, net163681, net163682, 
      net163683, net163684, net163685, net163686, net163687, net163688, 
      net163689, net163690, net163691, net163692 : std_logic;

begin
   en_iram <= en_iram_port;
   
   en_dram <= '1';
   cw_2_port <= '0';
   cw_3_port <= '0';
   cw_4_port <= '0';
   cw_5_port <= '0';
   cw_6_port <= '0';
   cw_7_port <= '0';
   cw_8_port <= '0';
   cw_9_port <= '0';
   cw_10_port <= '0';
   cw_11_port <= '0';
   cw_12_port <= '0';
   cw_13_port <= '0';
   cw_14_port <= '0';
   cw_15_port <= '0';
   cw_16_port <= '0';
   cw_17_port <= '0';
   cw_18_port <= '0';
   cw_19_port <= '0';
   CU0 : 
                           ControlUnit_ISTR_SIZE32_DATA_SIZE32_OPCD_SIZE6_FUNC_SIZE11_CWRD_SIZE20_CALU_SIZE5_ADDR_SIZE32 
                           port map( clk => clk, rst => rst, ir(31) => 
                           ir_31_port, ir(30) => ir_30_port, ir(29) => 
                           ir_29_port, ir(28) => ir_28_port, ir(27) => 
                           ir_27_port, ir(26) => ir_26_port, ir(25) => 
                           ir_25_port, ir(24) => ir_24_port, ir(23) => 
                           ir_23_port, ir(22) => ir_22_port, ir(21) => 
                           ir_21_port, ir(20) => ir_20_port, ir(19) => 
                           ir_19_port, ir(18) => ir_18_port, ir(17) => 
                           ir_17_port, ir(16) => ir_16_port, ir(15) => 
                           ir_15_port, ir(14) => ir_14_port, ir(13) => 
                           ir_13_port, ir(12) => ir_12_port, ir(11) => 
                           ir_11_port, ir(10) => ir_10_port, ir(9) => ir_9_port
                           , ir(8) => ir_8_port, ir(7) => ir_7_port, ir(6) => 
                           ir_6_port, ir(5) => ir_5_port, ir(4) => ir_4_port, 
                           ir(3) => ir_3_port, ir(2) => ir_2_port, ir(1) => 
                           ir_1_port, ir(0) => ir_0_port, pc(31) => pc_31_port,
                           pc(30) => pc_30_port, pc(29) => pc_29_port, pc(28) 
                           => pc_28_port, pc(27) => pc_27_port, pc(26) => 
                           pc_26_port, pc(25) => pc_25_port, pc(24) => 
                           pc_24_port, pc(23) => pc_23_port, pc(22) => 
                           pc_22_port, pc(21) => pc_21_port, pc(20) => 
                           pc_20_port, pc(19) => pc_19_port, pc(18) => 
                           pc_18_port, pc(17) => pc_17_port, pc(16) => 
                           pc_16_port, pc(15) => pc_15_port, pc(14) => 
                           pc_14_port, pc(13) => pc_13_port, pc(12) => 
                           pc_12_port, pc(11) => pc_11_port, pc(10) => 
                           pc_10_port, pc(9) => pc_9_port, pc(8) => pc_8_port, 
                           pc(7) => pc_7_port, pc(6) => pc_6_port, pc(5) => 
                           pc_5_port, pc(4) => pc_4_port, pc(3) => pc_3_port, 
                           pc(2) => pc_2_port, pc(1) => pc_1_port, pc(0) => 
                           pc_0_port, reg_a(31) => reg_a_val_31_port, reg_a(30)
                           => reg_a_val_30_port, reg_a(29) => reg_a_val_29_port
                           , reg_a(28) => reg_a_val_28_port, reg_a(27) => 
                           reg_a_val_27_port, reg_a(26) => reg_a_val_26_port, 
                           reg_a(25) => reg_a_val_25_port, reg_a(24) => 
                           reg_a_val_24_port, reg_a(23) => reg_a_val_23_port, 
                           reg_a(22) => reg_a_val_22_port, reg_a(21) => 
                           reg_a_val_21_port, reg_a(20) => reg_a_val_20_port, 
                           reg_a(19) => reg_a_val_19_port, reg_a(18) => 
                           reg_a_val_18_port, reg_a(17) => reg_a_val_17_port, 
                           reg_a(16) => reg_a_val_16_port, reg_a(15) => 
                           reg_a_val_15_port, reg_a(14) => reg_a_val_14_port, 
                           reg_a(13) => reg_a_val_13_port, reg_a(12) => 
                           reg_a_val_12_port, reg_a(11) => reg_a_val_11_port, 
                           reg_a(10) => reg_a_val_10_port, reg_a(9) => 
                           reg_a_val_9_port, reg_a(8) => reg_a_val_8_port, 
                           reg_a(7) => reg_a_val_7_port, reg_a(6) => 
                           reg_a_val_6_port, reg_a(5) => reg_a_val_5_port, 
                           reg_a(4) => reg_a_val_4_port, reg_a(3) => 
                           reg_a_val_3_port, reg_a(2) => reg_a_val_2_port, 
                           reg_a(1) => reg_a_val_1_port, reg_a(0) => 
                           reg_a_val_0_port, ld_a(31) => ld_a_val_31_port, 
                           ld_a(30) => ld_a_val_30_port, ld_a(29) => 
                           ld_a_val_29_port, ld_a(28) => ld_a_val_28_port, 
                           ld_a(27) => ld_a_val_27_port, ld_a(26) => 
                           ld_a_val_26_port, ld_a(25) => ld_a_val_25_port, 
                           ld_a(24) => ld_a_val_24_port, ld_a(23) => 
                           ld_a_val_23_port, ld_a(22) => ld_a_val_22_port, 
                           ld_a(21) => ld_a_val_21_port, ld_a(20) => 
                           ld_a_val_20_port, ld_a(19) => ld_a_val_19_port, 
                           ld_a(18) => ld_a_val_18_port, ld_a(17) => 
                           ld_a_val_17_port, ld_a(16) => ld_a_val_16_port, 
                           ld_a(15) => ld_a_val_15_port, ld_a(14) => 
                           ld_a_val_14_port, ld_a(13) => ld_a_val_13_port, 
                           ld_a(12) => ld_a_val_12_port, ld_a(11) => 
                           ld_a_val_11_port, ld_a(10) => ld_a_val_10_port, 
                           ld_a(9) => ld_a_val_9_port, ld_a(8) => 
                           ld_a_val_8_port, ld_a(7) => ld_a_val_7_port, ld_a(6)
                           => ld_a_val_6_port, ld_a(5) => ld_a_val_5_port, 
                           ld_a(4) => ld_a_val_4_port, ld_a(3) => 
                           ld_a_val_3_port, ld_a(2) => ld_a_val_2_port, ld_a(1)
                           => ld_a_val_1_port, ld_a(0) => ld_a_val_0_port, 
                           sig_bal => sig_bal, sig_bpw => sig_bpw, sig_jral => 
                           sig_jral, sig_ral => sig_ral, sig_mul => sig_mul, 
                           sig_div => sig_div, sig_sqrt => sig_sqrt, cw(19) => 
                           net163675, cw(18) => net163676, cw(17) => net163677,
                           cw(16) => net163678, cw(15) => net163679, cw(14) => 
                           net163680, cw(13) => net163681, cw(12) => net163682,
                           cw(11) => net163683, cw(10) => net163684, cw(9) => 
                           net163685, cw(8) => net163686, cw(7) => net163687, 
                           cw(6) => net163688, cw(5) => net163689, cw(4) => 
                           net163690, cw(3) => net163691, cw(2) => net163692, 
                           cw(1) => cw_1_port, cw(0) => en_iram_port, calu(4) 
                           => calu_4_port, calu(3) => calu_3_port, calu(2) => 
                           calu_2_port, calu(1) => calu_1_port, calu(0) => 
                           calu_0_port);
   DP0 : 
                           DataPath_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_OPCD_SIZE6_IMME_SIZE16_CWRD_SIZE20_CALU_SIZE5_DRCW_SIZE4 
                           port map( clk => clk, rst => rst, istr_addr(31) => 
                           pc_bus(31), istr_addr(30) => pc_bus(30), 
                           istr_addr(29) => pc_bus(29), istr_addr(28) => 
                           pc_bus(28), istr_addr(27) => pc_bus(27), 
                           istr_addr(26) => pc_bus(26), istr_addr(25) => 
                           pc_bus(25), istr_addr(24) => pc_bus(24), 
                           istr_addr(23) => pc_bus(23), istr_addr(22) => 
                           pc_bus(22), istr_addr(21) => pc_bus(21), 
                           istr_addr(20) => pc_bus(20), istr_addr(19) => 
                           pc_bus(19), istr_addr(18) => pc_bus(18), 
                           istr_addr(17) => pc_bus(17), istr_addr(16) => 
                           pc_bus(16), istr_addr(15) => pc_bus(15), 
                           istr_addr(14) => pc_bus(14), istr_addr(13) => 
                           pc_bus(13), istr_addr(12) => pc_bus(12), 
                           istr_addr(11) => pc_bus(11), istr_addr(10) => 
                           pc_bus(10), istr_addr(9) => pc_bus(9), istr_addr(8) 
                           => pc_bus(8), istr_addr(7) => pc_bus(7), 
                           istr_addr(6) => pc_bus(6), istr_addr(5) => pc_bus(5)
                           , istr_addr(4) => pc_bus(4), istr_addr(3) => 
                           pc_bus(3), istr_addr(2) => pc_bus(2), istr_addr(1) 
                           => pc_bus(1), istr_addr(0) => pc_bus(0), 
                           istr_val(31) => ir_bus(31), istr_val(30) => 
                           ir_bus(30), istr_val(29) => ir_bus(29), istr_val(28)
                           => ir_bus(28), istr_val(27) => ir_bus(27), 
                           istr_val(26) => ir_bus(26), istr_val(25) => 
                           ir_bus(25), istr_val(24) => ir_bus(24), istr_val(23)
                           => ir_bus(23), istr_val(22) => ir_bus(22), 
                           istr_val(21) => ir_bus(21), istr_val(20) => 
                           ir_bus(20), istr_val(19) => ir_bus(19), istr_val(18)
                           => ir_bus(18), istr_val(17) => ir_bus(17), 
                           istr_val(16) => ir_bus(16), istr_val(15) => 
                           ir_bus(15), istr_val(14) => ir_bus(14), istr_val(13)
                           => ir_bus(13), istr_val(12) => ir_bus(12), 
                           istr_val(11) => ir_bus(11), istr_val(10) => 
                           ir_bus(10), istr_val(9) => ir_bus(9), istr_val(8) =>
                           ir_bus(8), istr_val(7) => ir_bus(7), istr_val(6) => 
                           ir_bus(6), istr_val(5) => ir_bus(5), istr_val(4) => 
                           ir_bus(4), istr_val(3) => ir_bus(3), istr_val(2) => 
                           ir_bus(2), istr_val(1) => ir_bus(1), istr_val(0) => 
                           ir_bus(0), ir_out(31) => ir_31_port, ir_out(30) => 
                           ir_30_port, ir_out(29) => ir_29_port, ir_out(28) => 
                           ir_28_port, ir_out(27) => ir_27_port, ir_out(26) => 
                           ir_26_port, ir_out(25) => ir_25_port, ir_out(24) => 
                           ir_24_port, ir_out(23) => ir_23_port, ir_out(22) => 
                           ir_22_port, ir_out(21) => ir_21_port, ir_out(20) => 
                           ir_20_port, ir_out(19) => ir_19_port, ir_out(18) => 
                           ir_18_port, ir_out(17) => ir_17_port, ir_out(16) => 
                           ir_16_port, ir_out(15) => ir_15_port, ir_out(14) => 
                           ir_14_port, ir_out(13) => ir_13_port, ir_out(12) => 
                           ir_12_port, ir_out(11) => ir_11_port, ir_out(10) => 
                           ir_10_port, ir_out(9) => ir_9_port, ir_out(8) => 
                           ir_8_port, ir_out(7) => ir_7_port, ir_out(6) => 
                           ir_6_port, ir_out(5) => ir_5_port, ir_out(4) => 
                           ir_4_port, ir_out(3) => ir_3_port, ir_out(2) => 
                           ir_2_port, ir_out(1) => ir_1_port, ir_out(0) => 
                           ir_0_port, pc_out(31) => pc_31_port, pc_out(30) => 
                           pc_30_port, pc_out(29) => pc_29_port, pc_out(28) => 
                           pc_28_port, pc_out(27) => pc_27_port, pc_out(26) => 
                           pc_26_port, pc_out(25) => pc_25_port, pc_out(24) => 
                           pc_24_port, pc_out(23) => pc_23_port, pc_out(22) => 
                           pc_22_port, pc_out(21) => pc_21_port, pc_out(20) => 
                           pc_20_port, pc_out(19) => pc_19_port, pc_out(18) => 
                           pc_18_port, pc_out(17) => pc_17_port, pc_out(16) => 
                           pc_16_port, pc_out(15) => pc_15_port, pc_out(14) => 
                           pc_14_port, pc_out(13) => pc_13_port, pc_out(12) => 
                           pc_12_port, pc_out(11) => pc_11_port, pc_out(10) => 
                           pc_10_port, pc_out(9) => pc_9_port, pc_out(8) => 
                           pc_8_port, pc_out(7) => pc_7_port, pc_out(6) => 
                           pc_6_port, pc_out(5) => pc_5_port, pc_out(4) => 
                           pc_4_port, pc_out(3) => pc_3_port, pc_out(2) => 
                           pc_2_port, pc_out(1) => pc_1_port, pc_out(0) => 
                           pc_0_port, reg_a_out(31) => reg_a_val_31_port, 
                           reg_a_out(30) => reg_a_val_30_port, reg_a_out(29) =>
                           reg_a_val_29_port, reg_a_out(28) => 
                           reg_a_val_28_port, reg_a_out(27) => 
                           reg_a_val_27_port, reg_a_out(26) => 
                           reg_a_val_26_port, reg_a_out(25) => 
                           reg_a_val_25_port, reg_a_out(24) => 
                           reg_a_val_24_port, reg_a_out(23) => 
                           reg_a_val_23_port, reg_a_out(22) => 
                           reg_a_val_22_port, reg_a_out(21) => 
                           reg_a_val_21_port, reg_a_out(20) => 
                           reg_a_val_20_port, reg_a_out(19) => 
                           reg_a_val_19_port, reg_a_out(18) => 
                           reg_a_val_18_port, reg_a_out(17) => 
                           reg_a_val_17_port, reg_a_out(16) => 
                           reg_a_val_16_port, reg_a_out(15) => 
                           reg_a_val_15_port, reg_a_out(14) => 
                           reg_a_val_14_port, reg_a_out(13) => 
                           reg_a_val_13_port, reg_a_out(12) => 
                           reg_a_val_12_port, reg_a_out(11) => 
                           reg_a_val_11_port, reg_a_out(10) => 
                           reg_a_val_10_port, reg_a_out(9) => reg_a_val_9_port,
                           reg_a_out(8) => reg_a_val_8_port, reg_a_out(7) => 
                           reg_a_val_7_port, reg_a_out(6) => reg_a_val_6_port, 
                           reg_a_out(5) => reg_a_val_5_port, reg_a_out(4) => 
                           reg_a_val_4_port, reg_a_out(3) => reg_a_val_3_port, 
                           reg_a_out(2) => reg_a_val_2_port, reg_a_out(1) => 
                           reg_a_val_1_port, reg_a_out(0) => reg_a_val_0_port, 
                           ld_a_out(31) => ld_a_val_31_port, ld_a_out(30) => 
                           ld_a_val_30_port, ld_a_out(29) => ld_a_val_29_port, 
                           ld_a_out(28) => ld_a_val_28_port, ld_a_out(27) => 
                           ld_a_val_27_port, ld_a_out(26) => ld_a_val_26_port, 
                           ld_a_out(25) => ld_a_val_25_port, ld_a_out(24) => 
                           ld_a_val_24_port, ld_a_out(23) => ld_a_val_23_port, 
                           ld_a_out(22) => ld_a_val_22_port, ld_a_out(21) => 
                           ld_a_val_21_port, ld_a_out(20) => ld_a_val_20_port, 
                           ld_a_out(19) => ld_a_val_19_port, ld_a_out(18) => 
                           ld_a_val_18_port, ld_a_out(17) => ld_a_val_17_port, 
                           ld_a_out(16) => ld_a_val_16_port, ld_a_out(15) => 
                           ld_a_val_15_port, ld_a_out(14) => ld_a_val_14_port, 
                           ld_a_out(13) => ld_a_val_13_port, ld_a_out(12) => 
                           ld_a_val_12_port, ld_a_out(11) => ld_a_val_11_port, 
                           ld_a_out(10) => ld_a_val_10_port, ld_a_out(9) => 
                           ld_a_val_9_port, ld_a_out(8) => ld_a_val_8_port, 
                           ld_a_out(7) => ld_a_val_7_port, ld_a_out(6) => 
                           ld_a_val_6_port, ld_a_out(5) => ld_a_val_5_port, 
                           ld_a_out(4) => ld_a_val_4_port, ld_a_out(3) => 
                           ld_a_val_3_port, ld_a_out(2) => ld_a_val_2_port, 
                           ld_a_out(1) => ld_a_val_1_port, ld_a_out(0) => 
                           ld_a_val_0_port, data_addr(31) => addr_bus(31), 
                           data_addr(30) => addr_bus(30), data_addr(29) => 
                           addr_bus(29), data_addr(28) => addr_bus(28), 
                           data_addr(27) => addr_bus(27), data_addr(26) => 
                           addr_bus(26), data_addr(25) => addr_bus(25), 
                           data_addr(24) => addr_bus(24), data_addr(23) => 
                           addr_bus(23), data_addr(22) => addr_bus(22), 
                           data_addr(21) => addr_bus(21), data_addr(20) => 
                           addr_bus(20), data_addr(19) => addr_bus(19), 
                           data_addr(18) => addr_bus(18), data_addr(17) => 
                           addr_bus(17), data_addr(16) => addr_bus(16), 
                           data_addr(15) => addr_bus(15), data_addr(14) => 
                           addr_bus(14), data_addr(13) => addr_bus(13), 
                           data_addr(12) => addr_bus(12), data_addr(11) => 
                           addr_bus(11), data_addr(10) => addr_bus(10), 
                           data_addr(9) => addr_bus(9), data_addr(8) => 
                           addr_bus(8), data_addr(7) => addr_bus(7), 
                           data_addr(6) => addr_bus(6), data_addr(5) => 
                           addr_bus(5), data_addr(4) => addr_bus(4), 
                           data_addr(3) => addr_bus(3), data_addr(2) => 
                           addr_bus(2), data_addr(1) => addr_bus(1), 
                           data_addr(0) => addr_bus(0), data_i_val(31) => 
                           do_bus(31), data_i_val(30) => do_bus(30), 
                           data_i_val(29) => do_bus(29), data_i_val(28) => 
                           do_bus(28), data_i_val(27) => do_bus(27), 
                           data_i_val(26) => do_bus(26), data_i_val(25) => 
                           do_bus(25), data_i_val(24) => do_bus(24), 
                           data_i_val(23) => do_bus(23), data_i_val(22) => 
                           do_bus(22), data_i_val(21) => do_bus(21), 
                           data_i_val(20) => do_bus(20), data_i_val(19) => 
                           do_bus(19), data_i_val(18) => do_bus(18), 
                           data_i_val(17) => do_bus(17), data_i_val(16) => 
                           do_bus(16), data_i_val(15) => do_bus(15), 
                           data_i_val(14) => do_bus(14), data_i_val(13) => 
                           do_bus(13), data_i_val(12) => do_bus(12), 
                           data_i_val(11) => do_bus(11), data_i_val(10) => 
                           do_bus(10), data_i_val(9) => do_bus(9), 
                           data_i_val(8) => do_bus(8), data_i_val(7) => 
                           do_bus(7), data_i_val(6) => do_bus(6), data_i_val(5)
                           => do_bus(5), data_i_val(4) => do_bus(4), 
                           data_i_val(3) => do_bus(3), data_i_val(2) => 
                           do_bus(2), data_i_val(1) => do_bus(1), data_i_val(0)
                           => do_bus(0), data_o_val(31) => di_bus(31), 
                           data_o_val(30) => di_bus(30), data_o_val(29) => 
                           di_bus(29), data_o_val(28) => di_bus(28), 
                           data_o_val(27) => di_bus(27), data_o_val(26) => 
                           di_bus(26), data_o_val(25) => di_bus(25), 
                           data_o_val(24) => di_bus(24), data_o_val(23) => 
                           di_bus(23), data_o_val(22) => di_bus(22), 
                           data_o_val(21) => di_bus(21), data_o_val(20) => 
                           di_bus(20), data_o_val(19) => di_bus(19), 
                           data_o_val(18) => di_bus(18), data_o_val(17) => 
                           di_bus(17), data_o_val(16) => di_bus(16), 
                           data_o_val(15) => di_bus(15), data_o_val(14) => 
                           di_bus(14), data_o_val(13) => di_bus(13), 
                           data_o_val(12) => di_bus(12), data_o_val(11) => 
                           di_bus(11), data_o_val(10) => di_bus(10), 
                           data_o_val(9) => di_bus(9), data_o_val(8) => 
                           di_bus(8), data_o_val(7) => di_bus(7), data_o_val(6)
                           => di_bus(6), data_o_val(5) => di_bus(5), 
                           data_o_val(4) => di_bus(4), data_o_val(3) => 
                           di_bus(3), data_o_val(2) => di_bus(2), data_o_val(1)
                           => di_bus(1), data_o_val(0) => di_bus(0), cw(19) => 
                           cw_19_port, cw(18) => cw_18_port, cw(17) => 
                           cw_17_port, cw(16) => cw_16_port, cw(15) => 
                           cw_15_port, cw(14) => cw_14_port, cw(13) => 
                           cw_13_port, cw(12) => cw_12_port, cw(11) => 
                           cw_11_port, cw(10) => cw_10_port, cw(9) => cw_9_port
                           , cw(8) => cw_8_port, cw(7) => cw_7_port, cw(6) => 
                           cw_6_port, cw(5) => cw_5_port, cw(4) => cw_4_port, 
                           cw(3) => cw_3_port, cw(2) => cw_2_port, cw(1) => 
                           cw_1_port, cw(0) => en_iram_port, dr_cw(3) => 
                           dr_cw(3), dr_cw(2) => dr_cw(2), dr_cw(1) => dr_cw(1)
                           , dr_cw(0) => dr_cw(0), calu(4) => calu_4_port, 
                           calu(3) => calu_3_port, calu(2) => calu_2_port, 
                           calu(1) => calu_1_port, calu(0) => calu_0_port, 
                           sig_bal => sig_bal, sig_bpw => sig_bpw, sig_jral => 
                           sig_jral, sig_ral => sig_ral, sig_mul => sig_mul, 
                           sig_div => sig_div, sig_sqrt => sig_sqrt);

end SYN_dlx_arch;
