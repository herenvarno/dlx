
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity StallGenerator_CWRD_SIZE20_DW01_inc_5 is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end StallGenerator_CWRD_SIZE20_DW01_inc_5;

architecture SYN_rpl of StallGenerator_CWRD_SIZE20_DW01_inc_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port : std_logic;

begin
   
   U1_1_30 : HA_X1 port map( A => A(30), B => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_1_29 : HA_X1 port map( A => A(29), B => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_1_28 : HA_X1 port map( A => A(28), B => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_1_27 : HA_X1 port map( A => A(27), B => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_1_26 : HA_X1 port map( A => A(26), B => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_1_25 : HA_X1 port map( A => A(25), B => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_1_24 : HA_X1 port map( A => A(24), B => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_1_23 : HA_X1 port map( A => A(23), B => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_1_22 : HA_X1 port map( A => A(22), B => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_1_21 : HA_X1 port map( A => A(21), B => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_1_20 : HA_X1 port map( A => A(20), B => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_1_19 : HA_X1 port map( A => A(19), B => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_1_18 : HA_X1 port map( A => A(18), B => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_1_17 : HA_X1 port map( A => A(17), B => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_1_16 : HA_X1 port map( A => A(16), B => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_1_15 : HA_X1 port map( A => A(15), B => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : XOR2_X1 port map( A => carry_31_port, B => A(31), Z => SUM(31));
   U2 : INV_X1 port map( A => A(0), ZN => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity StallGenerator_CWRD_SIZE20_DW01_inc_4 is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end StallGenerator_CWRD_SIZE20_DW01_inc_4;

architecture SYN_rpl of StallGenerator_CWRD_SIZE20_DW01_inc_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port : std_logic;

begin
   
   U1_1_30 : HA_X1 port map( A => A(30), B => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_1_29 : HA_X1 port map( A => A(29), B => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_1_28 : HA_X1 port map( A => A(28), B => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_1_27 : HA_X1 port map( A => A(27), B => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_1_26 : HA_X1 port map( A => A(26), B => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_1_25 : HA_X1 port map( A => A(25), B => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_1_24 : HA_X1 port map( A => A(24), B => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_1_23 : HA_X1 port map( A => A(23), B => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_1_22 : HA_X1 port map( A => A(22), B => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_1_21 : HA_X1 port map( A => A(21), B => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_1_20 : HA_X1 port map( A => A(20), B => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_1_19 : HA_X1 port map( A => A(19), B => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_1_18 : HA_X1 port map( A => A(18), B => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_1_17 : HA_X1 port map( A => A(17), B => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_1_16 : HA_X1 port map( A => A(16), B => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_1_15 : HA_X1 port map( A => A(15), B => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : XOR2_X1 port map( A => carry_31_port, B => A(31), Z => SUM(31));
   U2 : INV_X1 port map( A => A(0), ZN => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity StallGenerator_CWRD_SIZE20_DW01_inc_3 is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end StallGenerator_CWRD_SIZE20_DW01_inc_3;

architecture SYN_rpl of StallGenerator_CWRD_SIZE20_DW01_inc_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port : std_logic;

begin
   
   U1_1_30 : HA_X1 port map( A => A(30), B => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_1_29 : HA_X1 port map( A => A(29), B => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_1_28 : HA_X1 port map( A => A(28), B => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_1_27 : HA_X1 port map( A => A(27), B => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_1_26 : HA_X1 port map( A => A(26), B => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_1_25 : HA_X1 port map( A => A(25), B => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_1_24 : HA_X1 port map( A => A(24), B => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_1_23 : HA_X1 port map( A => A(23), B => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_1_22 : HA_X1 port map( A => A(22), B => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_1_21 : HA_X1 port map( A => A(21), B => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_1_20 : HA_X1 port map( A => A(20), B => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_1_19 : HA_X1 port map( A => A(19), B => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_1_18 : HA_X1 port map( A => A(18), B => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_1_17 : HA_X1 port map( A => A(17), B => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_1_16 : HA_X1 port map( A => A(16), B => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_1_15 : HA_X1 port map( A => A(15), B => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : XOR2_X1 port map( A => carry_31_port, B => A(31), Z => SUM(31));
   U2 : INV_X1 port map( A => A(0), ZN => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity StallGenerator_CWRD_SIZE20_DW01_inc_2 is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end StallGenerator_CWRD_SIZE20_DW01_inc_2;

architecture SYN_rpl of StallGenerator_CWRD_SIZE20_DW01_inc_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port : std_logic;

begin
   
   U1_1_30 : HA_X1 port map( A => A(30), B => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_1_29 : HA_X1 port map( A => A(29), B => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_1_28 : HA_X1 port map( A => A(28), B => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_1_27 : HA_X1 port map( A => A(27), B => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_1_26 : HA_X1 port map( A => A(26), B => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_1_25 : HA_X1 port map( A => A(25), B => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_1_24 : HA_X1 port map( A => A(24), B => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_1_23 : HA_X1 port map( A => A(23), B => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_1_22 : HA_X1 port map( A => A(22), B => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_1_21 : HA_X1 port map( A => A(21), B => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_1_20 : HA_X1 port map( A => A(20), B => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_1_19 : HA_X1 port map( A => A(19), B => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_1_18 : HA_X1 port map( A => A(18), B => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_1_17 : HA_X1 port map( A => A(17), B => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_1_16 : HA_X1 port map( A => A(16), B => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_1_15 : HA_X1 port map( A => A(15), B => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : XOR2_X1 port map( A => carry_31_port, B => A(31), Z => SUM(31));
   U2 : INV_X1 port map( A => A(0), ZN => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity StallGenerator_CWRD_SIZE20_DW01_inc_1 is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end StallGenerator_CWRD_SIZE20_DW01_inc_1;

architecture SYN_rpl of StallGenerator_CWRD_SIZE20_DW01_inc_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port : std_logic;

begin
   
   U1_1_30 : HA_X1 port map( A => A(30), B => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_1_29 : HA_X1 port map( A => A(29), B => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_1_28 : HA_X1 port map( A => A(28), B => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_1_27 : HA_X1 port map( A => A(27), B => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_1_26 : HA_X1 port map( A => A(26), B => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_1_25 : HA_X1 port map( A => A(25), B => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_1_24 : HA_X1 port map( A => A(24), B => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_1_23 : HA_X1 port map( A => A(23), B => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_1_22 : HA_X1 port map( A => A(22), B => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_1_21 : HA_X1 port map( A => A(21), B => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_1_20 : HA_X1 port map( A => A(20), B => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_1_19 : HA_X1 port map( A => A(19), B => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_1_18 : HA_X1 port map( A => A(18), B => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_1_17 : HA_X1 port map( A => A(17), B => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_1_16 : HA_X1 port map( A => A(16), B => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_1_15 : HA_X1 port map( A => A(15), B => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : XOR2_X1 port map( A => carry_31_port, B => A(31), Z => SUM(31));
   U2 : INV_X1 port map( A => A(0), ZN => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity StallGenerator_CWRD_SIZE20_DW01_inc_0 is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end StallGenerator_CWRD_SIZE20_DW01_inc_0;

architecture SYN_rpl of StallGenerator_CWRD_SIZE20_DW01_inc_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port : std_logic;

begin
   
   U1_1_30 : HA_X1 port map( A => A(30), B => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_1_29 : HA_X1 port map( A => A(29), B => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_1_28 : HA_X1 port map( A => A(28), B => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_1_27 : HA_X1 port map( A => A(27), B => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_1_26 : HA_X1 port map( A => A(26), B => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_1_25 : HA_X1 port map( A => A(25), B => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_1_24 : HA_X1 port map( A => A(24), B => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_1_23 : HA_X1 port map( A => A(23), B => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_1_22 : HA_X1 port map( A => A(22), B => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_1_21 : HA_X1 port map( A => A(21), B => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_1_20 : HA_X1 port map( A => A(20), B => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_1_19 : HA_X1 port map( A => A(19), B => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_1_18 : HA_X1 port map( A => A(18), B => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_1_17 : HA_X1 port map( A => A(17), B => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_1_16 : HA_X1 port map( A => A(16), B => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_1_15 : HA_X1 port map( A => A(15), B => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : XOR2_X1 port map( A => carry_31_port, B => A(31), Z => SUM(31));
   U2 : INV_X1 port map( A => A(0), ZN => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Shifter_DATA_SIZE32_DW_rbsh_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end Shifter_DATA_SIZE32_DW_rbsh_0;

architecture SYN_mx2 of Shifter_DATA_SIZE32_DW_rbsh_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal MR_int_1_31_port, MR_int_1_30_port, MR_int_1_29_port, 
      MR_int_1_28_port, MR_int_1_27_port, MR_int_1_26_port, MR_int_1_25_port, 
      MR_int_1_24_port, MR_int_1_23_port, MR_int_1_22_port, MR_int_1_21_port, 
      MR_int_1_20_port, MR_int_1_19_port, MR_int_1_18_port, MR_int_1_17_port, 
      MR_int_1_16_port, MR_int_1_15_port, MR_int_1_14_port, MR_int_1_13_port, 
      MR_int_1_12_port, MR_int_1_11_port, MR_int_1_10_port, MR_int_1_9_port, 
      MR_int_1_8_port, MR_int_1_7_port, MR_int_1_6_port, MR_int_1_5_port, 
      MR_int_1_4_port, MR_int_1_3_port, MR_int_1_2_port, MR_int_1_1_port, 
      MR_int_1_0_port, MR_int_2_31_port, MR_int_2_30_port, MR_int_2_29_port, 
      MR_int_2_28_port, MR_int_2_27_port, MR_int_2_26_port, MR_int_2_25_port, 
      MR_int_2_24_port, MR_int_2_23_port, MR_int_2_22_port, MR_int_2_21_port, 
      MR_int_2_20_port, MR_int_2_19_port, MR_int_2_18_port, MR_int_2_17_port, 
      MR_int_2_16_port, MR_int_2_15_port, MR_int_2_14_port, MR_int_2_13_port, 
      MR_int_2_12_port, MR_int_2_11_port, MR_int_2_10_port, MR_int_2_9_port, 
      MR_int_2_8_port, MR_int_2_7_port, MR_int_2_6_port, MR_int_2_5_port, 
      MR_int_2_4_port, MR_int_2_3_port, MR_int_2_2_port, MR_int_2_1_port, 
      MR_int_2_0_port, MR_int_3_31_port, MR_int_3_30_port, MR_int_3_29_port, 
      MR_int_3_28_port, MR_int_3_27_port, MR_int_3_26_port, MR_int_3_25_port, 
      MR_int_3_24_port, MR_int_3_23_port, MR_int_3_22_port, MR_int_3_21_port, 
      MR_int_3_20_port, MR_int_3_19_port, MR_int_3_18_port, MR_int_3_17_port, 
      MR_int_3_16_port, MR_int_3_15_port, MR_int_3_14_port, MR_int_3_13_port, 
      MR_int_3_12_port, MR_int_3_11_port, MR_int_3_10_port, MR_int_3_9_port, 
      MR_int_3_8_port, MR_int_3_7_port, MR_int_3_6_port, MR_int_3_5_port, 
      MR_int_3_4_port, MR_int_3_3_port, MR_int_3_2_port, MR_int_3_1_port, 
      MR_int_3_0_port, MR_int_4_31_port, MR_int_4_30_port, MR_int_4_29_port, 
      MR_int_4_28_port, MR_int_4_27_port, MR_int_4_26_port, MR_int_4_25_port, 
      MR_int_4_24_port, MR_int_4_23_port, MR_int_4_22_port, MR_int_4_21_port, 
      MR_int_4_20_port, MR_int_4_19_port, MR_int_4_18_port, MR_int_4_17_port, 
      MR_int_4_16_port, MR_int_4_15_port, MR_int_4_14_port, MR_int_4_13_port, 
      MR_int_4_12_port, MR_int_4_11_port, MR_int_4_10_port, MR_int_4_9_port, 
      MR_int_4_8_port, MR_int_4_7_port, MR_int_4_6_port, MR_int_4_5_port, 
      MR_int_4_4_port, MR_int_4_3_port, MR_int_4_2_port, MR_int_4_1_port, 
      MR_int_4_0_port, n1, n2, n3 : std_logic;

begin
   
   M1_4_31 : MUX2_X1 port map( A => MR_int_4_31_port, B => MR_int_4_15_port, S 
                           => n3, Z => B(31));
   M1_4_30 : MUX2_X1 port map( A => MR_int_4_30_port, B => MR_int_4_14_port, S 
                           => n3, Z => B(30));
   M1_4_29 : MUX2_X1 port map( A => MR_int_4_29_port, B => MR_int_4_13_port, S 
                           => n3, Z => B(29));
   M1_4_28 : MUX2_X1 port map( A => MR_int_4_28_port, B => MR_int_4_12_port, S 
                           => n3, Z => B(28));
   M1_4_27 : MUX2_X1 port map( A => MR_int_4_27_port, B => MR_int_4_11_port, S 
                           => n3, Z => B(27));
   M1_4_26 : MUX2_X1 port map( A => MR_int_4_26_port, B => MR_int_4_10_port, S 
                           => n3, Z => B(26));
   M1_4_25 : MUX2_X1 port map( A => MR_int_4_25_port, B => MR_int_4_9_port, S 
                           => n3, Z => B(25));
   M1_4_24 : MUX2_X1 port map( A => MR_int_4_24_port, B => MR_int_4_8_port, S 
                           => n3, Z => B(24));
   M1_4_23 : MUX2_X1 port map( A => MR_int_4_23_port, B => MR_int_4_7_port, S 
                           => n2, Z => B(23));
   M1_4_22 : MUX2_X1 port map( A => MR_int_4_22_port, B => MR_int_4_6_port, S 
                           => n2, Z => B(22));
   M1_4_21 : MUX2_X1 port map( A => MR_int_4_21_port, B => MR_int_4_5_port, S 
                           => n2, Z => B(21));
   M1_4_20 : MUX2_X1 port map( A => MR_int_4_20_port, B => MR_int_4_4_port, S 
                           => n2, Z => B(20));
   M1_4_19 : MUX2_X1 port map( A => MR_int_4_19_port, B => MR_int_4_3_port, S 
                           => n2, Z => B(19));
   M1_4_18 : MUX2_X1 port map( A => MR_int_4_18_port, B => MR_int_4_2_port, S 
                           => n2, Z => B(18));
   M1_4_17 : MUX2_X1 port map( A => MR_int_4_17_port, B => MR_int_4_1_port, S 
                           => n2, Z => B(17));
   M1_4_16 : MUX2_X1 port map( A => MR_int_4_16_port, B => MR_int_4_0_port, S 
                           => n2, Z => B(16));
   M1_4_15 : MUX2_X1 port map( A => MR_int_4_15_port, B => MR_int_4_31_port, S 
                           => n2, Z => B(15));
   M1_4_14 : MUX2_X1 port map( A => MR_int_4_14_port, B => MR_int_4_30_port, S 
                           => n2, Z => B(14));
   M1_4_13 : MUX2_X1 port map( A => MR_int_4_13_port, B => MR_int_4_29_port, S 
                           => n2, Z => B(13));
   M1_4_12 : MUX2_X1 port map( A => MR_int_4_12_port, B => MR_int_4_28_port, S 
                           => n2, Z => B(12));
   M1_4_11 : MUX2_X1 port map( A => MR_int_4_11_port, B => MR_int_4_27_port, S 
                           => n1, Z => B(11));
   M1_4_10 : MUX2_X1 port map( A => MR_int_4_10_port, B => MR_int_4_26_port, S 
                           => n1, Z => B(10));
   M1_4_9 : MUX2_X1 port map( A => MR_int_4_9_port, B => MR_int_4_25_port, S =>
                           n1, Z => B(9));
   M1_4_8 : MUX2_X1 port map( A => MR_int_4_8_port, B => MR_int_4_24_port, S =>
                           n1, Z => B(8));
   M1_4_7 : MUX2_X1 port map( A => MR_int_4_7_port, B => MR_int_4_23_port, S =>
                           n1, Z => B(7));
   M1_4_6 : MUX2_X1 port map( A => MR_int_4_6_port, B => MR_int_4_22_port, S =>
                           n1, Z => B(6));
   M1_4_5 : MUX2_X1 port map( A => MR_int_4_5_port, B => MR_int_4_21_port, S =>
                           n1, Z => B(5));
   M1_4_4 : MUX2_X1 port map( A => MR_int_4_4_port, B => MR_int_4_20_port, S =>
                           n1, Z => B(4));
   M1_4_3 : MUX2_X1 port map( A => MR_int_4_3_port, B => MR_int_4_19_port, S =>
                           n1, Z => B(3));
   M1_4_2 : MUX2_X1 port map( A => MR_int_4_2_port, B => MR_int_4_18_port, S =>
                           n1, Z => B(2));
   M1_4_1 : MUX2_X1 port map( A => MR_int_4_1_port, B => MR_int_4_17_port, S =>
                           n1, Z => B(1));
   M1_4_0 : MUX2_X1 port map( A => MR_int_4_0_port, B => MR_int_4_16_port, S =>
                           n1, Z => B(0));
   M1_3_31_0 : MUX2_X1 port map( A => MR_int_3_31_port, B => MR_int_3_7_port, S
                           => SH(3), Z => MR_int_4_31_port);
   M1_3_30_0 : MUX2_X1 port map( A => MR_int_3_30_port, B => MR_int_3_6_port, S
                           => SH(3), Z => MR_int_4_30_port);
   M1_3_29_0 : MUX2_X1 port map( A => MR_int_3_29_port, B => MR_int_3_5_port, S
                           => SH(3), Z => MR_int_4_29_port);
   M1_3_28_0 : MUX2_X1 port map( A => MR_int_3_28_port, B => MR_int_3_4_port, S
                           => SH(3), Z => MR_int_4_28_port);
   M1_3_27_0 : MUX2_X1 port map( A => MR_int_3_27_port, B => MR_int_3_3_port, S
                           => SH(3), Z => MR_int_4_27_port);
   M1_3_26_0 : MUX2_X1 port map( A => MR_int_3_26_port, B => MR_int_3_2_port, S
                           => SH(3), Z => MR_int_4_26_port);
   M1_3_25_0 : MUX2_X1 port map( A => MR_int_3_25_port, B => MR_int_3_1_port, S
                           => SH(3), Z => MR_int_4_25_port);
   M1_3_24_0 : MUX2_X1 port map( A => MR_int_3_24_port, B => MR_int_3_0_port, S
                           => SH(3), Z => MR_int_4_24_port);
   M1_3_23_0 : MUX2_X1 port map( A => MR_int_3_23_port, B => MR_int_3_31_port, 
                           S => SH(3), Z => MR_int_4_23_port);
   M1_3_22_0 : MUX2_X1 port map( A => MR_int_3_22_port, B => MR_int_3_30_port, 
                           S => SH(3), Z => MR_int_4_22_port);
   M1_3_21_0 : MUX2_X1 port map( A => MR_int_3_21_port, B => MR_int_3_29_port, 
                           S => SH(3), Z => MR_int_4_21_port);
   M1_3_20_0 : MUX2_X1 port map( A => MR_int_3_20_port, B => MR_int_3_28_port, 
                           S => SH(3), Z => MR_int_4_20_port);
   M1_3_19_0 : MUX2_X1 port map( A => MR_int_3_19_port, B => MR_int_3_27_port, 
                           S => SH(3), Z => MR_int_4_19_port);
   M1_3_18_0 : MUX2_X1 port map( A => MR_int_3_18_port, B => MR_int_3_26_port, 
                           S => SH(3), Z => MR_int_4_18_port);
   M1_3_17_0 : MUX2_X1 port map( A => MR_int_3_17_port, B => MR_int_3_25_port, 
                           S => SH(3), Z => MR_int_4_17_port);
   M1_3_16_0 : MUX2_X1 port map( A => MR_int_3_16_port, B => MR_int_3_24_port, 
                           S => SH(3), Z => MR_int_4_16_port);
   M1_3_15_0 : MUX2_X1 port map( A => MR_int_3_15_port, B => MR_int_3_23_port, 
                           S => SH(3), Z => MR_int_4_15_port);
   M1_3_14_0 : MUX2_X1 port map( A => MR_int_3_14_port, B => MR_int_3_22_port, 
                           S => SH(3), Z => MR_int_4_14_port);
   M1_3_13_0 : MUX2_X1 port map( A => MR_int_3_13_port, B => MR_int_3_21_port, 
                           S => SH(3), Z => MR_int_4_13_port);
   M1_3_12_0 : MUX2_X1 port map( A => MR_int_3_12_port, B => MR_int_3_20_port, 
                           S => SH(3), Z => MR_int_4_12_port);
   M1_3_11_0 : MUX2_X1 port map( A => MR_int_3_11_port, B => MR_int_3_19_port, 
                           S => SH(3), Z => MR_int_4_11_port);
   M1_3_10_0 : MUX2_X1 port map( A => MR_int_3_10_port, B => MR_int_3_18_port, 
                           S => SH(3), Z => MR_int_4_10_port);
   M1_3_9_0 : MUX2_X1 port map( A => MR_int_3_9_port, B => MR_int_3_17_port, S 
                           => SH(3), Z => MR_int_4_9_port);
   M1_3_8_0 : MUX2_X1 port map( A => MR_int_3_8_port, B => MR_int_3_16_port, S 
                           => SH(3), Z => MR_int_4_8_port);
   M1_3_7 : MUX2_X1 port map( A => MR_int_3_7_port, B => MR_int_3_15_port, S =>
                           SH(3), Z => MR_int_4_7_port);
   M1_3_6 : MUX2_X1 port map( A => MR_int_3_6_port, B => MR_int_3_14_port, S =>
                           SH(3), Z => MR_int_4_6_port);
   M1_3_5 : MUX2_X1 port map( A => MR_int_3_5_port, B => MR_int_3_13_port, S =>
                           SH(3), Z => MR_int_4_5_port);
   M1_3_4 : MUX2_X1 port map( A => MR_int_3_4_port, B => MR_int_3_12_port, S =>
                           SH(3), Z => MR_int_4_4_port);
   M1_3_3 : MUX2_X1 port map( A => MR_int_3_3_port, B => MR_int_3_11_port, S =>
                           SH(3), Z => MR_int_4_3_port);
   M1_3_2 : MUX2_X1 port map( A => MR_int_3_2_port, B => MR_int_3_10_port, S =>
                           SH(3), Z => MR_int_4_2_port);
   M1_3_1 : MUX2_X1 port map( A => MR_int_3_1_port, B => MR_int_3_9_port, S => 
                           SH(3), Z => MR_int_4_1_port);
   M1_3_0 : MUX2_X1 port map( A => MR_int_3_0_port, B => MR_int_3_8_port, S => 
                           SH(3), Z => MR_int_4_0_port);
   M1_2_31_0 : MUX2_X1 port map( A => MR_int_2_31_port, B => MR_int_2_3_port, S
                           => SH(2), Z => MR_int_3_31_port);
   M1_2_30_0 : MUX2_X1 port map( A => MR_int_2_30_port, B => MR_int_2_2_port, S
                           => SH(2), Z => MR_int_3_30_port);
   M1_2_29_0 : MUX2_X1 port map( A => MR_int_2_29_port, B => MR_int_2_1_port, S
                           => SH(2), Z => MR_int_3_29_port);
   M1_2_28_0 : MUX2_X1 port map( A => MR_int_2_28_port, B => MR_int_2_0_port, S
                           => SH(2), Z => MR_int_3_28_port);
   M1_2_27_0 : MUX2_X1 port map( A => MR_int_2_27_port, B => MR_int_2_31_port, 
                           S => SH(2), Z => MR_int_3_27_port);
   M1_2_26_0 : MUX2_X1 port map( A => MR_int_2_26_port, B => MR_int_2_30_port, 
                           S => SH(2), Z => MR_int_3_26_port);
   M1_2_25_0 : MUX2_X1 port map( A => MR_int_2_25_port, B => MR_int_2_29_port, 
                           S => SH(2), Z => MR_int_3_25_port);
   M1_2_24_0 : MUX2_X1 port map( A => MR_int_2_24_port, B => MR_int_2_28_port, 
                           S => SH(2), Z => MR_int_3_24_port);
   M1_2_23_0 : MUX2_X1 port map( A => MR_int_2_23_port, B => MR_int_2_27_port, 
                           S => SH(2), Z => MR_int_3_23_port);
   M1_2_22_0 : MUX2_X1 port map( A => MR_int_2_22_port, B => MR_int_2_26_port, 
                           S => SH(2), Z => MR_int_3_22_port);
   M1_2_21_0 : MUX2_X1 port map( A => MR_int_2_21_port, B => MR_int_2_25_port, 
                           S => SH(2), Z => MR_int_3_21_port);
   M1_2_20_0 : MUX2_X1 port map( A => MR_int_2_20_port, B => MR_int_2_24_port, 
                           S => SH(2), Z => MR_int_3_20_port);
   M1_2_19_0 : MUX2_X1 port map( A => MR_int_2_19_port, B => MR_int_2_23_port, 
                           S => SH(2), Z => MR_int_3_19_port);
   M1_2_18_0 : MUX2_X1 port map( A => MR_int_2_18_port, B => MR_int_2_22_port, 
                           S => SH(2), Z => MR_int_3_18_port);
   M1_2_17_0 : MUX2_X1 port map( A => MR_int_2_17_port, B => MR_int_2_21_port, 
                           S => SH(2), Z => MR_int_3_17_port);
   M1_2_16_0 : MUX2_X1 port map( A => MR_int_2_16_port, B => MR_int_2_20_port, 
                           S => SH(2), Z => MR_int_3_16_port);
   M1_2_15_0 : MUX2_X1 port map( A => MR_int_2_15_port, B => MR_int_2_19_port, 
                           S => SH(2), Z => MR_int_3_15_port);
   M1_2_14_0 : MUX2_X1 port map( A => MR_int_2_14_port, B => MR_int_2_18_port, 
                           S => SH(2), Z => MR_int_3_14_port);
   M1_2_13_0 : MUX2_X1 port map( A => MR_int_2_13_port, B => MR_int_2_17_port, 
                           S => SH(2), Z => MR_int_3_13_port);
   M1_2_12_0 : MUX2_X1 port map( A => MR_int_2_12_port, B => MR_int_2_16_port, 
                           S => SH(2), Z => MR_int_3_12_port);
   M1_2_11_0 : MUX2_X1 port map( A => MR_int_2_11_port, B => MR_int_2_15_port, 
                           S => SH(2), Z => MR_int_3_11_port);
   M1_2_10_0 : MUX2_X1 port map( A => MR_int_2_10_port, B => MR_int_2_14_port, 
                           S => SH(2), Z => MR_int_3_10_port);
   M1_2_9_0 : MUX2_X1 port map( A => MR_int_2_9_port, B => MR_int_2_13_port, S 
                           => SH(2), Z => MR_int_3_9_port);
   M1_2_8_0 : MUX2_X1 port map( A => MR_int_2_8_port, B => MR_int_2_12_port, S 
                           => SH(2), Z => MR_int_3_8_port);
   M1_2_7_0 : MUX2_X1 port map( A => MR_int_2_7_port, B => MR_int_2_11_port, S 
                           => SH(2), Z => MR_int_3_7_port);
   M1_2_6_0 : MUX2_X1 port map( A => MR_int_2_6_port, B => MR_int_2_10_port, S 
                           => SH(2), Z => MR_int_3_6_port);
   M1_2_5_0 : MUX2_X1 port map( A => MR_int_2_5_port, B => MR_int_2_9_port, S 
                           => SH(2), Z => MR_int_3_5_port);
   M1_2_4_0 : MUX2_X1 port map( A => MR_int_2_4_port, B => MR_int_2_8_port, S 
                           => SH(2), Z => MR_int_3_4_port);
   M1_2_3 : MUX2_X1 port map( A => MR_int_2_3_port, B => MR_int_2_7_port, S => 
                           SH(2), Z => MR_int_3_3_port);
   M1_2_2 : MUX2_X1 port map( A => MR_int_2_2_port, B => MR_int_2_6_port, S => 
                           SH(2), Z => MR_int_3_2_port);
   M1_2_1 : MUX2_X1 port map( A => MR_int_2_1_port, B => MR_int_2_5_port, S => 
                           SH(2), Z => MR_int_3_1_port);
   M1_2_0 : MUX2_X1 port map( A => MR_int_2_0_port, B => MR_int_2_4_port, S => 
                           SH(2), Z => MR_int_3_0_port);
   M1_1_31_0 : MUX2_X1 port map( A => MR_int_1_31_port, B => MR_int_1_1_port, S
                           => SH(1), Z => MR_int_2_31_port);
   M1_1_30_0 : MUX2_X1 port map( A => MR_int_1_30_port, B => MR_int_1_0_port, S
                           => SH(1), Z => MR_int_2_30_port);
   M1_1_29_0 : MUX2_X1 port map( A => MR_int_1_29_port, B => MR_int_1_31_port, 
                           S => SH(1), Z => MR_int_2_29_port);
   M1_1_28_0 : MUX2_X1 port map( A => MR_int_1_28_port, B => MR_int_1_30_port, 
                           S => SH(1), Z => MR_int_2_28_port);
   M1_1_27_0 : MUX2_X1 port map( A => MR_int_1_27_port, B => MR_int_1_29_port, 
                           S => SH(1), Z => MR_int_2_27_port);
   M1_1_26_0 : MUX2_X1 port map( A => MR_int_1_26_port, B => MR_int_1_28_port, 
                           S => SH(1), Z => MR_int_2_26_port);
   M1_1_25_0 : MUX2_X1 port map( A => MR_int_1_25_port, B => MR_int_1_27_port, 
                           S => SH(1), Z => MR_int_2_25_port);
   M1_1_24_0 : MUX2_X1 port map( A => MR_int_1_24_port, B => MR_int_1_26_port, 
                           S => SH(1), Z => MR_int_2_24_port);
   M1_1_23_0 : MUX2_X1 port map( A => MR_int_1_23_port, B => MR_int_1_25_port, 
                           S => SH(1), Z => MR_int_2_23_port);
   M1_1_22_0 : MUX2_X1 port map( A => MR_int_1_22_port, B => MR_int_1_24_port, 
                           S => SH(1), Z => MR_int_2_22_port);
   M1_1_21_0 : MUX2_X1 port map( A => MR_int_1_21_port, B => MR_int_1_23_port, 
                           S => SH(1), Z => MR_int_2_21_port);
   M1_1_20_0 : MUX2_X1 port map( A => MR_int_1_20_port, B => MR_int_1_22_port, 
                           S => SH(1), Z => MR_int_2_20_port);
   M1_1_19_0 : MUX2_X1 port map( A => MR_int_1_19_port, B => MR_int_1_21_port, 
                           S => SH(1), Z => MR_int_2_19_port);
   M1_1_18_0 : MUX2_X1 port map( A => MR_int_1_18_port, B => MR_int_1_20_port, 
                           S => SH(1), Z => MR_int_2_18_port);
   M1_1_17_0 : MUX2_X1 port map( A => MR_int_1_17_port, B => MR_int_1_19_port, 
                           S => SH(1), Z => MR_int_2_17_port);
   M1_1_16_0 : MUX2_X1 port map( A => MR_int_1_16_port, B => MR_int_1_18_port, 
                           S => SH(1), Z => MR_int_2_16_port);
   M1_1_15_0 : MUX2_X1 port map( A => MR_int_1_15_port, B => MR_int_1_17_port, 
                           S => SH(1), Z => MR_int_2_15_port);
   M1_1_14_0 : MUX2_X1 port map( A => MR_int_1_14_port, B => MR_int_1_16_port, 
                           S => SH(1), Z => MR_int_2_14_port);
   M1_1_13_0 : MUX2_X1 port map( A => MR_int_1_13_port, B => MR_int_1_15_port, 
                           S => SH(1), Z => MR_int_2_13_port);
   M1_1_12_0 : MUX2_X1 port map( A => MR_int_1_12_port, B => MR_int_1_14_port, 
                           S => SH(1), Z => MR_int_2_12_port);
   M1_1_11_0 : MUX2_X1 port map( A => MR_int_1_11_port, B => MR_int_1_13_port, 
                           S => SH(1), Z => MR_int_2_11_port);
   M1_1_10_0 : MUX2_X1 port map( A => MR_int_1_10_port, B => MR_int_1_12_port, 
                           S => SH(1), Z => MR_int_2_10_port);
   M1_1_9_0 : MUX2_X1 port map( A => MR_int_1_9_port, B => MR_int_1_11_port, S 
                           => SH(1), Z => MR_int_2_9_port);
   M1_1_8_0 : MUX2_X1 port map( A => MR_int_1_8_port, B => MR_int_1_10_port, S 
                           => SH(1), Z => MR_int_2_8_port);
   M1_1_7_0 : MUX2_X1 port map( A => MR_int_1_7_port, B => MR_int_1_9_port, S 
                           => SH(1), Z => MR_int_2_7_port);
   M1_1_6_0 : MUX2_X1 port map( A => MR_int_1_6_port, B => MR_int_1_8_port, S 
                           => SH(1), Z => MR_int_2_6_port);
   M1_1_5_0 : MUX2_X1 port map( A => MR_int_1_5_port, B => MR_int_1_7_port, S 
                           => SH(1), Z => MR_int_2_5_port);
   M1_1_4_0 : MUX2_X1 port map( A => MR_int_1_4_port, B => MR_int_1_6_port, S 
                           => SH(1), Z => MR_int_2_4_port);
   M1_1_3_0 : MUX2_X1 port map( A => MR_int_1_3_port, B => MR_int_1_5_port, S 
                           => SH(1), Z => MR_int_2_3_port);
   M1_1_2_0 : MUX2_X1 port map( A => MR_int_1_2_port, B => MR_int_1_4_port, S 
                           => SH(1), Z => MR_int_2_2_port);
   M1_1_1 : MUX2_X1 port map( A => MR_int_1_1_port, B => MR_int_1_3_port, S => 
                           SH(1), Z => MR_int_2_1_port);
   M1_1_0 : MUX2_X1 port map( A => MR_int_1_0_port, B => MR_int_1_2_port, S => 
                           SH(1), Z => MR_int_2_0_port);
   M1_0_31_0 : MUX2_X1 port map( A => A(31), B => A(0), S => SH(0), Z => 
                           MR_int_1_31_port);
   M1_0_30_0 : MUX2_X1 port map( A => A(30), B => A(31), S => SH(0), Z => 
                           MR_int_1_30_port);
   M1_0_29_0 : MUX2_X1 port map( A => A(29), B => A(30), S => SH(0), Z => 
                           MR_int_1_29_port);
   M1_0_28_0 : MUX2_X1 port map( A => A(28), B => A(29), S => SH(0), Z => 
                           MR_int_1_28_port);
   M1_0_27_0 : MUX2_X1 port map( A => A(27), B => A(28), S => SH(0), Z => 
                           MR_int_1_27_port);
   M1_0_26_0 : MUX2_X1 port map( A => A(26), B => A(27), S => SH(0), Z => 
                           MR_int_1_26_port);
   M1_0_25_0 : MUX2_X1 port map( A => A(25), B => A(26), S => SH(0), Z => 
                           MR_int_1_25_port);
   M1_0_24_0 : MUX2_X1 port map( A => A(24), B => A(25), S => SH(0), Z => 
                           MR_int_1_24_port);
   M1_0_23_0 : MUX2_X1 port map( A => A(23), B => A(24), S => SH(0), Z => 
                           MR_int_1_23_port);
   M1_0_22_0 : MUX2_X1 port map( A => A(22), B => A(23), S => SH(0), Z => 
                           MR_int_1_22_port);
   M1_0_21_0 : MUX2_X1 port map( A => A(21), B => A(22), S => SH(0), Z => 
                           MR_int_1_21_port);
   M1_0_20_0 : MUX2_X1 port map( A => A(20), B => A(21), S => SH(0), Z => 
                           MR_int_1_20_port);
   M1_0_19_0 : MUX2_X1 port map( A => A(19), B => A(20), S => SH(0), Z => 
                           MR_int_1_19_port);
   M1_0_18_0 : MUX2_X1 port map( A => A(18), B => A(19), S => SH(0), Z => 
                           MR_int_1_18_port);
   M1_0_17_0 : MUX2_X1 port map( A => A(17), B => A(18), S => SH(0), Z => 
                           MR_int_1_17_port);
   M1_0_16_0 : MUX2_X1 port map( A => A(16), B => A(17), S => SH(0), Z => 
                           MR_int_1_16_port);
   M1_0_15_0 : MUX2_X1 port map( A => A(15), B => A(16), S => SH(0), Z => 
                           MR_int_1_15_port);
   M1_0_14_0 : MUX2_X1 port map( A => A(14), B => A(15), S => SH(0), Z => 
                           MR_int_1_14_port);
   M1_0_13_0 : MUX2_X1 port map( A => A(13), B => A(14), S => SH(0), Z => 
                           MR_int_1_13_port);
   M1_0_12_0 : MUX2_X1 port map( A => A(12), B => A(13), S => SH(0), Z => 
                           MR_int_1_12_port);
   M1_0_11_0 : MUX2_X1 port map( A => A(11), B => A(12), S => SH(0), Z => 
                           MR_int_1_11_port);
   M1_0_10_0 : MUX2_X1 port map( A => A(10), B => A(11), S => SH(0), Z => 
                           MR_int_1_10_port);
   M1_0_9_0 : MUX2_X1 port map( A => A(9), B => A(10), S => SH(0), Z => 
                           MR_int_1_9_port);
   M1_0_8_0 : MUX2_X1 port map( A => A(8), B => A(9), S => SH(0), Z => 
                           MR_int_1_8_port);
   M1_0_7_0 : MUX2_X1 port map( A => A(7), B => A(8), S => SH(0), Z => 
                           MR_int_1_7_port);
   M1_0_6_0 : MUX2_X1 port map( A => A(6), B => A(7), S => SH(0), Z => 
                           MR_int_1_6_port);
   M1_0_5_0 : MUX2_X1 port map( A => A(5), B => A(6), S => SH(0), Z => 
                           MR_int_1_5_port);
   M1_0_4_0 : MUX2_X1 port map( A => A(4), B => A(5), S => SH(0), Z => 
                           MR_int_1_4_port);
   M1_0_3_0 : MUX2_X1 port map( A => A(3), B => A(4), S => SH(0), Z => 
                           MR_int_1_3_port);
   M1_0_2_0 : MUX2_X1 port map( A => A(2), B => A(3), S => SH(0), Z => 
                           MR_int_1_2_port);
   M1_0_1_0 : MUX2_X1 port map( A => A(1), B => A(2), S => SH(0), Z => 
                           MR_int_1_1_port);
   M1_0_0 : MUX2_X1 port map( A => A(0), B => A(1), S => SH(0), Z => 
                           MR_int_1_0_port);
   U2 : BUF_X1 port map( A => SH(4), Z => n1);
   U3 : BUF_X1 port map( A => SH(4), Z => n2);
   U4 : BUF_X1 port map( A => SH(4), Z => n3);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Shifter_DATA_SIZE32_DW_lbsh_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end Shifter_DATA_SIZE32_DW_lbsh_0;

architecture SYN_mx2 of Shifter_DATA_SIZE32_DW_lbsh_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal ML_int_1_31_port, ML_int_1_30_port, ML_int_1_29_port, 
      ML_int_1_28_port, ML_int_1_27_port, ML_int_1_26_port, ML_int_1_25_port, 
      ML_int_1_24_port, ML_int_1_23_port, ML_int_1_22_port, ML_int_1_21_port, 
      ML_int_1_20_port, ML_int_1_19_port, ML_int_1_18_port, ML_int_1_17_port, 
      ML_int_1_16_port, ML_int_1_15_port, ML_int_1_14_port, ML_int_1_13_port, 
      ML_int_1_12_port, ML_int_1_11_port, ML_int_1_10_port, ML_int_1_9_port, 
      ML_int_1_8_port, ML_int_1_7_port, ML_int_1_6_port, ML_int_1_5_port, 
      ML_int_1_4_port, ML_int_1_3_port, ML_int_1_2_port, ML_int_1_1_port, 
      ML_int_1_0_port, ML_int_2_31_port, ML_int_2_30_port, ML_int_2_29_port, 
      ML_int_2_28_port, ML_int_2_27_port, ML_int_2_26_port, ML_int_2_25_port, 
      ML_int_2_24_port, ML_int_2_23_port, ML_int_2_22_port, ML_int_2_21_port, 
      ML_int_2_20_port, ML_int_2_19_port, ML_int_2_18_port, ML_int_2_17_port, 
      ML_int_2_16_port, ML_int_2_15_port, ML_int_2_14_port, ML_int_2_13_port, 
      ML_int_2_12_port, ML_int_2_11_port, ML_int_2_10_port, ML_int_2_9_port, 
      ML_int_2_8_port, ML_int_2_7_port, ML_int_2_6_port, ML_int_2_5_port, 
      ML_int_2_4_port, ML_int_2_3_port, ML_int_2_2_port, ML_int_2_1_port, 
      ML_int_2_0_port, ML_int_3_31_port, ML_int_3_30_port, ML_int_3_29_port, 
      ML_int_3_28_port, ML_int_3_27_port, ML_int_3_26_port, ML_int_3_25_port, 
      ML_int_3_24_port, ML_int_3_23_port, ML_int_3_22_port, ML_int_3_21_port, 
      ML_int_3_20_port, ML_int_3_19_port, ML_int_3_18_port, ML_int_3_17_port, 
      ML_int_3_16_port, ML_int_3_15_port, ML_int_3_14_port, ML_int_3_13_port, 
      ML_int_3_12_port, ML_int_3_11_port, ML_int_3_10_port, ML_int_3_9_port, 
      ML_int_3_8_port, ML_int_3_7_port, ML_int_3_6_port, ML_int_3_5_port, 
      ML_int_3_4_port, ML_int_3_3_port, ML_int_3_2_port, ML_int_3_1_port, 
      ML_int_3_0_port, ML_int_4_31_port, ML_int_4_30_port, ML_int_4_29_port, 
      ML_int_4_28_port, ML_int_4_27_port, ML_int_4_26_port, ML_int_4_25_port, 
      ML_int_4_24_port, ML_int_4_23_port, ML_int_4_22_port, ML_int_4_21_port, 
      ML_int_4_20_port, ML_int_4_19_port, ML_int_4_18_port, ML_int_4_17_port, 
      ML_int_4_16_port, ML_int_4_15_port, ML_int_4_14_port, ML_int_4_13_port, 
      ML_int_4_12_port, ML_int_4_11_port, ML_int_4_10_port, ML_int_4_9_port, 
      ML_int_4_8_port, ML_int_4_7_port, ML_int_4_6_port, ML_int_4_5_port, 
      ML_int_4_4_port, ML_int_4_3_port, ML_int_4_2_port, ML_int_4_1_port, 
      ML_int_4_0_port, n1, n2, n3 : std_logic;

begin
   
   M1_4_31 : MUX2_X1 port map( A => ML_int_4_31_port, B => ML_int_4_15_port, S 
                           => n3, Z => B(31));
   M1_4_30 : MUX2_X1 port map( A => ML_int_4_30_port, B => ML_int_4_14_port, S 
                           => n3, Z => B(30));
   M1_4_29 : MUX2_X1 port map( A => ML_int_4_29_port, B => ML_int_4_13_port, S 
                           => n3, Z => B(29));
   M1_4_28 : MUX2_X1 port map( A => ML_int_4_28_port, B => ML_int_4_12_port, S 
                           => n3, Z => B(28));
   M1_4_27 : MUX2_X1 port map( A => ML_int_4_27_port, B => ML_int_4_11_port, S 
                           => n3, Z => B(27));
   M1_4_26 : MUX2_X1 port map( A => ML_int_4_26_port, B => ML_int_4_10_port, S 
                           => n3, Z => B(26));
   M1_4_25 : MUX2_X1 port map( A => ML_int_4_25_port, B => ML_int_4_9_port, S 
                           => n3, Z => B(25));
   M1_4_24 : MUX2_X1 port map( A => ML_int_4_24_port, B => ML_int_4_8_port, S 
                           => n3, Z => B(24));
   M1_4_23 : MUX2_X1 port map( A => ML_int_4_23_port, B => ML_int_4_7_port, S 
                           => n2, Z => B(23));
   M1_4_22 : MUX2_X1 port map( A => ML_int_4_22_port, B => ML_int_4_6_port, S 
                           => n2, Z => B(22));
   M1_4_21 : MUX2_X1 port map( A => ML_int_4_21_port, B => ML_int_4_5_port, S 
                           => n2, Z => B(21));
   M1_4_20 : MUX2_X1 port map( A => ML_int_4_20_port, B => ML_int_4_4_port, S 
                           => n2, Z => B(20));
   M1_4_19 : MUX2_X1 port map( A => ML_int_4_19_port, B => ML_int_4_3_port, S 
                           => n2, Z => B(19));
   M1_4_18 : MUX2_X1 port map( A => ML_int_4_18_port, B => ML_int_4_2_port, S 
                           => n2, Z => B(18));
   M1_4_17 : MUX2_X1 port map( A => ML_int_4_17_port, B => ML_int_4_1_port, S 
                           => n2, Z => B(17));
   M1_4_16 : MUX2_X1 port map( A => ML_int_4_16_port, B => ML_int_4_0_port, S 
                           => n2, Z => B(16));
   M0_4_15 : MUX2_X1 port map( A => ML_int_4_15_port, B => ML_int_4_31_port, S 
                           => n2, Z => B(15));
   M0_4_14 : MUX2_X1 port map( A => ML_int_4_14_port, B => ML_int_4_30_port, S 
                           => n2, Z => B(14));
   M0_4_13 : MUX2_X1 port map( A => ML_int_4_13_port, B => ML_int_4_29_port, S 
                           => n2, Z => B(13));
   M0_4_12 : MUX2_X1 port map( A => ML_int_4_12_port, B => ML_int_4_28_port, S 
                           => n2, Z => B(12));
   M0_4_11 : MUX2_X1 port map( A => ML_int_4_11_port, B => ML_int_4_27_port, S 
                           => n1, Z => B(11));
   M0_4_10 : MUX2_X1 port map( A => ML_int_4_10_port, B => ML_int_4_26_port, S 
                           => n1, Z => B(10));
   M0_4_9 : MUX2_X1 port map( A => ML_int_4_9_port, B => ML_int_4_25_port, S =>
                           n1, Z => B(9));
   M0_4_8 : MUX2_X1 port map( A => ML_int_4_8_port, B => ML_int_4_24_port, S =>
                           n1, Z => B(8));
   M0_4_7 : MUX2_X1 port map( A => ML_int_4_7_port, B => ML_int_4_23_port, S =>
                           n1, Z => B(7));
   M0_4_6 : MUX2_X1 port map( A => ML_int_4_6_port, B => ML_int_4_22_port, S =>
                           n1, Z => B(6));
   M0_4_5 : MUX2_X1 port map( A => ML_int_4_5_port, B => ML_int_4_21_port, S =>
                           n1, Z => B(5));
   M0_4_4 : MUX2_X1 port map( A => ML_int_4_4_port, B => ML_int_4_20_port, S =>
                           n1, Z => B(4));
   M0_4_3 : MUX2_X1 port map( A => ML_int_4_3_port, B => ML_int_4_19_port, S =>
                           n1, Z => B(3));
   M0_4_2 : MUX2_X1 port map( A => ML_int_4_2_port, B => ML_int_4_18_port, S =>
                           n1, Z => B(2));
   M0_4_1 : MUX2_X1 port map( A => ML_int_4_1_port, B => ML_int_4_17_port, S =>
                           n1, Z => B(1));
   M0_4_0 : MUX2_X1 port map( A => ML_int_4_0_port, B => ML_int_4_16_port, S =>
                           n1, Z => B(0));
   M1_3_31 : MUX2_X1 port map( A => ML_int_3_31_port, B => ML_int_3_23_port, S 
                           => SH(3), Z => ML_int_4_31_port);
   M1_3_30 : MUX2_X1 port map( A => ML_int_3_30_port, B => ML_int_3_22_port, S 
                           => SH(3), Z => ML_int_4_30_port);
   M1_3_29 : MUX2_X1 port map( A => ML_int_3_29_port, B => ML_int_3_21_port, S 
                           => SH(3), Z => ML_int_4_29_port);
   M1_3_28 : MUX2_X1 port map( A => ML_int_3_28_port, B => ML_int_3_20_port, S 
                           => SH(3), Z => ML_int_4_28_port);
   M1_3_27 : MUX2_X1 port map( A => ML_int_3_27_port, B => ML_int_3_19_port, S 
                           => SH(3), Z => ML_int_4_27_port);
   M1_3_26 : MUX2_X1 port map( A => ML_int_3_26_port, B => ML_int_3_18_port, S 
                           => SH(3), Z => ML_int_4_26_port);
   M1_3_25 : MUX2_X1 port map( A => ML_int_3_25_port, B => ML_int_3_17_port, S 
                           => SH(3), Z => ML_int_4_25_port);
   M1_3_24 : MUX2_X1 port map( A => ML_int_3_24_port, B => ML_int_3_16_port, S 
                           => SH(3), Z => ML_int_4_24_port);
   M1_3_23 : MUX2_X1 port map( A => ML_int_3_23_port, B => ML_int_3_15_port, S 
                           => SH(3), Z => ML_int_4_23_port);
   M1_3_22 : MUX2_X1 port map( A => ML_int_3_22_port, B => ML_int_3_14_port, S 
                           => SH(3), Z => ML_int_4_22_port);
   M1_3_21 : MUX2_X1 port map( A => ML_int_3_21_port, B => ML_int_3_13_port, S 
                           => SH(3), Z => ML_int_4_21_port);
   M1_3_20 : MUX2_X1 port map( A => ML_int_3_20_port, B => ML_int_3_12_port, S 
                           => SH(3), Z => ML_int_4_20_port);
   M1_3_19 : MUX2_X1 port map( A => ML_int_3_19_port, B => ML_int_3_11_port, S 
                           => SH(3), Z => ML_int_4_19_port);
   M1_3_18 : MUX2_X1 port map( A => ML_int_3_18_port, B => ML_int_3_10_port, S 
                           => SH(3), Z => ML_int_4_18_port);
   M1_3_17 : MUX2_X1 port map( A => ML_int_3_17_port, B => ML_int_3_9_port, S 
                           => SH(3), Z => ML_int_4_17_port);
   M1_3_16 : MUX2_X1 port map( A => ML_int_3_16_port, B => ML_int_3_8_port, S 
                           => SH(3), Z => ML_int_4_16_port);
   M1_3_15 : MUX2_X1 port map( A => ML_int_3_15_port, B => ML_int_3_7_port, S 
                           => SH(3), Z => ML_int_4_15_port);
   M1_3_14 : MUX2_X1 port map( A => ML_int_3_14_port, B => ML_int_3_6_port, S 
                           => SH(3), Z => ML_int_4_14_port);
   M1_3_13 : MUX2_X1 port map( A => ML_int_3_13_port, B => ML_int_3_5_port, S 
                           => SH(3), Z => ML_int_4_13_port);
   M1_3_12 : MUX2_X1 port map( A => ML_int_3_12_port, B => ML_int_3_4_port, S 
                           => SH(3), Z => ML_int_4_12_port);
   M1_3_11 : MUX2_X1 port map( A => ML_int_3_11_port, B => ML_int_3_3_port, S 
                           => SH(3), Z => ML_int_4_11_port);
   M1_3_10 : MUX2_X1 port map( A => ML_int_3_10_port, B => ML_int_3_2_port, S 
                           => SH(3), Z => ML_int_4_10_port);
   M1_3_9 : MUX2_X1 port map( A => ML_int_3_9_port, B => ML_int_3_1_port, S => 
                           SH(3), Z => ML_int_4_9_port);
   M1_3_8 : MUX2_X1 port map( A => ML_int_3_8_port, B => ML_int_3_0_port, S => 
                           SH(3), Z => ML_int_4_8_port);
   M0_3_7 : MUX2_X1 port map( A => ML_int_3_7_port, B => ML_int_3_31_port, S =>
                           SH(3), Z => ML_int_4_7_port);
   M0_3_6 : MUX2_X1 port map( A => ML_int_3_6_port, B => ML_int_3_30_port, S =>
                           SH(3), Z => ML_int_4_6_port);
   M0_3_5 : MUX2_X1 port map( A => ML_int_3_5_port, B => ML_int_3_29_port, S =>
                           SH(3), Z => ML_int_4_5_port);
   M0_3_4 : MUX2_X1 port map( A => ML_int_3_4_port, B => ML_int_3_28_port, S =>
                           SH(3), Z => ML_int_4_4_port);
   M0_3_3 : MUX2_X1 port map( A => ML_int_3_3_port, B => ML_int_3_27_port, S =>
                           SH(3), Z => ML_int_4_3_port);
   M0_3_2 : MUX2_X1 port map( A => ML_int_3_2_port, B => ML_int_3_26_port, S =>
                           SH(3), Z => ML_int_4_2_port);
   M0_3_1 : MUX2_X1 port map( A => ML_int_3_1_port, B => ML_int_3_25_port, S =>
                           SH(3), Z => ML_int_4_1_port);
   M0_3_0 : MUX2_X1 port map( A => ML_int_3_0_port, B => ML_int_3_24_port, S =>
                           SH(3), Z => ML_int_4_0_port);
   M1_2_31 : MUX2_X1 port map( A => ML_int_2_31_port, B => ML_int_2_27_port, S 
                           => SH(2), Z => ML_int_3_31_port);
   M1_2_30 : MUX2_X1 port map( A => ML_int_2_30_port, B => ML_int_2_26_port, S 
                           => SH(2), Z => ML_int_3_30_port);
   M1_2_29 : MUX2_X1 port map( A => ML_int_2_29_port, B => ML_int_2_25_port, S 
                           => SH(2), Z => ML_int_3_29_port);
   M1_2_28 : MUX2_X1 port map( A => ML_int_2_28_port, B => ML_int_2_24_port, S 
                           => SH(2), Z => ML_int_3_28_port);
   M1_2_27 : MUX2_X1 port map( A => ML_int_2_27_port, B => ML_int_2_23_port, S 
                           => SH(2), Z => ML_int_3_27_port);
   M1_2_26 : MUX2_X1 port map( A => ML_int_2_26_port, B => ML_int_2_22_port, S 
                           => SH(2), Z => ML_int_3_26_port);
   M1_2_25 : MUX2_X1 port map( A => ML_int_2_25_port, B => ML_int_2_21_port, S 
                           => SH(2), Z => ML_int_3_25_port);
   M1_2_24 : MUX2_X1 port map( A => ML_int_2_24_port, B => ML_int_2_20_port, S 
                           => SH(2), Z => ML_int_3_24_port);
   M1_2_23 : MUX2_X1 port map( A => ML_int_2_23_port, B => ML_int_2_19_port, S 
                           => SH(2), Z => ML_int_3_23_port);
   M1_2_22 : MUX2_X1 port map( A => ML_int_2_22_port, B => ML_int_2_18_port, S 
                           => SH(2), Z => ML_int_3_22_port);
   M1_2_21 : MUX2_X1 port map( A => ML_int_2_21_port, B => ML_int_2_17_port, S 
                           => SH(2), Z => ML_int_3_21_port);
   M1_2_20 : MUX2_X1 port map( A => ML_int_2_20_port, B => ML_int_2_16_port, S 
                           => SH(2), Z => ML_int_3_20_port);
   M1_2_19 : MUX2_X1 port map( A => ML_int_2_19_port, B => ML_int_2_15_port, S 
                           => SH(2), Z => ML_int_3_19_port);
   M1_2_18 : MUX2_X1 port map( A => ML_int_2_18_port, B => ML_int_2_14_port, S 
                           => SH(2), Z => ML_int_3_18_port);
   M1_2_17 : MUX2_X1 port map( A => ML_int_2_17_port, B => ML_int_2_13_port, S 
                           => SH(2), Z => ML_int_3_17_port);
   M1_2_16 : MUX2_X1 port map( A => ML_int_2_16_port, B => ML_int_2_12_port, S 
                           => SH(2), Z => ML_int_3_16_port);
   M1_2_15 : MUX2_X1 port map( A => ML_int_2_15_port, B => ML_int_2_11_port, S 
                           => SH(2), Z => ML_int_3_15_port);
   M1_2_14 : MUX2_X1 port map( A => ML_int_2_14_port, B => ML_int_2_10_port, S 
                           => SH(2), Z => ML_int_3_14_port);
   M1_2_13 : MUX2_X1 port map( A => ML_int_2_13_port, B => ML_int_2_9_port, S 
                           => SH(2), Z => ML_int_3_13_port);
   M1_2_12 : MUX2_X1 port map( A => ML_int_2_12_port, B => ML_int_2_8_port, S 
                           => SH(2), Z => ML_int_3_12_port);
   M1_2_11 : MUX2_X1 port map( A => ML_int_2_11_port, B => ML_int_2_7_port, S 
                           => SH(2), Z => ML_int_3_11_port);
   M1_2_10 : MUX2_X1 port map( A => ML_int_2_10_port, B => ML_int_2_6_port, S 
                           => SH(2), Z => ML_int_3_10_port);
   M1_2_9 : MUX2_X1 port map( A => ML_int_2_9_port, B => ML_int_2_5_port, S => 
                           SH(2), Z => ML_int_3_9_port);
   M1_2_8 : MUX2_X1 port map( A => ML_int_2_8_port, B => ML_int_2_4_port, S => 
                           SH(2), Z => ML_int_3_8_port);
   M1_2_7 : MUX2_X1 port map( A => ML_int_2_7_port, B => ML_int_2_3_port, S => 
                           SH(2), Z => ML_int_3_7_port);
   M1_2_6 : MUX2_X1 port map( A => ML_int_2_6_port, B => ML_int_2_2_port, S => 
                           SH(2), Z => ML_int_3_6_port);
   M1_2_5 : MUX2_X1 port map( A => ML_int_2_5_port, B => ML_int_2_1_port, S => 
                           SH(2), Z => ML_int_3_5_port);
   M1_2_4 : MUX2_X1 port map( A => ML_int_2_4_port, B => ML_int_2_0_port, S => 
                           SH(2), Z => ML_int_3_4_port);
   M0_2_3 : MUX2_X1 port map( A => ML_int_2_3_port, B => ML_int_2_31_port, S =>
                           SH(2), Z => ML_int_3_3_port);
   M0_2_2 : MUX2_X1 port map( A => ML_int_2_2_port, B => ML_int_2_30_port, S =>
                           SH(2), Z => ML_int_3_2_port);
   M0_2_1 : MUX2_X1 port map( A => ML_int_2_1_port, B => ML_int_2_29_port, S =>
                           SH(2), Z => ML_int_3_1_port);
   M0_2_0 : MUX2_X1 port map( A => ML_int_2_0_port, B => ML_int_2_28_port, S =>
                           SH(2), Z => ML_int_3_0_port);
   M1_1_31 : MUX2_X1 port map( A => ML_int_1_31_port, B => ML_int_1_29_port, S 
                           => SH(1), Z => ML_int_2_31_port);
   M1_1_30 : MUX2_X1 port map( A => ML_int_1_30_port, B => ML_int_1_28_port, S 
                           => SH(1), Z => ML_int_2_30_port);
   M1_1_29 : MUX2_X1 port map( A => ML_int_1_29_port, B => ML_int_1_27_port, S 
                           => SH(1), Z => ML_int_2_29_port);
   M1_1_28 : MUX2_X1 port map( A => ML_int_1_28_port, B => ML_int_1_26_port, S 
                           => SH(1), Z => ML_int_2_28_port);
   M1_1_27 : MUX2_X1 port map( A => ML_int_1_27_port, B => ML_int_1_25_port, S 
                           => SH(1), Z => ML_int_2_27_port);
   M1_1_26 : MUX2_X1 port map( A => ML_int_1_26_port, B => ML_int_1_24_port, S 
                           => SH(1), Z => ML_int_2_26_port);
   M1_1_25 : MUX2_X1 port map( A => ML_int_1_25_port, B => ML_int_1_23_port, S 
                           => SH(1), Z => ML_int_2_25_port);
   M1_1_24 : MUX2_X1 port map( A => ML_int_1_24_port, B => ML_int_1_22_port, S 
                           => SH(1), Z => ML_int_2_24_port);
   M1_1_23 : MUX2_X1 port map( A => ML_int_1_23_port, B => ML_int_1_21_port, S 
                           => SH(1), Z => ML_int_2_23_port);
   M1_1_22 : MUX2_X1 port map( A => ML_int_1_22_port, B => ML_int_1_20_port, S 
                           => SH(1), Z => ML_int_2_22_port);
   M1_1_21 : MUX2_X1 port map( A => ML_int_1_21_port, B => ML_int_1_19_port, S 
                           => SH(1), Z => ML_int_2_21_port);
   M1_1_20 : MUX2_X1 port map( A => ML_int_1_20_port, B => ML_int_1_18_port, S 
                           => SH(1), Z => ML_int_2_20_port);
   M1_1_19 : MUX2_X1 port map( A => ML_int_1_19_port, B => ML_int_1_17_port, S 
                           => SH(1), Z => ML_int_2_19_port);
   M1_1_18 : MUX2_X1 port map( A => ML_int_1_18_port, B => ML_int_1_16_port, S 
                           => SH(1), Z => ML_int_2_18_port);
   M1_1_17 : MUX2_X1 port map( A => ML_int_1_17_port, B => ML_int_1_15_port, S 
                           => SH(1), Z => ML_int_2_17_port);
   M1_1_16 : MUX2_X1 port map( A => ML_int_1_16_port, B => ML_int_1_14_port, S 
                           => SH(1), Z => ML_int_2_16_port);
   M1_1_15 : MUX2_X1 port map( A => ML_int_1_15_port, B => ML_int_1_13_port, S 
                           => SH(1), Z => ML_int_2_15_port);
   M1_1_14 : MUX2_X1 port map( A => ML_int_1_14_port, B => ML_int_1_12_port, S 
                           => SH(1), Z => ML_int_2_14_port);
   M1_1_13 : MUX2_X1 port map( A => ML_int_1_13_port, B => ML_int_1_11_port, S 
                           => SH(1), Z => ML_int_2_13_port);
   M1_1_12 : MUX2_X1 port map( A => ML_int_1_12_port, B => ML_int_1_10_port, S 
                           => SH(1), Z => ML_int_2_12_port);
   M1_1_11 : MUX2_X1 port map( A => ML_int_1_11_port, B => ML_int_1_9_port, S 
                           => SH(1), Z => ML_int_2_11_port);
   M1_1_10 : MUX2_X1 port map( A => ML_int_1_10_port, B => ML_int_1_8_port, S 
                           => SH(1), Z => ML_int_2_10_port);
   M1_1_9 : MUX2_X1 port map( A => ML_int_1_9_port, B => ML_int_1_7_port, S => 
                           SH(1), Z => ML_int_2_9_port);
   M1_1_8 : MUX2_X1 port map( A => ML_int_1_8_port, B => ML_int_1_6_port, S => 
                           SH(1), Z => ML_int_2_8_port);
   M1_1_7 : MUX2_X1 port map( A => ML_int_1_7_port, B => ML_int_1_5_port, S => 
                           SH(1), Z => ML_int_2_7_port);
   M1_1_6 : MUX2_X1 port map( A => ML_int_1_6_port, B => ML_int_1_4_port, S => 
                           SH(1), Z => ML_int_2_6_port);
   M1_1_5 : MUX2_X1 port map( A => ML_int_1_5_port, B => ML_int_1_3_port, S => 
                           SH(1), Z => ML_int_2_5_port);
   M1_1_4 : MUX2_X1 port map( A => ML_int_1_4_port, B => ML_int_1_2_port, S => 
                           SH(1), Z => ML_int_2_4_port);
   M1_1_3 : MUX2_X1 port map( A => ML_int_1_3_port, B => ML_int_1_1_port, S => 
                           SH(1), Z => ML_int_2_3_port);
   M1_1_2 : MUX2_X1 port map( A => ML_int_1_2_port, B => ML_int_1_0_port, S => 
                           SH(1), Z => ML_int_2_2_port);
   M0_1_1 : MUX2_X1 port map( A => ML_int_1_1_port, B => ML_int_1_31_port, S =>
                           SH(1), Z => ML_int_2_1_port);
   M0_1_0 : MUX2_X1 port map( A => ML_int_1_0_port, B => ML_int_1_30_port, S =>
                           SH(1), Z => ML_int_2_0_port);
   M1_0_31 : MUX2_X1 port map( A => A(31), B => A(30), S => SH(0), Z => 
                           ML_int_1_31_port);
   M1_0_30 : MUX2_X1 port map( A => A(30), B => A(29), S => SH(0), Z => 
                           ML_int_1_30_port);
   M1_0_29 : MUX2_X1 port map( A => A(29), B => A(28), S => SH(0), Z => 
                           ML_int_1_29_port);
   M1_0_28 : MUX2_X1 port map( A => A(28), B => A(27), S => SH(0), Z => 
                           ML_int_1_28_port);
   M1_0_27 : MUX2_X1 port map( A => A(27), B => A(26), S => SH(0), Z => 
                           ML_int_1_27_port);
   M1_0_26 : MUX2_X1 port map( A => A(26), B => A(25), S => SH(0), Z => 
                           ML_int_1_26_port);
   M1_0_25 : MUX2_X1 port map( A => A(25), B => A(24), S => SH(0), Z => 
                           ML_int_1_25_port);
   M1_0_24 : MUX2_X1 port map( A => A(24), B => A(23), S => SH(0), Z => 
                           ML_int_1_24_port);
   M1_0_23 : MUX2_X1 port map( A => A(23), B => A(22), S => SH(0), Z => 
                           ML_int_1_23_port);
   M1_0_22 : MUX2_X1 port map( A => A(22), B => A(21), S => SH(0), Z => 
                           ML_int_1_22_port);
   M1_0_21 : MUX2_X1 port map( A => A(21), B => A(20), S => SH(0), Z => 
                           ML_int_1_21_port);
   M1_0_20 : MUX2_X1 port map( A => A(20), B => A(19), S => SH(0), Z => 
                           ML_int_1_20_port);
   M1_0_19 : MUX2_X1 port map( A => A(19), B => A(18), S => SH(0), Z => 
                           ML_int_1_19_port);
   M1_0_18 : MUX2_X1 port map( A => A(18), B => A(17), S => SH(0), Z => 
                           ML_int_1_18_port);
   M1_0_17 : MUX2_X1 port map( A => A(17), B => A(16), S => SH(0), Z => 
                           ML_int_1_17_port);
   M1_0_16 : MUX2_X1 port map( A => A(16), B => A(15), S => SH(0), Z => 
                           ML_int_1_16_port);
   M1_0_15 : MUX2_X1 port map( A => A(15), B => A(14), S => SH(0), Z => 
                           ML_int_1_15_port);
   M1_0_14 : MUX2_X1 port map( A => A(14), B => A(13), S => SH(0), Z => 
                           ML_int_1_14_port);
   M1_0_13 : MUX2_X1 port map( A => A(13), B => A(12), S => SH(0), Z => 
                           ML_int_1_13_port);
   M1_0_12 : MUX2_X1 port map( A => A(12), B => A(11), S => SH(0), Z => 
                           ML_int_1_12_port);
   M1_0_11 : MUX2_X1 port map( A => A(11), B => A(10), S => SH(0), Z => 
                           ML_int_1_11_port);
   M1_0_10 : MUX2_X1 port map( A => A(10), B => A(9), S => SH(0), Z => 
                           ML_int_1_10_port);
   M1_0_9 : MUX2_X1 port map( A => A(9), B => A(8), S => SH(0), Z => 
                           ML_int_1_9_port);
   M1_0_8 : MUX2_X1 port map( A => A(8), B => A(7), S => SH(0), Z => 
                           ML_int_1_8_port);
   M1_0_7 : MUX2_X1 port map( A => A(7), B => A(6), S => SH(0), Z => 
                           ML_int_1_7_port);
   M1_0_6 : MUX2_X1 port map( A => A(6), B => A(5), S => SH(0), Z => 
                           ML_int_1_6_port);
   M1_0_5 : MUX2_X1 port map( A => A(5), B => A(4), S => SH(0), Z => 
                           ML_int_1_5_port);
   M1_0_4 : MUX2_X1 port map( A => A(4), B => A(3), S => SH(0), Z => 
                           ML_int_1_4_port);
   M1_0_3 : MUX2_X1 port map( A => A(3), B => A(2), S => SH(0), Z => 
                           ML_int_1_3_port);
   M1_0_2 : MUX2_X1 port map( A => A(2), B => A(1), S => SH(0), Z => 
                           ML_int_1_2_port);
   M1_0_1 : MUX2_X1 port map( A => A(1), B => A(0), S => SH(0), Z => 
                           ML_int_1_1_port);
   M0_0_0 : MUX2_X1 port map( A => A(0), B => A(31), S => SH(0), Z => 
                           ML_int_1_0_port);
   U2 : BUF_X1 port map( A => SH(4), Z => n1);
   U3 : BUF_X1 port map( A => SH(4), Z => n2);
   U4 : BUF_X1 port map( A => SH(4), Z => n3);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Shifter_DATA_SIZE32_DW_sra_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end Shifter_DATA_SIZE32_DW_sra_0;

architecture SYN_mx2 of Shifter_DATA_SIZE32_DW_sra_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, B_25_port, 
      B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, B_19_port, 
      B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, B_13_port, 
      B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port, B_6_port, 
      B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, B_0_port, n1, n2, n3, 
      n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171 : std_logic;

begin
   B <= ( A(31), B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, 
      B_25_port, B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, 
      B_19_port, B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, 
      B_13_port, B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port,
      B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, B_0_port );
   
   U2 : NOR2_X2 port map( A1 => SH(2), A2 => SH(3), ZN => n73);
   U3 : INV_X1 port map( A => SH(4), ZN => n1);
   U4 : OAI221_X1 port map( B1 => n2, B2 => n3, C1 => n4, C2 => n1, A => n5, ZN
                           => B_9_port);
   U5 : AOI222_X1 port map( A1 => n6, A2 => n7, B1 => n8, B2 => n9, C1 => n10, 
                           C2 => n11, ZN => n5);
   U6 : INV_X1 port map( A => n12, ZN => n2);
   U7 : OAI221_X1 port map( B1 => n13, B2 => n3, C1 => n14, C2 => n1, A => n15,
                           ZN => B_8_port);
   U8 : AOI222_X1 port map( A1 => n6, A2 => n16, B1 => n8, B2 => n17, C1 => n10
                           , C2 => n18, ZN => n15);
   U9 : INV_X1 port map( A => n19, ZN => n13);
   U10 : OAI221_X1 port map( B1 => n20, B2 => n3, C1 => n21, C2 => n1, A => n22
                           , ZN => B_7_port);
   U11 : AOI222_X1 port map( A1 => n6, A2 => n23, B1 => n8, B2 => n24, C1 => 
                           n10, C2 => n25, ZN => n22);
   U12 : OAI221_X1 port map( B1 => n26, B2 => n3, C1 => n27, C2 => n1, A => n28
                           , ZN => B_6_port);
   U13 : AOI222_X1 port map( A1 => n6, A2 => n29, B1 => n8, B2 => n30, C1 => 
                           n10, C2 => n31, ZN => n28);
   U14 : OAI221_X1 port map( B1 => n32, B2 => n3, C1 => n33, C2 => n1, A => n34
                           , ZN => B_5_port);
   U15 : AOI222_X1 port map( A1 => n6, A2 => n12, B1 => n8, B2 => n7, C1 => n10
                           , C2 => n9, ZN => n34);
   U16 : OAI221_X1 port map( B1 => n35, B2 => n3, C1 => n36, C2 => n1, A => n37
                           , ZN => B_4_port);
   U17 : AOI222_X1 port map( A1 => n6, A2 => n19, B1 => n8, B2 => n16, C1 => 
                           n10, C2 => n17, ZN => n37);
   U18 : OAI221_X1 port map( B1 => n20, B2 => n38, C1 => n39, C2 => n1, A => 
                           n40, ZN => B_3_port);
   U19 : AOI222_X1 port map( A1 => n10, A2 => n24, B1 => n41, B2 => n42, C1 => 
                           n8, C2 => n23, ZN => n40);
   U20 : OAI221_X1 port map( B1 => n43, B2 => n44, C1 => n45, C2 => n46, A => 
                           n47, ZN => n42);
   U21 : AOI22_X1 port map( A1 => A(5), A2 => n48, B1 => A(6), B2 => n49, ZN =>
                           n47);
   U22 : INV_X1 port map( A => A(4), ZN => n44);
   U23 : AOI221_X1 port map( B1 => n50, B2 => A(8), C1 => n51, C2 => A(7), A =>
                           n52, ZN => n20);
   U24 : OAI22_X1 port map( A1 => n53, A2 => n54, B1 => n55, B2 => n56, ZN => 
                           n52);
   U25 : OAI21_X1 port map( B1 => SH(4), B2 => n57, A => n58, ZN => B_30_port);
   U26 : OAI221_X1 port map( B1 => n26, B2 => n38, C1 => n59, C2 => n1, A => 
                           n60, ZN => B_2_port);
   U27 : AOI222_X1 port map( A1 => n10, A2 => n30, B1 => n41, B2 => n61, C1 => 
                           n8, C2 => n29, ZN => n60);
   U28 : OAI221_X1 port map( B1 => n43, B2 => n46, C1 => n45, C2 => n62, A => 
                           n63, ZN => n61);
   U29 : AOI22_X1 port map( A1 => A(4), A2 => n48, B1 => A(5), B2 => n49, ZN =>
                           n63);
   U30 : AOI221_X1 port map( B1 => n50, B2 => A(7), C1 => n51, C2 => A(6), A =>
                           n64, ZN => n26);
   U31 : OAI22_X1 port map( A1 => n65, A2 => n54, B1 => n53, B2 => n56, ZN => 
                           n64);
   U32 : OAI21_X1 port map( B1 => SH(4), B2 => n66, A => n58, ZN => B_29_port);
   U33 : OAI21_X1 port map( B1 => SH(4), B2 => n67, A => n58, ZN => B_28_port);
   U34 : OAI21_X1 port map( B1 => SH(4), B2 => n68, A => n58, ZN => B_27_port);
   U35 : OAI21_X1 port map( B1 => SH(4), B2 => n69, A => n58, ZN => B_26_port);
   U36 : OAI21_X1 port map( B1 => SH(4), B2 => n4, A => n58, ZN => B_25_port);
   U37 : AOI221_X1 port map( B1 => n70, B2 => n71, C1 => n72, C2 => n73, A => 
                           n74, ZN => n4);
   U38 : OAI21_X1 port map( B1 => SH(4), B2 => n14, A => n58, ZN => B_24_port);
   U39 : AOI221_X1 port map( B1 => n75, B2 => n71, C1 => n76, C2 => n73, A => 
                           n74, ZN => n14);
   U40 : OAI21_X1 port map( B1 => SH(4), B2 => n21, A => n58, ZN => B_23_port);
   U41 : AOI221_X1 port map( B1 => n77, B2 => n71, C1 => n78, C2 => n73, A => 
                           n74, ZN => n21);
   U42 : OAI21_X1 port map( B1 => SH(4), B2 => n27, A => n58, ZN => B_22_port);
   U43 : AOI221_X1 port map( B1 => n79, B2 => n71, C1 => n80, C2 => n73, A => 
                           n81, ZN => n27);
   U44 : INV_X1 port map( A => n82, ZN => n81);
   U45 : AOI21_X1 port map( B1 => n83, B2 => n84, A => n85, ZN => n82);
   U46 : OAI21_X1 port map( B1 => SH(4), B2 => n33, A => n58, ZN => B_21_port);
   U47 : AOI221_X1 port map( B1 => n72, B2 => n71, C1 => n11, C2 => n73, A => 
                           n86, ZN => n33);
   U48 : INV_X1 port map( A => n87, ZN => n86);
   U49 : AOI21_X1 port map( B1 => n83, B2 => n70, A => n85, ZN => n87);
   U50 : OAI21_X1 port map( B1 => SH(4), B2 => n36, A => n58, ZN => B_20_port);
   U51 : AOI221_X1 port map( B1 => n76, B2 => n71, C1 => n18, C2 => n73, A => 
                           n88, ZN => n36);
   U52 : INV_X1 port map( A => n89, ZN => n88);
   U53 : AOI21_X1 port map( B1 => n83, B2 => n75, A => n85, ZN => n89);
   U54 : OAI221_X1 port map( B1 => n32, B2 => n38, C1 => n90, C2 => n1, A => 
                           n91, ZN => B_1_port);
   U55 : AOI222_X1 port map( A1 => n10, A2 => n7, B1 => n41, B2 => n92, C1 => 
                           n8, C2 => n12, ZN => n91);
   U56 : OAI221_X1 port map( B1 => n43, B2 => n55, C1 => n45, C2 => n53, A => 
                           n93, ZN => n12);
   U57 : AOI22_X1 port map( A1 => A(11), A2 => n48, B1 => A(12), B2 => n49, ZN 
                           => n93);
   U58 : OAI221_X1 port map( B1 => n43, B2 => n62, C1 => n45, C2 => n94, A => 
                           n95, ZN => n92);
   U59 : AOI22_X1 port map( A1 => A(3), A2 => n48, B1 => A(4), B2 => n49, ZN =>
                           n95);
   U60 : INV_X1 port map( A => A(1), ZN => n94);
   U61 : AOI221_X1 port map( B1 => n50, B2 => A(6), C1 => n51, C2 => A(5), A =>
                           n96, ZN => n32);
   U62 : OAI22_X1 port map( A1 => n97, A2 => n54, B1 => n65, B2 => n56, ZN => 
                           n96);
   U63 : OAI21_X1 port map( B1 => SH(4), B2 => n39, A => n58, ZN => B_19_port);
   U64 : AOI221_X1 port map( B1 => n78, B2 => n71, C1 => n25, C2 => n73, A => 
                           n98, ZN => n39);
   U65 : INV_X1 port map( A => n99, ZN => n98);
   U66 : AOI21_X1 port map( B1 => n83, B2 => n77, A => n85, ZN => n99);
   U67 : NOR2_X1 port map( A1 => n100, A2 => n101, ZN => n85);
   U68 : OAI21_X1 port map( B1 => SH(4), B2 => n59, A => n58, ZN => B_18_port);
   U69 : AOI221_X1 port map( B1 => n80, B2 => n71, C1 => n31, C2 => n73, A => 
                           n102, ZN => n59);
   U70 : INV_X1 port map( A => n103, ZN => n102);
   U71 : AOI22_X1 port map( A1 => n104, A2 => n84, B1 => n83, B2 => n79, ZN => 
                           n103);
   U72 : OAI21_X1 port map( B1 => SH(4), B2 => n90, A => n58, ZN => B_17_port);
   U73 : AOI221_X1 port map( B1 => n11, B2 => n71, C1 => n9, C2 => n73, A => 
                           n105, ZN => n90);
   U74 : INV_X1 port map( A => n106, ZN => n105);
   U75 : AOI22_X1 port map( A1 => n104, A2 => n70, B1 => n83, B2 => n72, ZN => 
                           n106);
   U76 : OAI21_X1 port map( B1 => SH(4), B2 => n107, A => n58, ZN => B_16_port)
                           ;
   U77 : OAI221_X1 port map( B1 => n108, B2 => n38, C1 => n109, C2 => n3, A => 
                           n110, ZN => B_15_port);
   U78 : AOI221_X1 port map( B1 => n10, B2 => n77, C1 => n8, C2 => n78, A => 
                           n111, ZN => n110);
   U79 : INV_X1 port map( A => n58, ZN => n111);
   U80 : NAND2_X1 port map( A1 => SH(4), A2 => A(31), ZN => n58);
   U81 : INV_X1 port map( A => n25, ZN => n108);
   U82 : OAI221_X1 port map( B1 => n112, B2 => n3, C1 => n57, C2 => n1, A => 
                           n113, ZN => B_14_port);
   U83 : AOI222_X1 port map( A1 => n6, A2 => n31, B1 => n8, B2 => n80, C1 => 
                           n10, C2 => n79, ZN => n113);
   U84 : AOI21_X1 port map( B1 => n84, B2 => n73, A => n114, ZN => n57);
   U85 : OAI221_X1 port map( B1 => n115, B2 => n3, C1 => n66, C2 => n1, A => 
                           n116, ZN => B_13_port);
   U86 : AOI222_X1 port map( A1 => n6, A2 => n9, B1 => n8, B2 => n11, C1 => n10
                           , C2 => n72, ZN => n116);
   U87 : OAI221_X1 port map( B1 => n43, B2 => n117, C1 => n45, C2 => n118, A =>
                           n119, ZN => n72);
   U88 : AOI22_X1 port map( A1 => A(27), A2 => n48, B1 => A(28), B2 => n49, ZN 
                           => n119);
   U89 : OAI221_X1 port map( B1 => n43, B2 => n120, C1 => n45, C2 => n121, A =>
                           n122, ZN => n11);
   U90 : AOI22_X1 port map( A1 => A(23), A2 => n48, B1 => A(24), B2 => n49, ZN 
                           => n122);
   U91 : OAI221_X1 port map( B1 => n43, B2 => n123, C1 => n45, C2 => n124, A =>
                           n125, ZN => n9);
   U92 : AOI22_X1 port map( A1 => A(19), A2 => n48, B1 => A(20), B2 => n49, ZN 
                           => n125);
   U93 : AOI21_X1 port map( B1 => n70, B2 => n73, A => n114, ZN => n66);
   U94 : INV_X1 port map( A => n126, ZN => n70);
   U95 : AOI222_X1 port map( A1 => n51, A2 => A(29), B1 => n50, B2 => A(30), C1
                           => SH(1), C2 => A(31), ZN => n126);
   U96 : INV_X1 port map( A => n7, ZN => n115);
   U97 : OAI221_X1 port map( B1 => n43, B2 => n127, C1 => n45, C2 => n128, A =>
                           n129, ZN => n7);
   U98 : AOI22_X1 port map( A1 => A(15), A2 => n48, B1 => A(16), B2 => n49, ZN 
                           => n129);
   U99 : INV_X1 port map( A => A(14), ZN => n127);
   U100 : OAI221_X1 port map( B1 => n130, B2 => n3, C1 => n67, C2 => n1, A => 
                           n131, ZN => B_12_port);
   U101 : AOI222_X1 port map( A1 => n6, A2 => n17, B1 => n8, B2 => n18, C1 => 
                           n10, C2 => n76, ZN => n131);
   U102 : AOI21_X1 port map( B1 => n75, B2 => n73, A => n114, ZN => n67);
   U103 : INV_X1 port map( A => n16, ZN => n130);
   U104 : OAI221_X1 port map( B1 => n132, B2 => n3, C1 => n68, C2 => n1, A => 
                           n133, ZN => B_11_port);
   U105 : AOI222_X1 port map( A1 => n6, A2 => n24, B1 => n8, B2 => n25, C1 => 
                           n10, C2 => n78, ZN => n133);
   U106 : OAI221_X1 port map( B1 => n43, B2 => n134, C1 => n45, C2 => n135, A 
                           => n136, ZN => n78);
   U107 : AOI22_X1 port map( A1 => A(25), A2 => n48, B1 => A(26), B2 => n49, ZN
                           => n136);
   U108 : OAI221_X1 port map( B1 => n137, B2 => n43, C1 => n138, C2 => n45, A 
                           => n139, ZN => n25);
   U109 : AOI22_X1 port map( A1 => A(21), A2 => n48, B1 => A(22), B2 => n49, ZN
                           => n139);
   U110 : INV_X1 port map( A => n109, ZN => n24);
   U111 : AOI221_X1 port map( B1 => n50, B2 => A(16), C1 => n51, C2 => A(15), A
                           => n140, ZN => n109);
   U112 : OAI22_X1 port map( A1 => n124, A2 => n54, B1 => n123, B2 => n56, ZN 
                           => n140);
   U113 : INV_X1 port map( A => A(17), ZN => n124);
   U114 : AOI21_X1 port map( B1 => n77, B2 => n73, A => n114, ZN => n68);
   U115 : OAI21_X1 port map( B1 => n101, B2 => n141, A => n100, ZN => n114);
   U116 : INV_X1 port map( A => A(31), ZN => n141);
   U117 : OAI221_X1 port map( B1 => n43, B2 => n142, C1 => n45, C2 => n143, A 
                           => n144, ZN => n77);
   U118 : AOI22_X1 port map( A1 => A(29), A2 => n48, B1 => A(30), B2 => n49, ZN
                           => n144);
   U119 : INV_X1 port map( A => n23, ZN => n132);
   U120 : OAI221_X1 port map( B1 => n43, B2 => n145, C1 => n45, C2 => n146, A 
                           => n147, ZN => n23);
   U121 : AOI22_X1 port map( A1 => A(13), A2 => n48, B1 => A(14), B2 => n49, ZN
                           => n147);
   U122 : OAI221_X1 port map( B1 => n148, B2 => n3, C1 => n69, C2 => n1, A => 
                           n149, ZN => B_10_port);
   U123 : AOI222_X1 port map( A1 => n6, A2 => n30, B1 => n8, B2 => n31, C1 => 
                           n10, C2 => n80, ZN => n149);
   U124 : OAI221_X1 port map( B1 => n43, B2 => n135, C1 => n45, C2 => n120, A 
                           => n150, ZN => n80);
   U125 : AOI22_X1 port map( A1 => A(24), A2 => n48, B1 => A(25), B2 => n49, ZN
                           => n150);
   U126 : INV_X1 port map( A => A(22), ZN => n120);
   U127 : INV_X1 port map( A => A(23), ZN => n135);
   U128 : OAI221_X1 port map( B1 => n138, B2 => n43, C1 => n123, C2 => n45, A 
                           => n151, ZN => n31);
   U129 : AOI22_X1 port map( A1 => A(20), A2 => n48, B1 => A(21), B2 => n49, ZN
                           => n151);
   U130 : INV_X1 port map( A => n112, ZN => n30);
   U131 : AOI221_X1 port map( B1 => n50, B2 => A(15), C1 => n51, C2 => A(14), A
                           => n152, ZN => n112);
   U132 : INV_X1 port map( A => n153, ZN => n152);
   U133 : AOI22_X1 port map( A1 => A(16), A2 => n48, B1 => A(17), B2 => n49, ZN
                           => n153);
   U134 : INV_X1 port map( A => n38, ZN => n6);
   U135 : AOI221_X1 port map( B1 => n84, B2 => n71, C1 => n79, C2 => n73, A => 
                           n74, ZN => n69);
   U136 : INV_X1 port map( A => n100, ZN => n74);
   U137 : NAND2_X1 port map( A1 => A(31), A2 => SH(3), ZN => n100);
   U138 : OAI221_X1 port map( B1 => n43, B2 => n143, C1 => n45, C2 => n117, A 
                           => n154, ZN => n79);
   U139 : AOI22_X1 port map( A1 => A(28), A2 => n48, B1 => A(29), B2 => n49, ZN
                           => n154);
   U140 : INV_X1 port map( A => A(26), ZN => n117);
   U141 : INV_X1 port map( A => A(27), ZN => n143);
   U142 : MUX2_X1 port map( A => A(31), B => A(30), S => n51, Z => n84);
   U143 : INV_X1 port map( A => n29, ZN => n148);
   U144 : OAI221_X1 port map( B1 => n43, B2 => n146, C1 => n45, C2 => n55, A =>
                           n155, ZN => n29);
   U145 : AOI22_X1 port map( A1 => A(12), A2 => n48, B1 => A(13), B2 => n49, ZN
                           => n155);
   U146 : INV_X1 port map( A => A(10), ZN => n55);
   U147 : INV_X1 port map( A => A(11), ZN => n146);
   U148 : OAI221_X1 port map( B1 => n35, B2 => n38, C1 => n107, C2 => n1, A => 
                           n156, ZN => B_0_port);
   U149 : AOI222_X1 port map( A1 => n10, A2 => n16, B1 => n41, B2 => n157, C1 
                           => n8, C2 => n19, ZN => n156);
   U150 : OAI221_X1 port map( B1 => n43, B2 => n53, C1 => n45, C2 => n65, A => 
                           n158, ZN => n19);
   U151 : AOI22_X1 port map( A1 => A(10), A2 => n48, B1 => A(11), B2 => n49, ZN
                           => n158);
   U152 : INV_X1 port map( A => A(8), ZN => n65);
   U153 : INV_X1 port map( A => A(9), ZN => n53);
   U154 : AND2_X1 port map( A1 => n159, A2 => n101, ZN => n8);
   U155 : OAI221_X1 port map( B1 => n54, B2 => n62, C1 => n56, C2 => n46, A => 
                           n160, ZN => n157);
   U156 : AOI22_X1 port map( A1 => A(1), A2 => n50, B1 => A(0), B2 => n51, ZN 
                           => n160);
   U157 : INV_X1 port map( A => A(3), ZN => n46);
   U158 : INV_X1 port map( A => A(2), ZN => n62);
   U159 : INV_X1 port map( A => n3, ZN => n41);
   U160 : NAND2_X1 port map( A1 => n73, A2 => n1, ZN => n3);
   U161 : OAI221_X1 port map( B1 => n43, B2 => n128, C1 => n45, C2 => n145, A 
                           => n161, ZN => n16);
   U162 : AOI22_X1 port map( A1 => A(14), A2 => n48, B1 => A(15), B2 => n49, ZN
                           => n161);
   U163 : INV_X1 port map( A => A(12), ZN => n145);
   U164 : INV_X1 port map( A => A(13), ZN => n128);
   U165 : AND2_X1 port map( A1 => SH(2), A2 => n159, ZN => n10);
   U166 : AND2_X1 port map( A1 => SH(3), A2 => n1, ZN => n159);
   U167 : AOI221_X1 port map( B1 => n18, B2 => n71, C1 => n17, C2 => n73, A => 
                           n162, ZN => n107);
   U168 : INV_X1 port map( A => n163, ZN => n162);
   U169 : AOI22_X1 port map( A1 => n104, A2 => n75, B1 => n83, B2 => n76, ZN =>
                           n163);
   U170 : OAI221_X1 port map( B1 => n43, B2 => n118, C1 => n45, C2 => n134, A 
                           => n164, ZN => n76);
   U171 : AOI22_X1 port map( A1 => A(26), A2 => n48, B1 => A(27), B2 => n49, ZN
                           => n164);
   U172 : INV_X1 port map( A => A(24), ZN => n134);
   U173 : INV_X1 port map( A => A(25), ZN => n118);
   U174 : AND2_X1 port map( A1 => SH(3), A2 => n101, ZN => n83);
   U175 : OAI221_X1 port map( B1 => n43, B2 => n165, C1 => n45, C2 => n142, A 
                           => n166, ZN => n75);
   U176 : AOI22_X1 port map( A1 => A(30), A2 => n48, B1 => A(31), B2 => n49, ZN
                           => n166);
   U177 : INV_X1 port map( A => A(28), ZN => n142);
   U178 : INV_X1 port map( A => A(29), ZN => n165);
   U179 : AND2_X1 port map( A1 => SH(2), A2 => SH(3), ZN => n104);
   U180 : OAI221_X1 port map( B1 => n54, B2 => n123, C1 => n138, C2 => n56, A 
                           => n167, ZN => n17);
   U181 : AOI22_X1 port map( A1 => A(17), A2 => n50, B1 => A(16), B2 => n51, ZN
                           => n167);
   U182 : INV_X1 port map( A => A(19), ZN => n138);
   U183 : INV_X1 port map( A => A(18), ZN => n123);
   U184 : OAI221_X1 port map( B1 => n43, B2 => n121, C1 => n137, C2 => n45, A 
                           => n168, ZN => n18);
   U185 : AOI22_X1 port map( A1 => A(22), A2 => n48, B1 => A(23), B2 => n49, ZN
                           => n168);
   U186 : INV_X1 port map( A => n56, ZN => n49);
   U187 : INV_X1 port map( A => n54, ZN => n48);
   U188 : INV_X1 port map( A => n51, ZN => n45);
   U189 : INV_X1 port map( A => A(20), ZN => n137);
   U190 : INV_X1 port map( A => A(21), ZN => n121);
   U191 : INV_X1 port map( A => n50, ZN => n43);
   U192 : NAND2_X1 port map( A1 => n71, A2 => n1, ZN => n38);
   U193 : NOR2_X1 port map( A1 => n101, A2 => SH(3), ZN => n71);
   U194 : INV_X1 port map( A => SH(2), ZN => n101);
   U195 : AOI221_X1 port map( B1 => n50, B2 => A(5), C1 => n51, C2 => A(4), A 
                           => n169, ZN => n35);
   U196 : OAI22_X1 port map( A1 => n170, A2 => n54, B1 => n97, B2 => n56, ZN =>
                           n169);
   U197 : NAND2_X1 port map( A1 => SH(0), A2 => SH(1), ZN => n56);
   U198 : INV_X1 port map( A => A(7), ZN => n97);
   U199 : NAND2_X1 port map( A1 => SH(1), A2 => n171, ZN => n54);
   U200 : INV_X1 port map( A => A(6), ZN => n170);
   U201 : NOR2_X1 port map( A1 => SH(0), A2 => SH(1), ZN => n51);
   U202 : NOR2_X1 port map( A1 => n171, A2 => SH(1), ZN => n50);
   U203 : INV_X1 port map( A => SH(0), ZN => n171);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Shifter_DATA_SIZE32_DW_rash_0 is

   port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH : 
         in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out 
         std_logic_vector (31 downto 0));

end Shifter_DATA_SIZE32_DW_rash_0;

architecture SYN_mx2 of Shifter_DATA_SIZE32_DW_rash_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162 : 
      std_logic;

begin
   
   U3 : NOR2_X2 port map( A1 => SH(0), A2 => SH(1), ZN => n50);
   U4 : NOR2_X2 port map( A1 => n162, A2 => SH(1), ZN => n49);
   U5 : INV_X1 port map( A => SH(4), ZN => n1);
   U6 : OAI221_X1 port map( B1 => n2, B2 => n3, C1 => n4, C2 => n1, A => n5, ZN
                           => B(9));
   U7 : AOI222_X1 port map( A1 => n6, A2 => n7, B1 => n8, B2 => n9, C1 => n10, 
                           C2 => n11, ZN => n5);
   U8 : OAI221_X1 port map( B1 => n12, B2 => n3, C1 => n13, C2 => n1, A => n14,
                           ZN => B(8));
   U9 : AOI222_X1 port map( A1 => n6, A2 => n15, B1 => n8, B2 => n16, C1 => n10
                           , C2 => n17, ZN => n14);
   U10 : OAI221_X1 port map( B1 => n18, B2 => n3, C1 => n19, C2 => n1, A => n20
                           , ZN => B(7));
   U11 : AOI222_X1 port map( A1 => n6, A2 => n21, B1 => n8, B2 => n22, C1 => 
                           n10, C2 => n23, ZN => n20);
   U12 : OAI221_X1 port map( B1 => n24, B2 => n3, C1 => n25, C2 => n1, A => n26
                           , ZN => B(6));
   U13 : AOI222_X1 port map( A1 => n6, A2 => n27, B1 => n8, B2 => n28, C1 => 
                           n10, C2 => n29, ZN => n26);
   U14 : OAI221_X1 port map( B1 => n30, B2 => n3, C1 => n31, C2 => n1, A => n32
                           , ZN => B(5));
   U15 : AOI222_X1 port map( A1 => n6, A2 => n33, B1 => n8, B2 => n7, C1 => n10
                           , C2 => n9, ZN => n32);
   U16 : OAI221_X1 port map( B1 => n34, B2 => n3, C1 => n35, C2 => n1, A => n36
                           , ZN => B(4));
   U17 : AOI222_X1 port map( A1 => n6, A2 => n37, B1 => n8, B2 => n15, C1 => 
                           n10, C2 => n16, ZN => n36);
   U18 : OAI221_X1 port map( B1 => n18, B2 => n38, C1 => n39, C2 => n1, A => 
                           n40, ZN => B(3));
   U19 : AOI222_X1 port map( A1 => n10, A2 => n22, B1 => n41, B2 => n42, C1 => 
                           n8, C2 => n21, ZN => n40);
   U20 : INV_X1 port map( A => n43, ZN => n21);
   U21 : OAI221_X1 port map( B1 => n44, B2 => n45, C1 => n46, C2 => n47, A => 
                           n48, ZN => n42);
   U22 : AOI22_X1 port map( A1 => A(4), A2 => n49, B1 => A(3), B2 => n50, ZN =>
                           n48);
   U23 : AOI221_X1 port map( B1 => n51, B2 => A(10), C1 => n52, C2 => A(9), A 
                           => n53, ZN => n18);
   U24 : OAI22_X1 port map( A1 => n54, A2 => n55, B1 => n56, B2 => n57, ZN => 
                           n53);
   U25 : AND2_X1 port map( A1 => n41, A2 => n58, ZN => B(31));
   U26 : AND2_X1 port map( A1 => n59, A2 => n41, ZN => B(30));
   U27 : OAI221_X1 port map( B1 => n24, B2 => n38, C1 => n60, C2 => n1, A => 
                           n61, ZN => B(2));
   U28 : AOI222_X1 port map( A1 => n10, A2 => n28, B1 => n41, B2 => n62, C1 => 
                           n8, C2 => n27, ZN => n61);
   U29 : INV_X1 port map( A => n63, ZN => n27);
   U30 : OAI221_X1 port map( B1 => n44, B2 => n47, C1 => n46, C2 => n64, A => 
                           n65, ZN => n62);
   U31 : AOI22_X1 port map( A1 => A(3), A2 => n49, B1 => A(2), B2 => n50, ZN =>
                           n65);
   U32 : AOI221_X1 port map( B1 => n51, B2 => A(9), C1 => n52, C2 => A(8), A =>
                           n66, ZN => n24);
   U33 : OAI22_X1 port map( A1 => n56, A2 => n55, B1 => n45, B2 => n57, ZN => 
                           n66);
   U34 : INV_X1 port map( A => A(7), ZN => n56);
   U35 : AND2_X1 port map( A1 => n67, A2 => n41, ZN => B(29));
   U36 : AND2_X1 port map( A1 => n68, A2 => n41, ZN => B(28));
   U37 : NOR3_X1 port map( A1 => n69, A2 => SH(4), A3 => SH(3), ZN => B(27));
   U38 : NOR2_X1 port map( A1 => SH(4), A2 => n70, ZN => B(26));
   U39 : NOR2_X1 port map( A1 => SH(4), A2 => n4, ZN => B(25));
   U40 : AOI22_X1 port map( A1 => n71, A2 => n72, B1 => n67, B2 => n73, ZN => 
                           n4);
   U41 : NOR2_X1 port map( A1 => SH(4), A2 => n13, ZN => B(24));
   U42 : AOI22_X1 port map( A1 => n74, A2 => n72, B1 => n68, B2 => n73, ZN => 
                           n13);
   U43 : NOR2_X1 port map( A1 => SH(4), A2 => n19, ZN => B(23));
   U44 : AOI222_X1 port map( A1 => n75, A2 => n73, B1 => n58, B2 => n76, C1 => 
                           n77, C2 => n72, ZN => n19);
   U45 : NOR2_X1 port map( A1 => SH(4), A2 => n25, ZN => B(22));
   U46 : AOI222_X1 port map( A1 => n78, A2 => n73, B1 => n59, B2 => n76, C1 => 
                           n79, C2 => n72, ZN => n25);
   U47 : NOR2_X1 port map( A1 => SH(4), A2 => n31, ZN => B(21));
   U48 : AOI222_X1 port map( A1 => n71, A2 => n73, B1 => n67, B2 => n76, C1 => 
                           n11, C2 => n72, ZN => n31);
   U49 : NOR2_X1 port map( A1 => SH(4), A2 => n35, ZN => B(20));
   U50 : AOI222_X1 port map( A1 => n74, A2 => n73, B1 => n68, B2 => n76, C1 => 
                           n17, C2 => n72, ZN => n35);
   U51 : OAI221_X1 port map( B1 => n30, B2 => n38, C1 => n80, C2 => n1, A => 
                           n81, ZN => B(1));
   U52 : AOI222_X1 port map( A1 => n10, A2 => n7, B1 => n41, B2 => n82, C1 => 
                           n8, C2 => n33, ZN => n81);
   U53 : INV_X1 port map( A => n2, ZN => n33);
   U54 : AOI221_X1 port map( B1 => n51, B2 => A(12), C1 => n52, C2 => A(11), A 
                           => n83, ZN => n2);
   U55 : OAI22_X1 port map( A1 => n84, A2 => n55, B1 => n85, B2 => n57, ZN => 
                           n83);
   U56 : OAI221_X1 port map( B1 => n44, B2 => n64, C1 => n46, C2 => n86, A => 
                           n87, ZN => n82);
   U57 : AOI22_X1 port map( A1 => A(2), A2 => n49, B1 => A(1), B2 => n50, ZN =>
                           n87);
   U58 : AOI221_X1 port map( B1 => n51, B2 => A(8), C1 => n52, C2 => A(7), A =>
                           n88, ZN => n30);
   U59 : OAI22_X1 port map( A1 => n45, A2 => n55, B1 => n47, B2 => n57, ZN => 
                           n88);
   U60 : INV_X1 port map( A => A(6), ZN => n45);
   U61 : NOR2_X1 port map( A1 => SH(4), A2 => n39, ZN => B(19));
   U62 : AOI222_X1 port map( A1 => n23, A2 => n72, B1 => n77, B2 => n73, C1 => 
                           n89, C2 => SH(3), ZN => n39);
   U63 : NOR2_X1 port map( A1 => SH(4), A2 => n60, ZN => B(18));
   U64 : AOI221_X1 port map( B1 => n79, B2 => n73, C1 => n29, C2 => n72, A => 
                           n90, ZN => n60);
   U65 : INV_X1 port map( A => n91, ZN => n90);
   U66 : AOI22_X1 port map( A1 => n92, A2 => n59, B1 => n76, B2 => n78, ZN => 
                           n91);
   U67 : NOR2_X1 port map( A1 => SH(4), A2 => n80, ZN => B(17));
   U68 : AOI221_X1 port map( B1 => n11, B2 => n73, C1 => n9, C2 => n72, A => 
                           n93, ZN => n80);
   U69 : INV_X1 port map( A => n94, ZN => n93);
   U70 : AOI22_X1 port map( A1 => n92, A2 => n67, B1 => n76, B2 => n71, ZN => 
                           n94);
   U71 : NOR2_X1 port map( A1 => SH(4), A2 => n95, ZN => B(16));
   U72 : OAI221_X1 port map( B1 => n96, B2 => n38, C1 => n97, C2 => n3, A => 
                           n98, ZN => B(15));
   U73 : AOI222_X1 port map( A1 => n10, A2 => n75, B1 => n99, B2 => n58, C1 => 
                           n8, C2 => n77, ZN => n98);
   U74 : INV_X1 port map( A => n23, ZN => n96);
   U75 : OAI221_X1 port map( B1 => n100, B2 => n38, C1 => n101, C2 => n3, A => 
                           n102, ZN => B(14));
   U76 : AOI222_X1 port map( A1 => n10, A2 => n78, B1 => n99, B2 => n59, C1 => 
                           n8, C2 => n79, ZN => n102);
   U77 : INV_X1 port map( A => n28, ZN => n101);
   U78 : INV_X1 port map( A => n29, ZN => n100);
   U79 : OAI221_X1 port map( B1 => n103, B2 => n38, C1 => n104, C2 => n3, A => 
                           n105, ZN => B(13));
   U80 : AOI222_X1 port map( A1 => n10, A2 => n71, B1 => n99, B2 => n67, C1 => 
                           n8, C2 => n11, ZN => n105);
   U81 : OAI221_X1 port map( B1 => n44, B2 => n106, C1 => n46, C2 => n107, A =>
                           n108, ZN => n11);
   U82 : AOI22_X1 port map( A1 => A(22), A2 => n49, B1 => A(21), B2 => n50, ZN 
                           => n108);
   U83 : INV_X1 port map( A => A(23), ZN => n107);
   U84 : OAI222_X1 port map( A1 => n55, A2 => n109, B1 => n46, B2 => n110, C1 
                           => n57, C2 => n111, ZN => n67);
   U85 : OAI221_X1 port map( B1 => n44, B2 => n112, C1 => n46, C2 => n113, A =>
                           n114, ZN => n71);
   U86 : AOI22_X1 port map( A1 => A(26), A2 => n49, B1 => A(25), B2 => n50, ZN 
                           => n114);
   U87 : INV_X1 port map( A => n7, ZN => n104);
   U88 : OAI221_X1 port map( B1 => n44, B2 => n115, C1 => n46, C2 => n116, A =>
                           n117, ZN => n7);
   U89 : AOI22_X1 port map( A1 => A(14), A2 => n49, B1 => A(13), B2 => n50, ZN 
                           => n117);
   U90 : INV_X1 port map( A => n9, ZN => n103);
   U91 : OAI221_X1 port map( B1 => n44, B2 => n118, C1 => n46, C2 => n119, A =>
                           n120, ZN => n9);
   U92 : AOI22_X1 port map( A1 => A(18), A2 => n49, B1 => A(17), B2 => n50, ZN 
                           => n120);
   U93 : INV_X1 port map( A => n121, ZN => B(12));
   U94 : AOI221_X1 port map( B1 => n16, B2 => n6, C1 => n15, C2 => n41, A => 
                           n122, ZN => n121);
   U95 : INV_X1 port map( A => n123, ZN => n122);
   U96 : AOI222_X1 port map( A1 => n10, A2 => n74, B1 => n99, B2 => n68, C1 => 
                           n8, C2 => n17, ZN => n123);
   U97 : NOR2_X1 port map( A1 => n1, A2 => n124, ZN => n99);
   U98 : OAI221_X1 port map( B1 => n97, B2 => n38, C1 => n43, C2 => n3, A => 
                           n125, ZN => B(11));
   U99 : AOI221_X1 port map( B1 => n10, B2 => n77, C1 => n8, C2 => n23, A => 
                           n126, ZN => n125);
   U100 : NOR3_X1 port map( A1 => n1, A2 => SH(3), A3 => n69, ZN => n126);
   U101 : INV_X1 port map( A => n89, ZN => n69);
   U102 : MUX2_X1 port map( A => n75, B => n58, S => SH(2), Z => n89);
   U103 : NOR2_X1 port map( A1 => n110, A2 => n57, ZN => n58);
   U104 : OAI221_X1 port map( B1 => n44, B2 => n109, C1 => n46, C2 => n111, A 
                           => n127, ZN => n75);
   U105 : AOI22_X1 port map( A1 => A(28), A2 => n49, B1 => A(27), B2 => n50, ZN
                           => n127);
   U106 : OAI221_X1 port map( B1 => n118, B2 => n55, C1 => n119, C2 => n57, A 
                           => n128, ZN => n23);
   U107 : AOI22_X1 port map( A1 => A(22), A2 => n51, B1 => A(21), B2 => n52, ZN
                           => n128);
   U108 : OAI221_X1 port map( B1 => n44, B2 => n129, C1 => n46, C2 => n130, A 
                           => n131, ZN => n77);
   U109 : AOI22_X1 port map( A1 => A(24), A2 => n49, B1 => A(23), B2 => n50, ZN
                           => n131);
   U110 : AOI221_X1 port map( B1 => n51, B2 => A(14), C1 => n52, C2 => A(13), A
                           => n132, ZN => n43);
   U111 : OAI22_X1 port map( A1 => n133, A2 => n55, B1 => n134, B2 => n57, ZN 
                           => n132);
   U112 : INV_X1 port map( A => A(12), ZN => n133);
   U113 : INV_X1 port map( A => n22, ZN => n97);
   U114 : OAI221_X1 port map( B1 => n44, B2 => n135, C1 => n46, C2 => n136, A 
                           => n137, ZN => n22);
   U115 : AOI22_X1 port map( A1 => A(16), A2 => n49, B1 => A(15), B2 => n50, ZN
                           => n137);
   U116 : OAI221_X1 port map( B1 => n63, B2 => n3, C1 => n70, C2 => n1, A => 
                           n138, ZN => B(10));
   U117 : AOI222_X1 port map( A1 => n6, A2 => n28, B1 => n8, B2 => n29, C1 => 
                           n10, C2 => n79, ZN => n138);
   U118 : OAI221_X1 port map( B1 => n44, B2 => n130, C1 => n46, C2 => n106, A 
                           => n139, ZN => n79);
   U119 : AOI22_X1 port map( A1 => A(23), A2 => n49, B1 => A(22), B2 => n50, ZN
                           => n139);
   U120 : INV_X1 port map( A => A(24), ZN => n106);
   U121 : INV_X1 port map( A => A(25), ZN => n130);
   U122 : OAI221_X1 port map( B1 => n119, B2 => n55, C1 => n135, C2 => n57, A 
                           => n140, ZN => n29);
   U123 : AOI22_X1 port map( A1 => A(21), A2 => n51, B1 => n52, B2 => A(20), ZN
                           => n140);
   U124 : OAI221_X1 port map( B1 => n44, B2 => n136, C1 => n46, C2 => n115, A 
                           => n141, ZN => n28);
   U125 : AOI22_X1 port map( A1 => A(15), A2 => n49, B1 => A(14), B2 => n50, ZN
                           => n141);
   U126 : INV_X1 port map( A => A(16), ZN => n115);
   U127 : INV_X1 port map( A => A(17), ZN => n136);
   U128 : INV_X1 port map( A => n38, ZN => n6);
   U129 : AOI22_X1 port map( A1 => n78, A2 => n72, B1 => n59, B2 => n73, ZN => 
                           n70);
   U130 : OAI22_X1 port map( A1 => n57, A2 => n109, B1 => n55, B2 => n110, ZN 
                           => n59);
   U131 : OAI221_X1 port map( B1 => n44, B2 => n111, C1 => n46, C2 => n112, A 
                           => n142, ZN => n78);
   U132 : AOI22_X1 port map( A1 => A(27), A2 => n49, B1 => A(26), B2 => n50, ZN
                           => n142);
   U133 : INV_X1 port map( A => A(28), ZN => n112);
   U134 : INV_X1 port map( A => A(29), ZN => n111);
   U135 : AOI221_X1 port map( B1 => n51, B2 => A(13), C1 => n52, C2 => A(12), A
                           => n143, ZN => n63);
   U136 : OAI22_X1 port map( A1 => n134, A2 => n55, B1 => n84, B2 => n57, ZN =>
                           n143);
   U137 : INV_X1 port map( A => A(10), ZN => n84);
   U138 : INV_X1 port map( A => A(11), ZN => n134);
   U139 : OAI221_X1 port map( B1 => n34, B2 => n38, C1 => n95, C2 => n1, A => 
                           n144, ZN => B(0));
   U140 : AOI222_X1 port map( A1 => n10, A2 => n15, B1 => n41, B2 => n145, C1 
                           => n8, C2 => n37, ZN => n144);
   U141 : INV_X1 port map( A => n12, ZN => n37);
   U142 : AOI221_X1 port map( B1 => n51, B2 => A(11), C1 => n52, C2 => A(10), A
                           => n146, ZN => n12);
   U143 : OAI22_X1 port map( A1 => n85, A2 => n55, B1 => n54, B2 => n57, ZN => 
                           n146);
   U144 : INV_X1 port map( A => A(8), ZN => n54);
   U145 : INV_X1 port map( A => A(9), ZN => n85);
   U146 : AND2_X1 port map( A1 => n147, A2 => n148, ZN => n8);
   U147 : OAI221_X1 port map( B1 => n44, B2 => n86, C1 => n46, C2 => n149, A =>
                           n150, ZN => n145);
   U148 : AOI22_X1 port map( A1 => A(1), A2 => n49, B1 => A(0), B2 => n50, ZN 
                           => n150);
   U149 : INV_X1 port map( A => A(2), ZN => n149);
   U150 : INV_X1 port map( A => A(3), ZN => n86);
   U151 : INV_X1 port map( A => n3, ZN => n41);
   U152 : NAND2_X1 port map( A1 => n72, A2 => n1, ZN => n3);
   U153 : OAI221_X1 port map( B1 => n44, B2 => n116, C1 => n46, C2 => n151, A 
                           => n152, ZN => n15);
   U154 : AOI22_X1 port map( A1 => A(13), A2 => n49, B1 => A(12), B2 => n50, ZN
                           => n152);
   U155 : INV_X1 port map( A => A(14), ZN => n151);
   U156 : INV_X1 port map( A => A(15), ZN => n116);
   U157 : AND2_X1 port map( A1 => SH(2), A2 => n147, ZN => n10);
   U158 : NOR2_X1 port map( A1 => n153, A2 => SH(4), ZN => n147);
   U159 : AOI221_X1 port map( B1 => n17, B2 => n73, C1 => n16, C2 => n72, A => 
                           n154, ZN => n95);
   U160 : INV_X1 port map( A => n155, ZN => n154);
   U161 : AOI22_X1 port map( A1 => n92, A2 => n68, B1 => n76, B2 => n74, ZN => 
                           n155);
   U162 : OAI221_X1 port map( B1 => n44, B2 => n113, C1 => n46, C2 => n129, A 
                           => n156, ZN => n74);
   U163 : AOI22_X1 port map( A1 => A(25), A2 => n49, B1 => A(24), B2 => n50, ZN
                           => n156);
   U164 : INV_X1 port map( A => A(26), ZN => n129);
   U165 : INV_X1 port map( A => A(27), ZN => n113);
   U166 : NOR2_X1 port map( A1 => n153, A2 => SH(2), ZN => n76);
   U167 : OAI221_X1 port map( B1 => n44, B2 => n110, C1 => n46, C2 => n109, A 
                           => n157, ZN => n68);
   U168 : AOI22_X1 port map( A1 => A(29), A2 => n49, B1 => A(28), B2 => n50, ZN
                           => n157);
   U169 : INV_X1 port map( A => A(30), ZN => n109);
   U170 : INV_X1 port map( A => A(31), ZN => n110);
   U171 : NOR2_X1 port map( A1 => n148, A2 => n153, ZN => n92);
   U172 : INV_X1 port map( A => n124, ZN => n72);
   U173 : NAND2_X1 port map( A1 => n148, A2 => n153, ZN => n124);
   U174 : INV_X1 port map( A => SH(3), ZN => n153);
   U175 : OAI221_X1 port map( B1 => n44, B2 => n119, C1 => n46, C2 => n135, A 
                           => n158, ZN => n16);
   U176 : AOI22_X1 port map( A1 => A(17), A2 => n49, B1 => A(16), B2 => n50, ZN
                           => n158);
   U177 : INV_X1 port map( A => A(18), ZN => n135);
   U178 : INV_X1 port map( A => A(19), ZN => n119);
   U179 : OAI221_X1 port map( B1 => n55, B2 => n159, C1 => n118, C2 => n57, A 
                           => n160, ZN => n17);
   U180 : AOI22_X1 port map( A1 => A(23), A2 => n51, B1 => A(22), B2 => n52, ZN
                           => n160);
   U181 : INV_X1 port map( A => A(20), ZN => n118);
   U182 : INV_X1 port map( A => A(21), ZN => n159);
   U183 : NAND2_X1 port map( A1 => n73, A2 => n1, ZN => n38);
   U184 : NOR2_X1 port map( A1 => n148, A2 => SH(3), ZN => n73);
   U185 : INV_X1 port map( A => SH(2), ZN => n148);
   U186 : AOI221_X1 port map( B1 => n51, B2 => A(7), C1 => n52, C2 => A(6), A 
                           => n161, ZN => n34);
   U187 : OAI22_X1 port map( A1 => n47, A2 => n55, B1 => n64, B2 => n57, ZN => 
                           n161);
   U188 : INV_X1 port map( A => n50, ZN => n57);
   U189 : INV_X1 port map( A => A(4), ZN => n64);
   U190 : INV_X1 port map( A => n49, ZN => n55);
   U191 : INV_X1 port map( A => A(5), ZN => n47);
   U192 : INV_X1 port map( A => n46, ZN => n52);
   U193 : NAND2_X1 port map( A1 => SH(1), A2 => n162, ZN => n46);
   U194 : INV_X1 port map( A => SH(0), ZN => n162);
   U195 : INV_X1 port map( A => n44, ZN => n51);
   U196 : NAND2_X1 port map( A1 => SH(1), A2 => SH(0), ZN => n44);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Shifter_DATA_SIZE32_DW_sla_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end Shifter_DATA_SIZE32_DW_sla_0;

architecture SYN_mx2 of Shifter_DATA_SIZE32_DW_sla_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal B_31_port, B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, 
      B_25_port, B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, 
      B_19_port, B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, 
      B_13_port, B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port,
      B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, n1, n2, n3, 
      n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n173 : std_logic;

begin
   B <= ( B_31_port, B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, 
      B_25_port, B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, 
      B_19_port, B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, 
      B_13_port, B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port,
      B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, A(0) );
   
   U2 : NOR2_X2 port map( A1 => SH(2), A2 => SH(3), ZN => n75);
   U3 : INV_X1 port map( A => SH(4), ZN => n1);
   U4 : OAI21_X1 port map( B1 => SH(4), B2 => n2, A => n3, ZN => B_9_port);
   U5 : OAI21_X1 port map( B1 => SH(4), B2 => n4, A => n3, ZN => B_8_port);
   U6 : OAI21_X1 port map( B1 => SH(4), B2 => n5, A => n3, ZN => B_7_port);
   U7 : OAI21_X1 port map( B1 => SH(4), B2 => n6, A => n3, ZN => B_6_port);
   U8 : OAI21_X1 port map( B1 => SH(4), B2 => n7, A => n3, ZN => B_5_port);
   U9 : OAI21_X1 port map( B1 => SH(4), B2 => n8, A => n3, ZN => B_4_port);
   U10 : OAI21_X1 port map( B1 => SH(4), B2 => n9, A => n3, ZN => B_3_port);
   U11 : OAI221_X1 port map( B1 => n10, B2 => n11, C1 => n12, C2 => n1, A => 
                           n13, ZN => B_31_port);
   U12 : AOI222_X1 port map( A1 => n14, A2 => n15, B1 => n16, B2 => n17, C1 => 
                           n18, C2 => n19, ZN => n13);
   U13 : OAI221_X1 port map( B1 => n20, B2 => n21, C1 => n22, C2 => n23, A => 
                           n24, ZN => n17);
   U14 : AOI22_X1 port map( A1 => A(30), A2 => n25, B1 => A(31), B2 => n26, ZN 
                           => n24);
   U15 : OAI221_X1 port map( B1 => n27, B2 => n11, C1 => n28, C2 => n1, A => 
                           n29, ZN => B_30_port);
   U16 : AOI222_X1 port map( A1 => n14, A2 => n30, B1 => n16, B2 => n31, C1 => 
                           n18, C2 => n32, ZN => n29);
   U17 : OAI221_X1 port map( B1 => n33, B2 => n21, C1 => n34, C2 => n35, A => 
                           n36, ZN => n31);
   U18 : AOI22_X1 port map( A1 => A(28), A2 => n37, B1 => A(27), B2 => n38, ZN 
                           => n36);
   U19 : INV_X1 port map( A => A(30), ZN => n35);
   U20 : OAI21_X1 port map( B1 => SH(4), B2 => n39, A => n3, ZN => B_2_port);
   U21 : OAI221_X1 port map( B1 => n40, B2 => n11, C1 => n41, C2 => n1, A => 
                           n42, ZN => B_29_port);
   U22 : AOI222_X1 port map( A1 => n14, A2 => n43, B1 => n16, B2 => n44, C1 => 
                           n18, C2 => n45, ZN => n42);
   U23 : OAI221_X1 port map( B1 => n33, B2 => n23, C1 => n34, C2 => n21, A => 
                           n46, ZN => n44);
   U24 : AOI22_X1 port map( A1 => A(27), A2 => n37, B1 => A(26), B2 => n38, ZN 
                           => n46);
   U25 : INV_X1 port map( A => A(29), ZN => n21);
   U26 : OAI221_X1 port map( B1 => n47, B2 => n11, C1 => n48, C2 => n1, A => 
                           n49, ZN => B_28_port);
   U27 : AOI222_X1 port map( A1 => n14, A2 => n50, B1 => n16, B2 => n51, C1 => 
                           n18, C2 => n52, ZN => n49);
   U28 : OAI221_X1 port map( B1 => n33, B2 => n53, C1 => n34, C2 => n23, A => 
                           n54, ZN => n51);
   U29 : AOI22_X1 port map( A1 => A(26), A2 => n37, B1 => A(25), B2 => n38, ZN 
                           => n54);
   U30 : INV_X1 port map( A => A(28), ZN => n23);
   U31 : INV_X1 port map( A => A(27), ZN => n53);
   U32 : INV_X1 port map( A => n55, ZN => n16);
   U33 : OAI221_X1 port map( B1 => n10, B2 => n55, C1 => n56, C2 => n1, A => 
                           n57, ZN => B_27_port);
   U34 : AOI222_X1 port map( A1 => n58, A2 => n19, B1 => n18, B2 => n15, C1 => 
                           n14, C2 => n59, ZN => n57);
   U35 : INV_X1 port map( A => n60, ZN => n19);
   U36 : AOI221_X1 port map( B1 => n25, B2 => A(26), C1 => n26, C2 => A(27), A 
                           => n61, ZN => n10);
   U37 : INV_X1 port map( A => n62, ZN => n61);
   U38 : AOI22_X1 port map( A1 => A(25), A2 => n37, B1 => A(24), B2 => n38, ZN 
                           => n62);
   U39 : OAI221_X1 port map( B1 => n27, B2 => n55, C1 => n63, C2 => n1, A => 
                           n64, ZN => B_26_port);
   U40 : AOI222_X1 port map( A1 => n58, A2 => n32, B1 => n18, B2 => n30, C1 => 
                           n14, C2 => n65, ZN => n64);
   U41 : INV_X1 port map( A => n66, ZN => n32);
   U42 : AOI221_X1 port map( B1 => n25, B2 => A(25), C1 => n26, C2 => A(26), A 
                           => n67, ZN => n27);
   U43 : INV_X1 port map( A => n68, ZN => n67);
   U44 : AOI22_X1 port map( A1 => A(24), A2 => n37, B1 => A(23), B2 => n38, ZN 
                           => n68);
   U45 : OAI221_X1 port map( B1 => n40, B2 => n55, C1 => n2, C2 => n1, A => n69
                           , ZN => B_25_port);
   U46 : AOI222_X1 port map( A1 => n58, A2 => n45, B1 => n18, B2 => n43, C1 => 
                           n14, C2 => n70, ZN => n69);
   U47 : INV_X1 port map( A => n71, ZN => n45);
   U48 : AOI221_X1 port map( B1 => n72, B2 => n73, C1 => n74, C2 => n75, A => 
                           n76, ZN => n2);
   U49 : INV_X1 port map( A => n77, ZN => n76);
   U50 : AOI21_X1 port map( B1 => n78, B2 => n79, A => n80, ZN => n77);
   U51 : AOI221_X1 port map( B1 => n25, B2 => A(24), C1 => n26, C2 => A(25), A 
                           => n81, ZN => n40);
   U52 : INV_X1 port map( A => n82, ZN => n81);
   U53 : AOI22_X1 port map( A1 => A(23), A2 => n37, B1 => A(22), B2 => n38, ZN 
                           => n82);
   U54 : OAI221_X1 port map( B1 => n47, B2 => n55, C1 => n4, C2 => n1, A => n83
                           , ZN => B_24_port);
   U55 : AOI222_X1 port map( A1 => n58, A2 => n52, B1 => n18, B2 => n50, C1 => 
                           n14, C2 => n84, ZN => n83);
   U56 : INV_X1 port map( A => n85, ZN => n52);
   U57 : AOI221_X1 port map( B1 => n86, B2 => n73, C1 => n87, C2 => n75, A => 
                           n88, ZN => n4);
   U58 : AOI221_X1 port map( B1 => n25, B2 => A(23), C1 => n26, C2 => A(24), A 
                           => n89, ZN => n47);
   U59 : INV_X1 port map( A => n90, ZN => n89);
   U60 : AOI22_X1 port map( A1 => A(22), A2 => n37, B1 => A(21), B2 => n38, ZN 
                           => n90);
   U61 : OAI221_X1 port map( B1 => n60, B2 => n55, C1 => n5, C2 => n1, A => n91
                           , ZN => B_23_port);
   U62 : AOI222_X1 port map( A1 => n58, A2 => n15, B1 => n18, B2 => n59, C1 => 
                           n14, C2 => n92, ZN => n91);
   U63 : INV_X1 port map( A => n93, ZN => n15);
   U64 : AOI221_X1 port map( B1 => n94, B2 => n73, C1 => n95, C2 => n75, A => 
                           n88, ZN => n5);
   U65 : AOI221_X1 port map( B1 => n25, B2 => A(22), C1 => n26, C2 => A(23), A 
                           => n96, ZN => n60);
   U66 : INV_X1 port map( A => n97, ZN => n96);
   U67 : AOI22_X1 port map( A1 => A(21), A2 => n37, B1 => A(20), B2 => n38, ZN 
                           => n97);
   U68 : OAI221_X1 port map( B1 => n66, B2 => n55, C1 => n6, C2 => n1, A => n98
                           , ZN => B_22_port);
   U69 : AOI222_X1 port map( A1 => n58, A2 => n30, B1 => n18, B2 => n65, C1 => 
                           n14, C2 => n99, ZN => n98);
   U70 : INV_X1 port map( A => n100, ZN => n30);
   U71 : AOI221_X1 port map( B1 => n101, B2 => n73, C1 => n102, C2 => n75, A =>
                           n88, ZN => n6);
   U72 : AOI221_X1 port map( B1 => n25, B2 => A(21), C1 => n26, C2 => A(22), A 
                           => n103, ZN => n66);
   U73 : INV_X1 port map( A => n104, ZN => n103);
   U74 : AOI22_X1 port map( A1 => A(20), A2 => n37, B1 => A(19), B2 => n38, ZN 
                           => n104);
   U75 : OAI221_X1 port map( B1 => n71, B2 => n55, C1 => n7, C2 => n1, A => 
                           n105, ZN => B_21_port);
   U76 : AOI222_X1 port map( A1 => n58, A2 => n43, B1 => n18, B2 => n70, C1 => 
                           n14, C2 => n74, ZN => n105);
   U77 : INV_X1 port map( A => n106, ZN => n43);
   U78 : AOI221_X1 port map( B1 => n79, B2 => n73, C1 => n72, C2 => n75, A => 
                           n88, ZN => n7);
   U79 : INV_X1 port map( A => n107, ZN => n88);
   U80 : AOI221_X1 port map( B1 => n25, B2 => A(20), C1 => n26, C2 => A(21), A 
                           => n108, ZN => n71);
   U81 : OAI22_X1 port map( A1 => n109, A2 => n20, B1 => n110, B2 => n22, ZN =>
                           n108);
   U82 : INV_X1 port map( A => A(19), ZN => n109);
   U83 : OAI221_X1 port map( B1 => n85, B2 => n55, C1 => n8, C2 => n1, A => 
                           n111, ZN => B_20_port);
   U84 : AOI222_X1 port map( A1 => n58, A2 => n50, B1 => n18, B2 => n84, C1 => 
                           n14, C2 => n87, ZN => n111);
   U85 : INV_X1 port map( A => n112, ZN => n50);
   U86 : AOI21_X1 port map( B1 => n86, B2 => n75, A => n113, ZN => n8);
   U87 : AOI221_X1 port map( B1 => n25, B2 => A(19), C1 => n26, C2 => A(20), A 
                           => n114, ZN => n85);
   U88 : OAI22_X1 port map( A1 => n110, A2 => n20, B1 => n115, B2 => n22, ZN =>
                           n114);
   U89 : INV_X1 port map( A => A(18), ZN => n110);
   U90 : OAI21_X1 port map( B1 => SH(4), B2 => n116, A => n3, ZN => B_1_port);
   U91 : OAI221_X1 port map( B1 => n93, B2 => n55, C1 => n9, C2 => n1, A => 
                           n117, ZN => B_19_port);
   U92 : AOI222_X1 port map( A1 => n58, A2 => n59, B1 => n18, B2 => n92, C1 => 
                           n14, C2 => n95, ZN => n117);
   U93 : AOI21_X1 port map( B1 => n94, B2 => n75, A => n113, ZN => n9);
   U94 : AOI221_X1 port map( B1 => n25, B2 => A(18), C1 => n26, C2 => A(19), A 
                           => n118, ZN => n93);
   U95 : OAI22_X1 port map( A1 => n115, A2 => n20, B1 => n119, B2 => n22, ZN =>
                           n118);
   U96 : INV_X1 port map( A => A(17), ZN => n115);
   U97 : OAI221_X1 port map( B1 => n100, B2 => n55, C1 => n39, C2 => n1, A => 
                           n120, ZN => B_18_port);
   U98 : AOI222_X1 port map( A1 => n58, A2 => n65, B1 => n18, B2 => n99, C1 => 
                           n14, C2 => n102, ZN => n120);
   U99 : AOI21_X1 port map( B1 => n101, B2 => n75, A => n113, ZN => n39);
   U100 : AOI221_X1 port map( B1 => n25, B2 => A(17), C1 => n26, C2 => A(18), A
                           => n121, ZN => n100);
   U101 : OAI22_X1 port map( A1 => n119, A2 => n20, B1 => n122, B2 => n22, ZN 
                           => n121);
   U102 : INV_X1 port map( A => A(16), ZN => n119);
   U103 : OAI221_X1 port map( B1 => n106, B2 => n55, C1 => n116, C2 => n1, A =>
                           n123, ZN => B_17_port);
   U104 : AOI222_X1 port map( A1 => n58, A2 => n70, B1 => n18, B2 => n74, C1 =>
                           n14, C2 => n72, ZN => n123);
   U105 : INV_X1 port map( A => n11, ZN => n58);
   U106 : AOI21_X1 port map( B1 => n79, B2 => n75, A => n113, ZN => n116);
   U107 : OAI21_X1 port map( B1 => n124, B2 => n125, A => n107, ZN => n113);
   U108 : AOI221_X1 port map( B1 => n25, B2 => A(16), C1 => n26, C2 => A(17), A
                           => n126, ZN => n106);
   U109 : OAI22_X1 port map( A1 => n122, A2 => n20, B1 => n127, B2 => n22, ZN 
                           => n126);
   U110 : OAI221_X1 port map( B1 => n128, B2 => n11, C1 => n112, C2 => n55, A 
                           => n129, ZN => B_16_port);
   U111 : AOI221_X1 port map( B1 => n14, B2 => n86, C1 => n18, C2 => n87, A => 
                           n130, ZN => n129);
   U112 : INV_X1 port map( A => n3, ZN => n130);
   U113 : AND2_X1 port map( A1 => n131, A2 => n125, ZN => n18);
   U114 : AND2_X1 port map( A1 => n131, A2 => SH(2), ZN => n14);
   U115 : AND2_X1 port map( A1 => SH(3), A2 => n1, ZN => n131);
   U116 : NAND2_X1 port map( A1 => n75, A2 => n1, ZN => n55);
   U117 : AOI221_X1 port map( B1 => n25, B2 => A(15), C1 => n26, C2 => A(16), A
                           => n132, ZN => n112);
   U118 : OAI22_X1 port map( A1 => n127, A2 => n20, B1 => n133, B2 => n22, ZN 
                           => n132);
   U119 : NAND2_X1 port map( A1 => n73, A2 => n1, ZN => n11);
   U120 : INV_X1 port map( A => n84, ZN => n128);
   U121 : OAI21_X1 port map( B1 => SH(4), B2 => n12, A => n3, ZN => B_15_port);
   U122 : AOI221_X1 port map( B1 => n92, B2 => n73, C1 => n59, C2 => n75, A => 
                           n134, ZN => n12);
   U123 : INV_X1 port map( A => n135, ZN => n134);
   U124 : AOI22_X1 port map( A1 => n136, A2 => n94, B1 => n78, B2 => n95, ZN =>
                           n135);
   U125 : OAI221_X1 port map( B1 => n33, B2 => n127, C1 => n34, C2 => n122, A 
                           => n137, ZN => n59);
   U126 : AOI22_X1 port map( A1 => A(13), A2 => n37, B1 => A(12), B2 => n38, ZN
                           => n137);
   U127 : INV_X1 port map( A => A(15), ZN => n122);
   U128 : OAI21_X1 port map( B1 => SH(4), B2 => n28, A => n3, ZN => B_14_port);
   U129 : AOI221_X1 port map( B1 => n99, B2 => n73, C1 => n65, C2 => n75, A => 
                           n138, ZN => n28);
   U130 : INV_X1 port map( A => n139, ZN => n138);
   U131 : AOI22_X1 port map( A1 => n136, A2 => n101, B1 => n78, B2 => n102, ZN 
                           => n139);
   U132 : OAI221_X1 port map( B1 => n33, B2 => n133, C1 => n34, C2 => n127, A 
                           => n140, ZN => n65);
   U133 : AOI22_X1 port map( A1 => A(12), A2 => n37, B1 => A(11), B2 => n38, ZN
                           => n140);
   U134 : INV_X1 port map( A => A(14), ZN => n127);
   U135 : OAI21_X1 port map( B1 => SH(4), B2 => n41, A => n3, ZN => B_13_port);
   U136 : AOI221_X1 port map( B1 => n74, B2 => n73, C1 => n70, C2 => n75, A => 
                           n141, ZN => n41);
   U137 : INV_X1 port map( A => n142, ZN => n141);
   U138 : AOI22_X1 port map( A1 => n136, A2 => n79, B1 => n78, B2 => n72, ZN =>
                           n142);
   U139 : OAI221_X1 port map( B1 => n33, B2 => n143, C1 => n34, C2 => n144, A 
                           => n145, ZN => n72);
   U140 : AOI22_X1 port map( A1 => A(3), A2 => n37, B1 => A(2), B2 => n38, ZN 
                           => n145);
   U141 : INV_X1 port map( A => A(4), ZN => n143);
   U142 : MUX2_X1 port map( A => A(1), B => A(0), S => n34, Z => n79);
   U143 : AND2_X1 port map( A1 => SH(2), A2 => SH(3), ZN => n136);
   U144 : OAI221_X1 port map( B1 => n33, B2 => n146, C1 => n34, C2 => n133, A 
                           => n147, ZN => n70);
   U145 : AOI22_X1 port map( A1 => A(11), A2 => n37, B1 => A(10), B2 => n38, ZN
                           => n147);
   U146 : INV_X1 port map( A => A(13), ZN => n133);
   U147 : OAI221_X1 port map( B1 => n33, B2 => n148, C1 => n34, C2 => n149, A 
                           => n150, ZN => n74);
   U148 : AOI22_X1 port map( A1 => A(7), A2 => n37, B1 => A(6), B2 => n38, ZN 
                           => n150);
   U149 : OAI21_X1 port map( B1 => SH(4), B2 => n48, A => n3, ZN => B_12_port);
   U150 : AOI221_X1 port map( B1 => n87, B2 => n73, C1 => n84, C2 => n75, A => 
                           n151, ZN => n48);
   U151 : INV_X1 port map( A => n152, ZN => n151);
   U152 : AOI21_X1 port map( B1 => n78, B2 => n86, A => n80, ZN => n152);
   U153 : OAI221_X1 port map( B1 => n20, B2 => n153, C1 => n154, C2 => n22, A 
                           => n155, ZN => n86);
   U154 : AOI22_X1 port map( A1 => n25, A2 => A(3), B1 => A(4), B2 => n26, ZN 
                           => n155);
   U155 : OAI221_X1 port map( B1 => n33, B2 => n156, C1 => n34, C2 => n146, A 
                           => n157, ZN => n84);
   U156 : AOI22_X1 port map( A1 => A(10), A2 => n37, B1 => A(9), B2 => n38, ZN 
                           => n157);
   U157 : INV_X1 port map( A => A(12), ZN => n146);
   U158 : OAI221_X1 port map( B1 => n33, B2 => n158, C1 => n34, C2 => n148, A 
                           => n159, ZN => n87);
   U159 : AOI22_X1 port map( A1 => A(6), A2 => n37, B1 => A(5), B2 => n38, ZN 
                           => n159);
   U160 : INV_X1 port map( A => A(8), ZN => n148);
   U161 : OAI21_X1 port map( B1 => SH(4), B2 => n56, A => n3, ZN => B_11_port);
   U162 : AOI221_X1 port map( B1 => n95, B2 => n73, C1 => n92, C2 => n75, A => 
                           n160, ZN => n56);
   U163 : INV_X1 port map( A => n161, ZN => n160);
   U164 : AOI21_X1 port map( B1 => n78, B2 => n94, A => n80, ZN => n161);
   U165 : OAI221_X1 port map( B1 => n154, B2 => n20, C1 => n124, C2 => n22, A 
                           => n162, ZN => n94);
   U166 : AOI22_X1 port map( A1 => n25, A2 => A(2), B1 => A(3), B2 => n26, ZN 
                           => n162);
   U167 : INV_X1 port map( A => n34, ZN => n26);
   U168 : INV_X1 port map( A => n33, ZN => n25);
   U169 : OAI221_X1 port map( B1 => n33, B2 => n163, C1 => n34, C2 => n156, A 
                           => n164, ZN => n92);
   U170 : AOI22_X1 port map( A1 => A(9), A2 => n37, B1 => A(8), B2 => n38, ZN 
                           => n164);
   U171 : INV_X1 port map( A => A(11), ZN => n156);
   U172 : OAI221_X1 port map( B1 => n33, B2 => n165, C1 => n34, C2 => n158, A 
                           => n166, ZN => n95);
   U173 : AOI22_X1 port map( A1 => A(5), A2 => n37, B1 => A(4), B2 => n38, ZN 
                           => n166);
   U174 : INV_X1 port map( A => A(7), ZN => n158);
   U175 : OAI21_X1 port map( B1 => SH(4), B2 => n63, A => n3, ZN => B_10_port);
   U176 : NAND2_X1 port map( A1 => SH(4), A2 => A(0), ZN => n3);
   U177 : AOI221_X1 port map( B1 => n102, B2 => n73, C1 => n99, C2 => n75, A =>
                           n167, ZN => n63);
   U178 : INV_X1 port map( A => n168, ZN => n167);
   U179 : AOI21_X1 port map( B1 => n78, B2 => n101, A => n80, ZN => n168);
   U180 : NOR2_X1 port map( A1 => n125, A2 => n107, ZN => n80);
   U181 : NAND2_X1 port map( A1 => SH(3), A2 => A(0), ZN => n107);
   U182 : OAI222_X1 port map( A1 => n34, A2 => n153, B1 => n154, B2 => n33, C1 
                           => n124, C2 => n169, ZN => n101);
   U183 : INV_X1 port map( A => A(0), ZN => n124);
   U184 : INV_X1 port map( A => A(1), ZN => n154);
   U185 : INV_X1 port map( A => A(2), ZN => n153);
   U186 : AND2_X1 port map( A1 => SH(3), A2 => n125, ZN => n78);
   U187 : OAI221_X1 port map( B1 => n33, B2 => n149, C1 => n34, C2 => n163, A 
                           => n170, ZN => n99);
   U188 : AOI22_X1 port map( A1 => A(8), A2 => n37, B1 => A(7), B2 => n38, ZN 
                           => n170);
   U189 : INV_X1 port map( A => A(10), ZN => n163);
   U190 : INV_X1 port map( A => A(9), ZN => n149);
   U191 : NOR2_X1 port map( A1 => n125, A2 => SH(3), ZN => n73);
   U192 : INV_X1 port map( A => SH(2), ZN => n125);
   U193 : INV_X1 port map( A => n171, ZN => n102);
   U194 : AOI221_X1 port map( B1 => n37, B2 => A(4), C1 => A(3), C2 => n38, A 
                           => n172, ZN => n171);
   U195 : OAI22_X1 port map( A1 => n144, A2 => n33, B1 => n165, B2 => n34, ZN 
                           => n172);
   U196 : NAND2_X1 port map( A1 => n173, A2 => n169, ZN => n34);
   U197 : INV_X1 port map( A => A(6), ZN => n165);
   U198 : NAND2_X1 port map( A1 => SH(0), A2 => n169, ZN => n33);
   U199 : INV_X1 port map( A => SH(1), ZN => n169);
   U200 : INV_X1 port map( A => A(5), ZN => n144);
   U201 : INV_X1 port map( A => n22, ZN => n38);
   U202 : NAND2_X1 port map( A1 => SH(0), A2 => SH(1), ZN => n22);
   U203 : INV_X1 port map( A => n20, ZN => n37);
   U204 : NAND2_X1 port map( A1 => SH(1), A2 => n173, ZN => n20);
   U205 : INV_X1 port map( A => SH(0), ZN => n173);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Shifter_DATA_SIZE32_DW01_ash_0 is

   port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH : 
         in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out 
         std_logic_vector (31 downto 0));

end Shifter_DATA_SIZE32_DW01_ash_0;

architecture SYN_mx2 of Shifter_DATA_SIZE32_DW01_ash_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal SHMAG_3_port, SHMAG_2_port, SHMAG_1_port, SHMAG_0_port, 
      ML_int_1_31_port, ML_int_1_30_port, ML_int_1_29_port, ML_int_1_28_port, 
      ML_int_1_27_port, ML_int_1_26_port, ML_int_1_25_port, ML_int_1_24_port, 
      ML_int_1_23_port, ML_int_1_22_port, ML_int_1_21_port, ML_int_1_20_port, 
      ML_int_1_19_port, ML_int_1_18_port, ML_int_1_17_port, ML_int_1_16_port, 
      ML_int_1_15_port, ML_int_1_14_port, ML_int_1_13_port, ML_int_1_12_port, 
      ML_int_1_11_port, ML_int_1_10_port, ML_int_1_9_port, ML_int_1_8_port, 
      ML_int_1_7_port, ML_int_1_6_port, ML_int_1_5_port, ML_int_1_4_port, 
      ML_int_1_3_port, ML_int_1_2_port, ML_int_1_1_port, ML_int_1_0_port, 
      ML_int_2_31_port, ML_int_2_30_port, ML_int_2_29_port, ML_int_2_28_port, 
      ML_int_2_27_port, ML_int_2_26_port, ML_int_2_25_port, ML_int_2_24_port, 
      ML_int_2_23_port, ML_int_2_22_port, ML_int_2_21_port, ML_int_2_20_port, 
      ML_int_2_19_port, ML_int_2_18_port, ML_int_2_17_port, ML_int_2_16_port, 
      ML_int_2_15_port, ML_int_2_14_port, ML_int_2_13_port, ML_int_2_12_port, 
      ML_int_2_11_port, ML_int_2_10_port, ML_int_2_9_port, ML_int_2_8_port, 
      ML_int_2_7_port, ML_int_2_6_port, ML_int_2_5_port, ML_int_2_4_port, 
      ML_int_2_3_port, ML_int_2_2_port, ML_int_2_1_port, ML_int_2_0_port, 
      ML_int_3_31_port, ML_int_3_30_port, ML_int_3_29_port, ML_int_3_28_port, 
      ML_int_3_27_port, ML_int_3_26_port, ML_int_3_25_port, ML_int_3_24_port, 
      ML_int_3_23_port, ML_int_3_22_port, ML_int_3_21_port, ML_int_3_20_port, 
      ML_int_3_19_port, ML_int_3_18_port, ML_int_3_17_port, ML_int_3_16_port, 
      ML_int_3_15_port, ML_int_3_14_port, ML_int_3_13_port, ML_int_3_12_port, 
      ML_int_3_11_port, ML_int_3_10_port, ML_int_3_9_port, ML_int_3_8_port, 
      ML_int_3_7_port, ML_int_3_6_port, ML_int_3_5_port, ML_int_3_4_port, 
      ML_int_3_3_port, ML_int_3_2_port, ML_int_3_1_port, ML_int_3_0_port, 
      ML_int_4_31_port, ML_int_4_30_port, ML_int_4_29_port, ML_int_4_28_port, 
      ML_int_4_27_port, ML_int_4_26_port, ML_int_4_25_port, ML_int_4_24_port, 
      ML_int_4_23_port, ML_int_4_22_port, ML_int_4_21_port, ML_int_4_20_port, 
      ML_int_4_19_port, ML_int_4_18_port, ML_int_4_17_port, ML_int_4_16_port, 
      ML_int_4_15_port, ML_int_4_14_port, ML_int_4_13_port, ML_int_4_12_port, 
      ML_int_4_11_port, ML_int_4_10_port, ML_int_4_9_port, ML_int_4_8_port, 
      ML_int_4_7_port, ML_int_4_6_port, ML_int_4_5_port, ML_int_4_4_port, 
      ML_int_4_3_port, ML_int_4_2_port, ML_int_4_1_port, ML_int_4_0_port, n1, 
      n2, n3, n4, n5, n6, n7, n8, n9, n10 : std_logic;

begin
   
   M1_4_31 : MUX2_X1 port map( A => ML_int_4_31_port, B => ML_int_4_15_port, S 
                           => n1, Z => B(31));
   M1_4_30 : MUX2_X1 port map( A => ML_int_4_30_port, B => ML_int_4_14_port, S 
                           => n1, Z => B(30));
   M1_4_29 : MUX2_X1 port map( A => ML_int_4_29_port, B => ML_int_4_13_port, S 
                           => n1, Z => B(29));
   M1_4_28 : MUX2_X1 port map( A => ML_int_4_28_port, B => ML_int_4_12_port, S 
                           => n1, Z => B(28));
   M1_4_27 : MUX2_X1 port map( A => ML_int_4_27_port, B => ML_int_4_11_port, S 
                           => n1, Z => B(27));
   M1_4_26 : MUX2_X1 port map( A => ML_int_4_26_port, B => ML_int_4_10_port, S 
                           => n1, Z => B(26));
   M1_4_25 : MUX2_X1 port map( A => ML_int_4_25_port, B => ML_int_4_9_port, S 
                           => n1, Z => B(25));
   M1_4_24 : MUX2_X1 port map( A => ML_int_4_24_port, B => ML_int_4_8_port, S 
                           => n1, Z => B(24));
   M1_4_23 : MUX2_X1 port map( A => ML_int_4_23_port, B => ML_int_4_7_port, S 
                           => n1, Z => B(23));
   M1_4_22 : MUX2_X1 port map( A => ML_int_4_22_port, B => ML_int_4_6_port, S 
                           => n1, Z => B(22));
   M1_4_21 : MUX2_X1 port map( A => ML_int_4_21_port, B => ML_int_4_5_port, S 
                           => n1, Z => B(21));
   M1_4_20 : MUX2_X1 port map( A => ML_int_4_20_port, B => ML_int_4_4_port, S 
                           => n1, Z => B(20));
   M1_4_19 : MUX2_X1 port map( A => ML_int_4_19_port, B => ML_int_4_3_port, S 
                           => n1, Z => B(19));
   M1_4_18 : MUX2_X1 port map( A => ML_int_4_18_port, B => ML_int_4_2_port, S 
                           => n1, Z => B(18));
   M1_4_17 : MUX2_X1 port map( A => ML_int_4_17_port, B => ML_int_4_1_port, S 
                           => n1, Z => B(17));
   M1_4_16 : MUX2_X1 port map( A => ML_int_4_16_port, B => ML_int_4_0_port, S 
                           => n1, Z => B(16));
   M1_3_31 : MUX2_X1 port map( A => ML_int_3_31_port, B => ML_int_3_23_port, S 
                           => SH(3), Z => ML_int_4_31_port);
   M1_3_30 : MUX2_X1 port map( A => ML_int_3_30_port, B => ML_int_3_22_port, S 
                           => SH(3), Z => ML_int_4_30_port);
   M1_3_29 : MUX2_X1 port map( A => ML_int_3_29_port, B => ML_int_3_21_port, S 
                           => SH(3), Z => ML_int_4_29_port);
   M1_3_28 : MUX2_X1 port map( A => ML_int_3_28_port, B => ML_int_3_20_port, S 
                           => SH(3), Z => ML_int_4_28_port);
   M1_3_27 : MUX2_X1 port map( A => ML_int_3_27_port, B => ML_int_3_19_port, S 
                           => SH(3), Z => ML_int_4_27_port);
   M1_3_26 : MUX2_X1 port map( A => ML_int_3_26_port, B => ML_int_3_18_port, S 
                           => SH(3), Z => ML_int_4_26_port);
   M1_3_25 : MUX2_X1 port map( A => ML_int_3_25_port, B => ML_int_3_17_port, S 
                           => SH(3), Z => ML_int_4_25_port);
   M1_3_24 : MUX2_X1 port map( A => ML_int_3_24_port, B => ML_int_3_16_port, S 
                           => SH(3), Z => ML_int_4_24_port);
   M1_3_23 : MUX2_X1 port map( A => ML_int_3_23_port, B => ML_int_3_15_port, S 
                           => SH(3), Z => ML_int_4_23_port);
   M1_3_22 : MUX2_X1 port map( A => ML_int_3_22_port, B => ML_int_3_14_port, S 
                           => SH(3), Z => ML_int_4_22_port);
   M1_3_21 : MUX2_X1 port map( A => ML_int_3_21_port, B => ML_int_3_13_port, S 
                           => SH(3), Z => ML_int_4_21_port);
   M1_3_20 : MUX2_X1 port map( A => ML_int_3_20_port, B => ML_int_3_12_port, S 
                           => SH(3), Z => ML_int_4_20_port);
   M1_3_19 : MUX2_X1 port map( A => ML_int_3_19_port, B => ML_int_3_11_port, S 
                           => SH(3), Z => ML_int_4_19_port);
   M1_3_18 : MUX2_X1 port map( A => ML_int_3_18_port, B => ML_int_3_10_port, S 
                           => SH(3), Z => ML_int_4_18_port);
   M1_3_17 : MUX2_X1 port map( A => ML_int_3_17_port, B => ML_int_3_9_port, S 
                           => SH(3), Z => ML_int_4_17_port);
   M1_3_16 : MUX2_X1 port map( A => ML_int_3_16_port, B => ML_int_3_8_port, S 
                           => SH(3), Z => ML_int_4_16_port);
   M1_3_15 : MUX2_X1 port map( A => ML_int_3_15_port, B => ML_int_3_7_port, S 
                           => SH(3), Z => ML_int_4_15_port);
   M1_3_14 : MUX2_X1 port map( A => ML_int_3_14_port, B => ML_int_3_6_port, S 
                           => SH(3), Z => ML_int_4_14_port);
   M1_3_13 : MUX2_X1 port map( A => ML_int_3_13_port, B => ML_int_3_5_port, S 
                           => SH(3), Z => ML_int_4_13_port);
   M1_3_12 : MUX2_X1 port map( A => ML_int_3_12_port, B => ML_int_3_4_port, S 
                           => SH(3), Z => ML_int_4_12_port);
   M1_3_11 : MUX2_X1 port map( A => ML_int_3_11_port, B => ML_int_3_3_port, S 
                           => SH(3), Z => ML_int_4_11_port);
   M1_3_10 : MUX2_X1 port map( A => ML_int_3_10_port, B => ML_int_3_2_port, S 
                           => SH(3), Z => ML_int_4_10_port);
   M1_3_9 : MUX2_X1 port map( A => ML_int_3_9_port, B => ML_int_3_1_port, S => 
                           SH(3), Z => ML_int_4_9_port);
   M1_3_8 : MUX2_X1 port map( A => ML_int_3_8_port, B => ML_int_3_0_port, S => 
                           SH(3), Z => ML_int_4_8_port);
   M1_2_31 : MUX2_X1 port map( A => ML_int_2_31_port, B => ML_int_2_27_port, S 
                           => SH(2), Z => ML_int_3_31_port);
   M1_2_30 : MUX2_X1 port map( A => ML_int_2_30_port, B => ML_int_2_26_port, S 
                           => SH(2), Z => ML_int_3_30_port);
   M1_2_29 : MUX2_X1 port map( A => ML_int_2_29_port, B => ML_int_2_25_port, S 
                           => SH(2), Z => ML_int_3_29_port);
   M1_2_28 : MUX2_X1 port map( A => ML_int_2_28_port, B => ML_int_2_24_port, S 
                           => SH(2), Z => ML_int_3_28_port);
   M1_2_27 : MUX2_X1 port map( A => ML_int_2_27_port, B => ML_int_2_23_port, S 
                           => SH(2), Z => ML_int_3_27_port);
   M1_2_26 : MUX2_X1 port map( A => ML_int_2_26_port, B => ML_int_2_22_port, S 
                           => SH(2), Z => ML_int_3_26_port);
   M1_2_25 : MUX2_X1 port map( A => ML_int_2_25_port, B => ML_int_2_21_port, S 
                           => SH(2), Z => ML_int_3_25_port);
   M1_2_24 : MUX2_X1 port map( A => ML_int_2_24_port, B => ML_int_2_20_port, S 
                           => SH(2), Z => ML_int_3_24_port);
   M1_2_23 : MUX2_X1 port map( A => ML_int_2_23_port, B => ML_int_2_19_port, S 
                           => SH(2), Z => ML_int_3_23_port);
   M1_2_22 : MUX2_X1 port map( A => ML_int_2_22_port, B => ML_int_2_18_port, S 
                           => SH(2), Z => ML_int_3_22_port);
   M1_2_21 : MUX2_X1 port map( A => ML_int_2_21_port, B => ML_int_2_17_port, S 
                           => SH(2), Z => ML_int_3_21_port);
   M1_2_20 : MUX2_X1 port map( A => ML_int_2_20_port, B => ML_int_2_16_port, S 
                           => SH(2), Z => ML_int_3_20_port);
   M1_2_19 : MUX2_X1 port map( A => ML_int_2_19_port, B => ML_int_2_15_port, S 
                           => SH(2), Z => ML_int_3_19_port);
   M1_2_18 : MUX2_X1 port map( A => ML_int_2_18_port, B => ML_int_2_14_port, S 
                           => SH(2), Z => ML_int_3_18_port);
   M1_2_17 : MUX2_X1 port map( A => ML_int_2_17_port, B => ML_int_2_13_port, S 
                           => SH(2), Z => ML_int_3_17_port);
   M1_2_16 : MUX2_X1 port map( A => ML_int_2_16_port, B => ML_int_2_12_port, S 
                           => SH(2), Z => ML_int_3_16_port);
   M1_2_15 : MUX2_X1 port map( A => ML_int_2_15_port, B => ML_int_2_11_port, S 
                           => SH(2), Z => ML_int_3_15_port);
   M1_2_14 : MUX2_X1 port map( A => ML_int_2_14_port, B => ML_int_2_10_port, S 
                           => SH(2), Z => ML_int_3_14_port);
   M1_2_13 : MUX2_X1 port map( A => ML_int_2_13_port, B => ML_int_2_9_port, S 
                           => SH(2), Z => ML_int_3_13_port);
   M1_2_12 : MUX2_X1 port map( A => ML_int_2_12_port, B => ML_int_2_8_port, S 
                           => SH(2), Z => ML_int_3_12_port);
   M1_2_11 : MUX2_X1 port map( A => ML_int_2_11_port, B => ML_int_2_7_port, S 
                           => SH(2), Z => ML_int_3_11_port);
   M1_2_10 : MUX2_X1 port map( A => ML_int_2_10_port, B => ML_int_2_6_port, S 
                           => SH(2), Z => ML_int_3_10_port);
   M1_2_9 : MUX2_X1 port map( A => ML_int_2_9_port, B => ML_int_2_5_port, S => 
                           SH(2), Z => ML_int_3_9_port);
   M1_2_8 : MUX2_X1 port map( A => ML_int_2_8_port, B => ML_int_2_4_port, S => 
                           SH(2), Z => ML_int_3_8_port);
   M1_2_7 : MUX2_X1 port map( A => ML_int_2_7_port, B => ML_int_2_3_port, S => 
                           SH(2), Z => ML_int_3_7_port);
   M1_2_6 : MUX2_X1 port map( A => ML_int_2_6_port, B => ML_int_2_2_port, S => 
                           SH(2), Z => ML_int_3_6_port);
   M1_2_5 : MUX2_X1 port map( A => ML_int_2_5_port, B => ML_int_2_1_port, S => 
                           SH(2), Z => ML_int_3_5_port);
   M1_2_4 : MUX2_X1 port map( A => ML_int_2_4_port, B => ML_int_2_0_port, S => 
                           SH(2), Z => ML_int_3_4_port);
   M1_1_31 : MUX2_X1 port map( A => ML_int_1_31_port, B => ML_int_1_29_port, S 
                           => SH(1), Z => ML_int_2_31_port);
   M1_1_30 : MUX2_X1 port map( A => ML_int_1_30_port, B => ML_int_1_28_port, S 
                           => SH(1), Z => ML_int_2_30_port);
   M1_1_29 : MUX2_X1 port map( A => ML_int_1_29_port, B => ML_int_1_27_port, S 
                           => SH(1), Z => ML_int_2_29_port);
   M1_1_28 : MUX2_X1 port map( A => ML_int_1_28_port, B => ML_int_1_26_port, S 
                           => SH(1), Z => ML_int_2_28_port);
   M1_1_27 : MUX2_X1 port map( A => ML_int_1_27_port, B => ML_int_1_25_port, S 
                           => SH(1), Z => ML_int_2_27_port);
   M1_1_26 : MUX2_X1 port map( A => ML_int_1_26_port, B => ML_int_1_24_port, S 
                           => SH(1), Z => ML_int_2_26_port);
   M1_1_25 : MUX2_X1 port map( A => ML_int_1_25_port, B => ML_int_1_23_port, S 
                           => SH(1), Z => ML_int_2_25_port);
   M1_1_24 : MUX2_X1 port map( A => ML_int_1_24_port, B => ML_int_1_22_port, S 
                           => SH(1), Z => ML_int_2_24_port);
   M1_1_23 : MUX2_X1 port map( A => ML_int_1_23_port, B => ML_int_1_21_port, S 
                           => SH(1), Z => ML_int_2_23_port);
   M1_1_22 : MUX2_X1 port map( A => ML_int_1_22_port, B => ML_int_1_20_port, S 
                           => SH(1), Z => ML_int_2_22_port);
   M1_1_21 : MUX2_X1 port map( A => ML_int_1_21_port, B => ML_int_1_19_port, S 
                           => SH(1), Z => ML_int_2_21_port);
   M1_1_20 : MUX2_X1 port map( A => ML_int_1_20_port, B => ML_int_1_18_port, S 
                           => SH(1), Z => ML_int_2_20_port);
   M1_1_19 : MUX2_X1 port map( A => ML_int_1_19_port, B => ML_int_1_17_port, S 
                           => SH(1), Z => ML_int_2_19_port);
   M1_1_18 : MUX2_X1 port map( A => ML_int_1_18_port, B => ML_int_1_16_port, S 
                           => SH(1), Z => ML_int_2_18_port);
   M1_1_17 : MUX2_X1 port map( A => ML_int_1_17_port, B => ML_int_1_15_port, S 
                           => SH(1), Z => ML_int_2_17_port);
   M1_1_16 : MUX2_X1 port map( A => ML_int_1_16_port, B => ML_int_1_14_port, S 
                           => SH(1), Z => ML_int_2_16_port);
   M1_1_15 : MUX2_X1 port map( A => ML_int_1_15_port, B => ML_int_1_13_port, S 
                           => SH(1), Z => ML_int_2_15_port);
   M1_1_14 : MUX2_X1 port map( A => ML_int_1_14_port, B => ML_int_1_12_port, S 
                           => SH(1), Z => ML_int_2_14_port);
   M1_1_13 : MUX2_X1 port map( A => ML_int_1_13_port, B => ML_int_1_11_port, S 
                           => SH(1), Z => ML_int_2_13_port);
   M1_1_12 : MUX2_X1 port map( A => ML_int_1_12_port, B => ML_int_1_10_port, S 
                           => SH(1), Z => ML_int_2_12_port);
   M1_1_11 : MUX2_X1 port map( A => ML_int_1_11_port, B => ML_int_1_9_port, S 
                           => SH(1), Z => ML_int_2_11_port);
   M1_1_10 : MUX2_X1 port map( A => ML_int_1_10_port, B => ML_int_1_8_port, S 
                           => SH(1), Z => ML_int_2_10_port);
   M1_1_9 : MUX2_X1 port map( A => ML_int_1_9_port, B => ML_int_1_7_port, S => 
                           SH(1), Z => ML_int_2_9_port);
   M1_1_8 : MUX2_X1 port map( A => ML_int_1_8_port, B => ML_int_1_6_port, S => 
                           SH(1), Z => ML_int_2_8_port);
   M1_1_7 : MUX2_X1 port map( A => ML_int_1_7_port, B => ML_int_1_5_port, S => 
                           SH(1), Z => ML_int_2_7_port);
   M1_1_6 : MUX2_X1 port map( A => ML_int_1_6_port, B => ML_int_1_4_port, S => 
                           SH(1), Z => ML_int_2_6_port);
   M1_1_5 : MUX2_X1 port map( A => ML_int_1_5_port, B => ML_int_1_3_port, S => 
                           SH(1), Z => ML_int_2_5_port);
   M1_1_4 : MUX2_X1 port map( A => ML_int_1_4_port, B => ML_int_1_2_port, S => 
                           SH(1), Z => ML_int_2_4_port);
   M1_1_3 : MUX2_X1 port map( A => ML_int_1_3_port, B => ML_int_1_1_port, S => 
                           SH(1), Z => ML_int_2_3_port);
   M1_1_2 : MUX2_X1 port map( A => ML_int_1_2_port, B => ML_int_1_0_port, S => 
                           SH(1), Z => ML_int_2_2_port);
   M1_0_31 : MUX2_X1 port map( A => A(31), B => A(30), S => SH(0), Z => 
                           ML_int_1_31_port);
   M1_0_30 : MUX2_X1 port map( A => A(30), B => A(29), S => SH(0), Z => 
                           ML_int_1_30_port);
   M1_0_29 : MUX2_X1 port map( A => A(29), B => A(28), S => SH(0), Z => 
                           ML_int_1_29_port);
   M1_0_28 : MUX2_X1 port map( A => A(28), B => A(27), S => SH(0), Z => 
                           ML_int_1_28_port);
   M1_0_27 : MUX2_X1 port map( A => A(27), B => A(26), S => SH(0), Z => 
                           ML_int_1_27_port);
   M1_0_26 : MUX2_X1 port map( A => A(26), B => A(25), S => SH(0), Z => 
                           ML_int_1_26_port);
   M1_0_25 : MUX2_X1 port map( A => A(25), B => A(24), S => SH(0), Z => 
                           ML_int_1_25_port);
   M1_0_24 : MUX2_X1 port map( A => A(24), B => A(23), S => SH(0), Z => 
                           ML_int_1_24_port);
   M1_0_23 : MUX2_X1 port map( A => A(23), B => A(22), S => SH(0), Z => 
                           ML_int_1_23_port);
   M1_0_22 : MUX2_X1 port map( A => A(22), B => A(21), S => SH(0), Z => 
                           ML_int_1_22_port);
   M1_0_21 : MUX2_X1 port map( A => A(21), B => A(20), S => SH(0), Z => 
                           ML_int_1_21_port);
   M1_0_20 : MUX2_X1 port map( A => A(20), B => A(19), S => SH(0), Z => 
                           ML_int_1_20_port);
   M1_0_19 : MUX2_X1 port map( A => A(19), B => A(18), S => SH(0), Z => 
                           ML_int_1_19_port);
   M1_0_18 : MUX2_X1 port map( A => A(18), B => A(17), S => SH(0), Z => 
                           ML_int_1_18_port);
   M1_0_17 : MUX2_X1 port map( A => A(17), B => A(16), S => SH(0), Z => 
                           ML_int_1_17_port);
   M1_0_16 : MUX2_X1 port map( A => A(16), B => A(15), S => SH(0), Z => 
                           ML_int_1_16_port);
   M1_0_15 : MUX2_X1 port map( A => A(15), B => A(14), S => SH(0), Z => 
                           ML_int_1_15_port);
   M1_0_14 : MUX2_X1 port map( A => A(14), B => A(13), S => SH(0), Z => 
                           ML_int_1_14_port);
   M1_0_13 : MUX2_X1 port map( A => A(13), B => A(12), S => SH(0), Z => 
                           ML_int_1_13_port);
   M1_0_12 : MUX2_X1 port map( A => A(12), B => A(11), S => SH(0), Z => 
                           ML_int_1_12_port);
   M1_0_11 : MUX2_X1 port map( A => A(11), B => A(10), S => SH(0), Z => 
                           ML_int_1_11_port);
   M1_0_10 : MUX2_X1 port map( A => A(10), B => A(9), S => SH(0), Z => 
                           ML_int_1_10_port);
   M1_0_9 : MUX2_X1 port map( A => A(9), B => A(8), S => SH(0), Z => 
                           ML_int_1_9_port);
   M1_0_8 : MUX2_X1 port map( A => A(8), B => A(7), S => SH(0), Z => 
                           ML_int_1_8_port);
   M1_0_7 : MUX2_X1 port map( A => A(7), B => A(6), S => SH(0), Z => 
                           ML_int_1_7_port);
   M1_0_6 : MUX2_X1 port map( A => A(6), B => A(5), S => SH(0), Z => 
                           ML_int_1_6_port);
   M1_0_5 : MUX2_X1 port map( A => A(5), B => A(4), S => SH(0), Z => 
                           ML_int_1_5_port);
   M1_0_4 : MUX2_X1 port map( A => A(4), B => A(3), S => SH(0), Z => 
                           ML_int_1_4_port);
   M1_0_3 : MUX2_X1 port map( A => A(3), B => A(2), S => SH(0), Z => 
                           ML_int_1_3_port);
   M1_0_2 : MUX2_X1 port map( A => A(2), B => A(1), S => SH(0), Z => 
                           ML_int_1_2_port);
   M1_0_1 : MUX2_X1 port map( A => A(1), B => A(0), S => SH(0), Z => 
                           ML_int_1_1_port);
   U3 : INV_X1 port map( A => n2, ZN => n1);
   U4 : INV_X1 port map( A => SH(4), ZN => n2);
   U5 : AND2_X1 port map( A1 => ML_int_4_9_port, A2 => n2, ZN => B(9));
   U6 : AND2_X1 port map( A1 => ML_int_4_8_port, A2 => n2, ZN => B(8));
   U7 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => B(7));
   U8 : NOR2_X1 port map( A1 => n1, A2 => n4, ZN => B(6));
   U9 : NOR2_X1 port map( A1 => n1, A2 => n5, ZN => B(5));
   U10 : NOR2_X1 port map( A1 => n1, A2 => n6, ZN => B(4));
   U11 : NOR2_X1 port map( A1 => n1, A2 => n7, ZN => B(3));
   U12 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => B(2));
   U13 : NOR2_X1 port map( A1 => n1, A2 => n9, ZN => B(1));
   U14 : AND2_X1 port map( A1 => ML_int_4_15_port, A2 => n2, ZN => B(15));
   U15 : AND2_X1 port map( A1 => ML_int_4_14_port, A2 => n2, ZN => B(14));
   U16 : AND2_X1 port map( A1 => ML_int_4_13_port, A2 => n2, ZN => B(13));
   U17 : AND2_X1 port map( A1 => ML_int_4_12_port, A2 => n2, ZN => B(12));
   U18 : AND2_X1 port map( A1 => ML_int_4_11_port, A2 => n2, ZN => B(11));
   U19 : AND2_X1 port map( A1 => ML_int_4_10_port, A2 => n2, ZN => B(10));
   U20 : NOR2_X1 port map( A1 => SH(4), A2 => n10, ZN => B(0));
   U21 : INV_X1 port map( A => n3, ZN => ML_int_4_7_port);
   U22 : NAND2_X1 port map( A1 => ML_int_3_7_port, A2 => SHMAG_3_port, ZN => n3
                           );
   U23 : INV_X1 port map( A => n4, ZN => ML_int_4_6_port);
   U24 : NAND2_X1 port map( A1 => ML_int_3_6_port, A2 => SHMAG_3_port, ZN => n4
                           );
   U25 : INV_X1 port map( A => n5, ZN => ML_int_4_5_port);
   U26 : NAND2_X1 port map( A1 => ML_int_3_5_port, A2 => SHMAG_3_port, ZN => n5
                           );
   U27 : INV_X1 port map( A => n6, ZN => ML_int_4_4_port);
   U28 : NAND2_X1 port map( A1 => ML_int_3_4_port, A2 => SHMAG_3_port, ZN => n6
                           );
   U29 : INV_X1 port map( A => n7, ZN => ML_int_4_3_port);
   U30 : NAND2_X1 port map( A1 => ML_int_3_3_port, A2 => SHMAG_3_port, ZN => n7
                           );
   U31 : INV_X1 port map( A => n8, ZN => ML_int_4_2_port);
   U32 : NAND2_X1 port map( A1 => ML_int_3_2_port, A2 => SHMAG_3_port, ZN => n8
                           );
   U33 : INV_X1 port map( A => n9, ZN => ML_int_4_1_port);
   U34 : NAND2_X1 port map( A1 => ML_int_3_1_port, A2 => SHMAG_3_port, ZN => n9
                           );
   U35 : INV_X1 port map( A => n10, ZN => ML_int_4_0_port);
   U36 : NAND2_X1 port map( A1 => ML_int_3_0_port, A2 => SHMAG_3_port, ZN => 
                           n10);
   U37 : INV_X1 port map( A => SH(3), ZN => SHMAG_3_port);
   U38 : AND2_X1 port map( A1 => ML_int_2_3_port, A2 => SHMAG_2_port, ZN => 
                           ML_int_3_3_port);
   U39 : AND2_X1 port map( A1 => ML_int_2_2_port, A2 => SHMAG_2_port, ZN => 
                           ML_int_3_2_port);
   U40 : AND2_X1 port map( A1 => ML_int_2_1_port, A2 => SHMAG_2_port, ZN => 
                           ML_int_3_1_port);
   U41 : AND2_X1 port map( A1 => ML_int_2_0_port, A2 => SHMAG_2_port, ZN => 
                           ML_int_3_0_port);
   U42 : INV_X1 port map( A => SH(2), ZN => SHMAG_2_port);
   U43 : AND2_X1 port map( A1 => ML_int_1_1_port, A2 => SHMAG_1_port, ZN => 
                           ML_int_2_1_port);
   U44 : AND2_X1 port map( A1 => ML_int_1_0_port, A2 => SHMAG_1_port, ZN => 
                           ML_int_2_0_port);
   U45 : INV_X1 port map( A => SH(1), ZN => SHMAG_1_port);
   U46 : AND2_X1 port map( A1 => A(0), A2 => SHMAG_0_port, ZN => 
                           ML_int_1_0_port);
   U47 : INV_X1 port map( A => SH(0), ZN => SHMAG_0_port);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity BoothMul_DATA_SIZE16_STAGE10_DW01_inc_0 is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end BoothMul_DATA_SIZE16_STAGE10_DW01_inc_0;

architecture SYN_rpl of BoothMul_DATA_SIZE16_STAGE10_DW01_inc_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port : std_logic;

begin
   
   U1_1_30 : HA_X1 port map( A => A(30), B => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_1_29 : HA_X1 port map( A => A(29), B => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_1_28 : HA_X1 port map( A => A(28), B => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_1_27 : HA_X1 port map( A => A(27), B => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_1_26 : HA_X1 port map( A => A(26), B => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_1_25 : HA_X1 port map( A => A(25), B => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_1_24 : HA_X1 port map( A => A(24), B => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_1_23 : HA_X1 port map( A => A(23), B => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_1_22 : HA_X1 port map( A => A(22), B => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_1_21 : HA_X1 port map( A => A(21), B => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_1_20 : HA_X1 port map( A => A(20), B => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_1_19 : HA_X1 port map( A => A(19), B => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_1_18 : HA_X1 port map( A => A(18), B => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_1_17 : HA_X1 port map( A => A(17), B => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_1_16 : HA_X1 port map( A => A(16), B => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_1_15 : HA_X1 port map( A => A(15), B => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : XOR2_X1 port map( A => carry_31_port, B => A(31), Z => SUM(31));
   U2 : INV_X1 port map( A => A(0), ZN => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Div_DATA_SIZE32_DIV_STAGE34_SQRT_STAGE18_DW01_inc_0 is

   port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector (31
         downto 0));

end Div_DATA_SIZE32_DIV_STAGE34_SQRT_STAGE18_DW01_inc_0;

architecture SYN_rpl of Div_DATA_SIZE32_DIV_STAGE34_SQRT_STAGE18_DW01_inc_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component HA_X1
      port( A, B : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port : std_logic;

begin
   
   U1_1_30 : HA_X1 port map( A => A(30), B => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_1_29 : HA_X1 port map( A => A(29), B => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_1_28 : HA_X1 port map( A => A(28), B => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_1_27 : HA_X1 port map( A => A(27), B => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_1_26 : HA_X1 port map( A => A(26), B => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_1_25 : HA_X1 port map( A => A(25), B => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_1_24 : HA_X1 port map( A => A(24), B => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_1_23 : HA_X1 port map( A => A(23), B => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_1_22 : HA_X1 port map( A => A(22), B => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_1_21 : HA_X1 port map( A => A(21), B => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_1_20 : HA_X1 port map( A => A(20), B => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_1_19 : HA_X1 port map( A => A(19), B => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_1_18 : HA_X1 port map( A => A(18), B => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_1_17 : HA_X1 port map( A => A(17), B => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_1_16 : HA_X1 port map( A => A(16), B => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_1_15 : HA_X1 port map( A => A(15), B => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_1_14 : HA_X1 port map( A => A(14), B => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_1_13 : HA_X1 port map( A => A(13), B => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_1_12 : HA_X1 port map( A => A(12), B => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_1_11 : HA_X1 port map( A => A(11), B => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_1_10 : HA_X1 port map( A => A(10), B => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_1_9 : HA_X1 port map( A => A(9), B => carry_9_port, CO => carry_10_port, 
                           S => SUM(9));
   U1_1_8 : HA_X1 port map( A => A(8), B => carry_8_port, CO => carry_9_port, S
                           => SUM(8));
   U1_1_7 : HA_X1 port map( A => A(7), B => carry_7_port, CO => carry_8_port, S
                           => SUM(7));
   U1_1_6 : HA_X1 port map( A => A(6), B => carry_6_port, CO => carry_7_port, S
                           => SUM(6));
   U1_1_5 : HA_X1 port map( A => A(5), B => carry_5_port, CO => carry_6_port, S
                           => SUM(5));
   U1_1_4 : HA_X1 port map( A => A(4), B => carry_4_port, CO => carry_5_port, S
                           => SUM(4));
   U1_1_3 : HA_X1 port map( A => A(3), B => carry_3_port, CO => carry_4_port, S
                           => SUM(3));
   U1_1_2 : HA_X1 port map( A => A(2), B => carry_2_port, CO => carry_3_port, S
                           => SUM(2));
   U1_1_1 : HA_X1 port map( A => A(1), B => A(0), CO => carry_2_port, S => 
                           SUM(1));
   U1 : XOR2_X1 port map( A => carry_31_port, B => A(31), Z => SUM(31));
   U2 : INV_X1 port map( A => A(0), ZN => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_671 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_671;

architecture SYN_full_adder_arch of FullAdder_671 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_670 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_670;

architecture SYN_full_adder_arch of FullAdder_670 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_669 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_669;

architecture SYN_full_adder_arch of FullAdder_669 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_668 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_668;

architecture SYN_full_adder_arch of FullAdder_668 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_667 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_667;

architecture SYN_full_adder_arch of FullAdder_667 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_666 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_666;

architecture SYN_full_adder_arch of FullAdder_666 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_665 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_665;

architecture SYN_full_adder_arch of FullAdder_665 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_664 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_664;

architecture SYN_full_adder_arch of FullAdder_664 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_663 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_663;

architecture SYN_full_adder_arch of FullAdder_663 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_662 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_662;

architecture SYN_full_adder_arch of FullAdder_662 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_661 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_661;

architecture SYN_full_adder_arch of FullAdder_661 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_660 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_660;

architecture SYN_full_adder_arch of FullAdder_660 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_659 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_659;

architecture SYN_full_adder_arch of FullAdder_659 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_658 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_658;

architecture SYN_full_adder_arch of FullAdder_658 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_657 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_657;

architecture SYN_full_adder_arch of FullAdder_657 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_656 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_656;

architecture SYN_full_adder_arch of FullAdder_656 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_655 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_655;

architecture SYN_full_adder_arch of FullAdder_655 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_654 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_654;

architecture SYN_full_adder_arch of FullAdder_654 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_653 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_653;

architecture SYN_full_adder_arch of FullAdder_653 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_652 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_652;

architecture SYN_full_adder_arch of FullAdder_652 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_651 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_651;

architecture SYN_full_adder_arch of FullAdder_651 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_650 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_650;

architecture SYN_full_adder_arch of FullAdder_650 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_649 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_649;

architecture SYN_full_adder_arch of FullAdder_649 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_648 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_648;

architecture SYN_full_adder_arch of FullAdder_648 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_647 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_647;

architecture SYN_full_adder_arch of FullAdder_647 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_646 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_646;

architecture SYN_full_adder_arch of FullAdder_646 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_645 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_645;

architecture SYN_full_adder_arch of FullAdder_645 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_644 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_644;

architecture SYN_full_adder_arch of FullAdder_644 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_643 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_643;

architecture SYN_full_adder_arch of FullAdder_643 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_642 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_642;

architecture SYN_full_adder_arch of FullAdder_642 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_641 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_641;

architecture SYN_full_adder_arch of FullAdder_641 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_640 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_640;

architecture SYN_full_adder_arch of FullAdder_640 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_639 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_639;

architecture SYN_full_adder_arch of FullAdder_639 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_638 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_638;

architecture SYN_full_adder_arch of FullAdder_638 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_637 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_637;

architecture SYN_full_adder_arch of FullAdder_637 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_636 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_636;

architecture SYN_full_adder_arch of FullAdder_636 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_635 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_635;

architecture SYN_full_adder_arch of FullAdder_635 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_634 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_634;

architecture SYN_full_adder_arch of FullAdder_634 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_633 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_633;

architecture SYN_full_adder_arch of FullAdder_633 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_632 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_632;

architecture SYN_full_adder_arch of FullAdder_632 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_631 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_631;

architecture SYN_full_adder_arch of FullAdder_631 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_630 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_630;

architecture SYN_full_adder_arch of FullAdder_630 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_629 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_629;

architecture SYN_full_adder_arch of FullAdder_629 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_628 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_628;

architecture SYN_full_adder_arch of FullAdder_628 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_627 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_627;

architecture SYN_full_adder_arch of FullAdder_627 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_626 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_626;

architecture SYN_full_adder_arch of FullAdder_626 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_625 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_625;

architecture SYN_full_adder_arch of FullAdder_625 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_624 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_624;

architecture SYN_full_adder_arch of FullAdder_624 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_623 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_623;

architecture SYN_full_adder_arch of FullAdder_623 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_622 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_622;

architecture SYN_full_adder_arch of FullAdder_622 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_621 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_621;

architecture SYN_full_adder_arch of FullAdder_621 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_620 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_620;

architecture SYN_full_adder_arch of FullAdder_620 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_619 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_619;

architecture SYN_full_adder_arch of FullAdder_619 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_618 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_618;

architecture SYN_full_adder_arch of FullAdder_618 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_617 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_617;

architecture SYN_full_adder_arch of FullAdder_617 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_616 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_616;

architecture SYN_full_adder_arch of FullAdder_616 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_615 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_615;

architecture SYN_full_adder_arch of FullAdder_615 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_614 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_614;

architecture SYN_full_adder_arch of FullAdder_614 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_613 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_613;

architecture SYN_full_adder_arch of FullAdder_613 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_612 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_612;

architecture SYN_full_adder_arch of FullAdder_612 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_611 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_611;

architecture SYN_full_adder_arch of FullAdder_611 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_610 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_610;

architecture SYN_full_adder_arch of FullAdder_610 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_609 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_609;

architecture SYN_full_adder_arch of FullAdder_609 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_608 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_608;

architecture SYN_full_adder_arch of FullAdder_608 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_607 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_607;

architecture SYN_full_adder_arch of FullAdder_607 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_606 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_606;

architecture SYN_full_adder_arch of FullAdder_606 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_605 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_605;

architecture SYN_full_adder_arch of FullAdder_605 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_604 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_604;

architecture SYN_full_adder_arch of FullAdder_604 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_603 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_603;

architecture SYN_full_adder_arch of FullAdder_603 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_602 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_602;

architecture SYN_full_adder_arch of FullAdder_602 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_601 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_601;

architecture SYN_full_adder_arch of FullAdder_601 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_600 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_600;

architecture SYN_full_adder_arch of FullAdder_600 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_599 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_599;

architecture SYN_full_adder_arch of FullAdder_599 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_598 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_598;

architecture SYN_full_adder_arch of FullAdder_598 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_597 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_597;

architecture SYN_full_adder_arch of FullAdder_597 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_596 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_596;

architecture SYN_full_adder_arch of FullAdder_596 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_595 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_595;

architecture SYN_full_adder_arch of FullAdder_595 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_594 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_594;

architecture SYN_full_adder_arch of FullAdder_594 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_593 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_593;

architecture SYN_full_adder_arch of FullAdder_593 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_592 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_592;

architecture SYN_full_adder_arch of FullAdder_592 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_591 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_591;

architecture SYN_full_adder_arch of FullAdder_591 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_590 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_590;

architecture SYN_full_adder_arch of FullAdder_590 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_589 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_589;

architecture SYN_full_adder_arch of FullAdder_589 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_588 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_588;

architecture SYN_full_adder_arch of FullAdder_588 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_587 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_587;

architecture SYN_full_adder_arch of FullAdder_587 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_586 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_586;

architecture SYN_full_adder_arch of FullAdder_586 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_585 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_585;

architecture SYN_full_adder_arch of FullAdder_585 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_584 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_584;

architecture SYN_full_adder_arch of FullAdder_584 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_583 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_583;

architecture SYN_full_adder_arch of FullAdder_583 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_582 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_582;

architecture SYN_full_adder_arch of FullAdder_582 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_581 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_581;

architecture SYN_full_adder_arch of FullAdder_581 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_580 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_580;

architecture SYN_full_adder_arch of FullAdder_580 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_579 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_579;

architecture SYN_full_adder_arch of FullAdder_579 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_578 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_578;

architecture SYN_full_adder_arch of FullAdder_578 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_577 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_577;

architecture SYN_full_adder_arch of FullAdder_577 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_576 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_576;

architecture SYN_full_adder_arch of FullAdder_576 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_575 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_575;

architecture SYN_full_adder_arch of FullAdder_575 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_574 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_574;

architecture SYN_full_adder_arch of FullAdder_574 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_573 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_573;

architecture SYN_full_adder_arch of FullAdder_573 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_572 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_572;

architecture SYN_full_adder_arch of FullAdder_572 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_571 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_571;

architecture SYN_full_adder_arch of FullAdder_571 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_570 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_570;

architecture SYN_full_adder_arch of FullAdder_570 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_569 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_569;

architecture SYN_full_adder_arch of FullAdder_569 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_568 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_568;

architecture SYN_full_adder_arch of FullAdder_568 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_567 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_567;

architecture SYN_full_adder_arch of FullAdder_567 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_566 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_566;

architecture SYN_full_adder_arch of FullAdder_566 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_565 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_565;

architecture SYN_full_adder_arch of FullAdder_565 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_564 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_564;

architecture SYN_full_adder_arch of FullAdder_564 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_563 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_563;

architecture SYN_full_adder_arch of FullAdder_563 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_562 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_562;

architecture SYN_full_adder_arch of FullAdder_562 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_561 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_561;

architecture SYN_full_adder_arch of FullAdder_561 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_560 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_560;

architecture SYN_full_adder_arch of FullAdder_560 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_559 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_559;

architecture SYN_full_adder_arch of FullAdder_559 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_558 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_558;

architecture SYN_full_adder_arch of FullAdder_558 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_557 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_557;

architecture SYN_full_adder_arch of FullAdder_557 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_556 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_556;

architecture SYN_full_adder_arch of FullAdder_556 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_555 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_555;

architecture SYN_full_adder_arch of FullAdder_555 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_554 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_554;

architecture SYN_full_adder_arch of FullAdder_554 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_553 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_553;

architecture SYN_full_adder_arch of FullAdder_553 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_552 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_552;

architecture SYN_full_adder_arch of FullAdder_552 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_551 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_551;

architecture SYN_full_adder_arch of FullAdder_551 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_550 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_550;

architecture SYN_full_adder_arch of FullAdder_550 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_549 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_549;

architecture SYN_full_adder_arch of FullAdder_549 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_548 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_548;

architecture SYN_full_adder_arch of FullAdder_548 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_547 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_547;

architecture SYN_full_adder_arch of FullAdder_547 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_546 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_546;

architecture SYN_full_adder_arch of FullAdder_546 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_545 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_545;

architecture SYN_full_adder_arch of FullAdder_545 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_544 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_544;

architecture SYN_full_adder_arch of FullAdder_544 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_543 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_543;

architecture SYN_full_adder_arch of FullAdder_543 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_542 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_542;

architecture SYN_full_adder_arch of FullAdder_542 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_541 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_541;

architecture SYN_full_adder_arch of FullAdder_541 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_540 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_540;

architecture SYN_full_adder_arch of FullAdder_540 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_539 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_539;

architecture SYN_full_adder_arch of FullAdder_539 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_538 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_538;

architecture SYN_full_adder_arch of FullAdder_538 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_537 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_537;

architecture SYN_full_adder_arch of FullAdder_537 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_536 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_536;

architecture SYN_full_adder_arch of FullAdder_536 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_535 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_535;

architecture SYN_full_adder_arch of FullAdder_535 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_534 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_534;

architecture SYN_full_adder_arch of FullAdder_534 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_533 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_533;

architecture SYN_full_adder_arch of FullAdder_533 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_532 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_532;

architecture SYN_full_adder_arch of FullAdder_532 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_531 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_531;

architecture SYN_full_adder_arch of FullAdder_531 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_530 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_530;

architecture SYN_full_adder_arch of FullAdder_530 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_529 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_529;

architecture SYN_full_adder_arch of FullAdder_529 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_528 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_528;

architecture SYN_full_adder_arch of FullAdder_528 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_527 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_527;

architecture SYN_full_adder_arch of FullAdder_527 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_526 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_526;

architecture SYN_full_adder_arch of FullAdder_526 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_525 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_525;

architecture SYN_full_adder_arch of FullAdder_525 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_524 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_524;

architecture SYN_full_adder_arch of FullAdder_524 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_523 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_523;

architecture SYN_full_adder_arch of FullAdder_523 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_522 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_522;

architecture SYN_full_adder_arch of FullAdder_522 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_521 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_521;

architecture SYN_full_adder_arch of FullAdder_521 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_520 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_520;

architecture SYN_full_adder_arch of FullAdder_520 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_519 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_519;

architecture SYN_full_adder_arch of FullAdder_519 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_518 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_518;

architecture SYN_full_adder_arch of FullAdder_518 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_517 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_517;

architecture SYN_full_adder_arch of FullAdder_517 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_516 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_516;

architecture SYN_full_adder_arch of FullAdder_516 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_515 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_515;

architecture SYN_full_adder_arch of FullAdder_515 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_514 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_514;

architecture SYN_full_adder_arch of FullAdder_514 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_513 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_513;

architecture SYN_full_adder_arch of FullAdder_513 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_512 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_512;

architecture SYN_full_adder_arch of FullAdder_512 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_511 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_511;

architecture SYN_full_adder_arch of FullAdder_511 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_510 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_510;

architecture SYN_full_adder_arch of FullAdder_510 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_509 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_509;

architecture SYN_full_adder_arch of FullAdder_509 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_508 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_508;

architecture SYN_full_adder_arch of FullAdder_508 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_507 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_507;

architecture SYN_full_adder_arch of FullAdder_507 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_506 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_506;

architecture SYN_full_adder_arch of FullAdder_506 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_505 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_505;

architecture SYN_full_adder_arch of FullAdder_505 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_504 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_504;

architecture SYN_full_adder_arch of FullAdder_504 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_503 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_503;

architecture SYN_full_adder_arch of FullAdder_503 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_502 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_502;

architecture SYN_full_adder_arch of FullAdder_502 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_501 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_501;

architecture SYN_full_adder_arch of FullAdder_501 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_500 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_500;

architecture SYN_full_adder_arch of FullAdder_500 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_499 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_499;

architecture SYN_full_adder_arch of FullAdder_499 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_498 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_498;

architecture SYN_full_adder_arch of FullAdder_498 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_497 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_497;

architecture SYN_full_adder_arch of FullAdder_497 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_496 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_496;

architecture SYN_full_adder_arch of FullAdder_496 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_495 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_495;

architecture SYN_full_adder_arch of FullAdder_495 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_494 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_494;

architecture SYN_full_adder_arch of FullAdder_494 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_493 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_493;

architecture SYN_full_adder_arch of FullAdder_493 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_492 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_492;

architecture SYN_full_adder_arch of FullAdder_492 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_491 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_491;

architecture SYN_full_adder_arch of FullAdder_491 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_490 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_490;

architecture SYN_full_adder_arch of FullAdder_490 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_489 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_489;

architecture SYN_full_adder_arch of FullAdder_489 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_488 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_488;

architecture SYN_full_adder_arch of FullAdder_488 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_487 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_487;

architecture SYN_full_adder_arch of FullAdder_487 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_486 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_486;

architecture SYN_full_adder_arch of FullAdder_486 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_485 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_485;

architecture SYN_full_adder_arch of FullAdder_485 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_484 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_484;

architecture SYN_full_adder_arch of FullAdder_484 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_483 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_483;

architecture SYN_full_adder_arch of FullAdder_483 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_482 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_482;

architecture SYN_full_adder_arch of FullAdder_482 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_481 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_481;

architecture SYN_full_adder_arch of FullAdder_481 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_480 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_480;

architecture SYN_full_adder_arch of FullAdder_480 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_479 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_479;

architecture SYN_full_adder_arch of FullAdder_479 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_478 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_478;

architecture SYN_full_adder_arch of FullAdder_478 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_477 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_477;

architecture SYN_full_adder_arch of FullAdder_477 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_476 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_476;

architecture SYN_full_adder_arch of FullAdder_476 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_475 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_475;

architecture SYN_full_adder_arch of FullAdder_475 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_474 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_474;

architecture SYN_full_adder_arch of FullAdder_474 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_473 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_473;

architecture SYN_full_adder_arch of FullAdder_473 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_472 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_472;

architecture SYN_full_adder_arch of FullAdder_472 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_471 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_471;

architecture SYN_full_adder_arch of FullAdder_471 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_470 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_470;

architecture SYN_full_adder_arch of FullAdder_470 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_469 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_469;

architecture SYN_full_adder_arch of FullAdder_469 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_468 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_468;

architecture SYN_full_adder_arch of FullAdder_468 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_467 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_467;

architecture SYN_full_adder_arch of FullAdder_467 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_466 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_466;

architecture SYN_full_adder_arch of FullAdder_466 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_465 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_465;

architecture SYN_full_adder_arch of FullAdder_465 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_464 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_464;

architecture SYN_full_adder_arch of FullAdder_464 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_463 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_463;

architecture SYN_full_adder_arch of FullAdder_463 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_462 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_462;

architecture SYN_full_adder_arch of FullAdder_462 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_461 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_461;

architecture SYN_full_adder_arch of FullAdder_461 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_460 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_460;

architecture SYN_full_adder_arch of FullAdder_460 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_459 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_459;

architecture SYN_full_adder_arch of FullAdder_459 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_458 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_458;

architecture SYN_full_adder_arch of FullAdder_458 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_457 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_457;

architecture SYN_full_adder_arch of FullAdder_457 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_456 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_456;

architecture SYN_full_adder_arch of FullAdder_456 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_455 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_455;

architecture SYN_full_adder_arch of FullAdder_455 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_454 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_454;

architecture SYN_full_adder_arch of FullAdder_454 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_453 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_453;

architecture SYN_full_adder_arch of FullAdder_453 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_452 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_452;

architecture SYN_full_adder_arch of FullAdder_452 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_451 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_451;

architecture SYN_full_adder_arch of FullAdder_451 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_450 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_450;

architecture SYN_full_adder_arch of FullAdder_450 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_449 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_449;

architecture SYN_full_adder_arch of FullAdder_449 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_448 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_448;

architecture SYN_full_adder_arch of FullAdder_448 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_447 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_447;

architecture SYN_full_adder_arch of FullAdder_447 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_446 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_446;

architecture SYN_full_adder_arch of FullAdder_446 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_445 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_445;

architecture SYN_full_adder_arch of FullAdder_445 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_444 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_444;

architecture SYN_full_adder_arch of FullAdder_444 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_443 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_443;

architecture SYN_full_adder_arch of FullAdder_443 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_442 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_442;

architecture SYN_full_adder_arch of FullAdder_442 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_441 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_441;

architecture SYN_full_adder_arch of FullAdder_441 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_440 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_440;

architecture SYN_full_adder_arch of FullAdder_440 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_439 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_439;

architecture SYN_full_adder_arch of FullAdder_439 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_438 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_438;

architecture SYN_full_adder_arch of FullAdder_438 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_437 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_437;

architecture SYN_full_adder_arch of FullAdder_437 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_436 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_436;

architecture SYN_full_adder_arch of FullAdder_436 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_435 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_435;

architecture SYN_full_adder_arch of FullAdder_435 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_434 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_434;

architecture SYN_full_adder_arch of FullAdder_434 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_433 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_433;

architecture SYN_full_adder_arch of FullAdder_433 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_432 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_432;

architecture SYN_full_adder_arch of FullAdder_432 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_431 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_431;

architecture SYN_full_adder_arch of FullAdder_431 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_430 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_430;

architecture SYN_full_adder_arch of FullAdder_430 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_429 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_429;

architecture SYN_full_adder_arch of FullAdder_429 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_428 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_428;

architecture SYN_full_adder_arch of FullAdder_428 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_427 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_427;

architecture SYN_full_adder_arch of FullAdder_427 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_426 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_426;

architecture SYN_full_adder_arch of FullAdder_426 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_425 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_425;

architecture SYN_full_adder_arch of FullAdder_425 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_424 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_424;

architecture SYN_full_adder_arch of FullAdder_424 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_423 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_423;

architecture SYN_full_adder_arch of FullAdder_423 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_422 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_422;

architecture SYN_full_adder_arch of FullAdder_422 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_421 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_421;

architecture SYN_full_adder_arch of FullAdder_421 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_420 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_420;

architecture SYN_full_adder_arch of FullAdder_420 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_419 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_419;

architecture SYN_full_adder_arch of FullAdder_419 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_418 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_418;

architecture SYN_full_adder_arch of FullAdder_418 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_417 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_417;

architecture SYN_full_adder_arch of FullAdder_417 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_416 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_416;

architecture SYN_full_adder_arch of FullAdder_416 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_415 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_415;

architecture SYN_full_adder_arch of FullAdder_415 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_414 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_414;

architecture SYN_full_adder_arch of FullAdder_414 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_413 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_413;

architecture SYN_full_adder_arch of FullAdder_413 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_412 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_412;

architecture SYN_full_adder_arch of FullAdder_412 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_411 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_411;

architecture SYN_full_adder_arch of FullAdder_411 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_410 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_410;

architecture SYN_full_adder_arch of FullAdder_410 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_409 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_409;

architecture SYN_full_adder_arch of FullAdder_409 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_408 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_408;

architecture SYN_full_adder_arch of FullAdder_408 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_407 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_407;

architecture SYN_full_adder_arch of FullAdder_407 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_406 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_406;

architecture SYN_full_adder_arch of FullAdder_406 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_405 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_405;

architecture SYN_full_adder_arch of FullAdder_405 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_404 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_404;

architecture SYN_full_adder_arch of FullAdder_404 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_403 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_403;

architecture SYN_full_adder_arch of FullAdder_403 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_402 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_402;

architecture SYN_full_adder_arch of FullAdder_402 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_401 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_401;

architecture SYN_full_adder_arch of FullAdder_401 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_400 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_400;

architecture SYN_full_adder_arch of FullAdder_400 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_399 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_399;

architecture SYN_full_adder_arch of FullAdder_399 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_398 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_398;

architecture SYN_full_adder_arch of FullAdder_398 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_397 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_397;

architecture SYN_full_adder_arch of FullAdder_397 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_396 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_396;

architecture SYN_full_adder_arch of FullAdder_396 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_395 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_395;

architecture SYN_full_adder_arch of FullAdder_395 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_394 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_394;

architecture SYN_full_adder_arch of FullAdder_394 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_393 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_393;

architecture SYN_full_adder_arch of FullAdder_393 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_392 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_392;

architecture SYN_full_adder_arch of FullAdder_392 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_391 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_391;

architecture SYN_full_adder_arch of FullAdder_391 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_390 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_390;

architecture SYN_full_adder_arch of FullAdder_390 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_389 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_389;

architecture SYN_full_adder_arch of FullAdder_389 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_388 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_388;

architecture SYN_full_adder_arch of FullAdder_388 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_387 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_387;

architecture SYN_full_adder_arch of FullAdder_387 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_386 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_386;

architecture SYN_full_adder_arch of FullAdder_386 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_385 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_385;

architecture SYN_full_adder_arch of FullAdder_385 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_384 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_384;

architecture SYN_full_adder_arch of FullAdder_384 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_383 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_383;

architecture SYN_full_adder_arch of FullAdder_383 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_382 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_382;

architecture SYN_full_adder_arch of FullAdder_382 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_381 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_381;

architecture SYN_full_adder_arch of FullAdder_381 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_380 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_380;

architecture SYN_full_adder_arch of FullAdder_380 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_379 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_379;

architecture SYN_full_adder_arch of FullAdder_379 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_378 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_378;

architecture SYN_full_adder_arch of FullAdder_378 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_377 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_377;

architecture SYN_full_adder_arch of FullAdder_377 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_376 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_376;

architecture SYN_full_adder_arch of FullAdder_376 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_375 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_375;

architecture SYN_full_adder_arch of FullAdder_375 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_374 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_374;

architecture SYN_full_adder_arch of FullAdder_374 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_373 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_373;

architecture SYN_full_adder_arch of FullAdder_373 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_372 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_372;

architecture SYN_full_adder_arch of FullAdder_372 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_371 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_371;

architecture SYN_full_adder_arch of FullAdder_371 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_370 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_370;

architecture SYN_full_adder_arch of FullAdder_370 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_369 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_369;

architecture SYN_full_adder_arch of FullAdder_369 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_368 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_368;

architecture SYN_full_adder_arch of FullAdder_368 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_367 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_367;

architecture SYN_full_adder_arch of FullAdder_367 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_366 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_366;

architecture SYN_full_adder_arch of FullAdder_366 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_365 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_365;

architecture SYN_full_adder_arch of FullAdder_365 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_364 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_364;

architecture SYN_full_adder_arch of FullAdder_364 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_363 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_363;

architecture SYN_full_adder_arch of FullAdder_363 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_362 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_362;

architecture SYN_full_adder_arch of FullAdder_362 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_361 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_361;

architecture SYN_full_adder_arch of FullAdder_361 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_360 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_360;

architecture SYN_full_adder_arch of FullAdder_360 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_359 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_359;

architecture SYN_full_adder_arch of FullAdder_359 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_358 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_358;

architecture SYN_full_adder_arch of FullAdder_358 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_357 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_357;

architecture SYN_full_adder_arch of FullAdder_357 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_356 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_356;

architecture SYN_full_adder_arch of FullAdder_356 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_355 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_355;

architecture SYN_full_adder_arch of FullAdder_355 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_354 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_354;

architecture SYN_full_adder_arch of FullAdder_354 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_353 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_353;

architecture SYN_full_adder_arch of FullAdder_353 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_352 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_352;

architecture SYN_full_adder_arch of FullAdder_352 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_351 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_351;

architecture SYN_full_adder_arch of FullAdder_351 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_350 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_350;

architecture SYN_full_adder_arch of FullAdder_350 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_349 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_349;

architecture SYN_full_adder_arch of FullAdder_349 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_348 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_348;

architecture SYN_full_adder_arch of FullAdder_348 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_347 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_347;

architecture SYN_full_adder_arch of FullAdder_347 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_346 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_346;

architecture SYN_full_adder_arch of FullAdder_346 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_345 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_345;

architecture SYN_full_adder_arch of FullAdder_345 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_344 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_344;

architecture SYN_full_adder_arch of FullAdder_344 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_343 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_343;

architecture SYN_full_adder_arch of FullAdder_343 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_342 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_342;

architecture SYN_full_adder_arch of FullAdder_342 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_341 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_341;

architecture SYN_full_adder_arch of FullAdder_341 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_340 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_340;

architecture SYN_full_adder_arch of FullAdder_340 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_339 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_339;

architecture SYN_full_adder_arch of FullAdder_339 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_338 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_338;

architecture SYN_full_adder_arch of FullAdder_338 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_337 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_337;

architecture SYN_full_adder_arch of FullAdder_337 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_336 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_336;

architecture SYN_full_adder_arch of FullAdder_336 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_335 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_335;

architecture SYN_full_adder_arch of FullAdder_335 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_334 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_334;

architecture SYN_full_adder_arch of FullAdder_334 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_333 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_333;

architecture SYN_full_adder_arch of FullAdder_333 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_332 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_332;

architecture SYN_full_adder_arch of FullAdder_332 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_331 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_331;

architecture SYN_full_adder_arch of FullAdder_331 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_330 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_330;

architecture SYN_full_adder_arch of FullAdder_330 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_329 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_329;

architecture SYN_full_adder_arch of FullAdder_329 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_328 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_328;

architecture SYN_full_adder_arch of FullAdder_328 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_327 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_327;

architecture SYN_full_adder_arch of FullAdder_327 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_326 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_326;

architecture SYN_full_adder_arch of FullAdder_326 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_325 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_325;

architecture SYN_full_adder_arch of FullAdder_325 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_324 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_324;

architecture SYN_full_adder_arch of FullAdder_324 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_323 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_323;

architecture SYN_full_adder_arch of FullAdder_323 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_322 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_322;

architecture SYN_full_adder_arch of FullAdder_322 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_321 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_321;

architecture SYN_full_adder_arch of FullAdder_321 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_320 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_320;

architecture SYN_full_adder_arch of FullAdder_320 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_319 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_319;

architecture SYN_full_adder_arch of FullAdder_319 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_318 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_318;

architecture SYN_full_adder_arch of FullAdder_318 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_317 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_317;

architecture SYN_full_adder_arch of FullAdder_317 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_316 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_316;

architecture SYN_full_adder_arch of FullAdder_316 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_315 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_315;

architecture SYN_full_adder_arch of FullAdder_315 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_314 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_314;

architecture SYN_full_adder_arch of FullAdder_314 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_313 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_313;

architecture SYN_full_adder_arch of FullAdder_313 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_312 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_312;

architecture SYN_full_adder_arch of FullAdder_312 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_311 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_311;

architecture SYN_full_adder_arch of FullAdder_311 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_310 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_310;

architecture SYN_full_adder_arch of FullAdder_310 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_309 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_309;

architecture SYN_full_adder_arch of FullAdder_309 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_308 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_308;

architecture SYN_full_adder_arch of FullAdder_308 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_307 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_307;

architecture SYN_full_adder_arch of FullAdder_307 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_306 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_306;

architecture SYN_full_adder_arch of FullAdder_306 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_305 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_305;

architecture SYN_full_adder_arch of FullAdder_305 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_304 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_304;

architecture SYN_full_adder_arch of FullAdder_304 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_303 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_303;

architecture SYN_full_adder_arch of FullAdder_303 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_302 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_302;

architecture SYN_full_adder_arch of FullAdder_302 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_301 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_301;

architecture SYN_full_adder_arch of FullAdder_301 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_300 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_300;

architecture SYN_full_adder_arch of FullAdder_300 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_299 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_299;

architecture SYN_full_adder_arch of FullAdder_299 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_298 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_298;

architecture SYN_full_adder_arch of FullAdder_298 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_297 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_297;

architecture SYN_full_adder_arch of FullAdder_297 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_296 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_296;

architecture SYN_full_adder_arch of FullAdder_296 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_295 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_295;

architecture SYN_full_adder_arch of FullAdder_295 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_294 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_294;

architecture SYN_full_adder_arch of FullAdder_294 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_293 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_293;

architecture SYN_full_adder_arch of FullAdder_293 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_292 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_292;

architecture SYN_full_adder_arch of FullAdder_292 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_291 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_291;

architecture SYN_full_adder_arch of FullAdder_291 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_290 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_290;

architecture SYN_full_adder_arch of FullAdder_290 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_289 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_289;

architecture SYN_full_adder_arch of FullAdder_289 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_288 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_288;

architecture SYN_full_adder_arch of FullAdder_288 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_287 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_287;

architecture SYN_full_adder_arch of FullAdder_287 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_286 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_286;

architecture SYN_full_adder_arch of FullAdder_286 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_285 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_285;

architecture SYN_full_adder_arch of FullAdder_285 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_284 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_284;

architecture SYN_full_adder_arch of FullAdder_284 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_283 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_283;

architecture SYN_full_adder_arch of FullAdder_283 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_282 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_282;

architecture SYN_full_adder_arch of FullAdder_282 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_281 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_281;

architecture SYN_full_adder_arch of FullAdder_281 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_280 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_280;

architecture SYN_full_adder_arch of FullAdder_280 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_279 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_279;

architecture SYN_full_adder_arch of FullAdder_279 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_278 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_278;

architecture SYN_full_adder_arch of FullAdder_278 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_277 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_277;

architecture SYN_full_adder_arch of FullAdder_277 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_276 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_276;

architecture SYN_full_adder_arch of FullAdder_276 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_275 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_275;

architecture SYN_full_adder_arch of FullAdder_275 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_274 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_274;

architecture SYN_full_adder_arch of FullAdder_274 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_273 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_273;

architecture SYN_full_adder_arch of FullAdder_273 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_272 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_272;

architecture SYN_full_adder_arch of FullAdder_272 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_271 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_271;

architecture SYN_full_adder_arch of FullAdder_271 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_270 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_270;

architecture SYN_full_adder_arch of FullAdder_270 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_269 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_269;

architecture SYN_full_adder_arch of FullAdder_269 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_268 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_268;

architecture SYN_full_adder_arch of FullAdder_268 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_267 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_267;

architecture SYN_full_adder_arch of FullAdder_267 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_266 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_266;

architecture SYN_full_adder_arch of FullAdder_266 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_265 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_265;

architecture SYN_full_adder_arch of FullAdder_265 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_264 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_264;

architecture SYN_full_adder_arch of FullAdder_264 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_263 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_263;

architecture SYN_full_adder_arch of FullAdder_263 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_262 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_262;

architecture SYN_full_adder_arch of FullAdder_262 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_261 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_261;

architecture SYN_full_adder_arch of FullAdder_261 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_260 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_260;

architecture SYN_full_adder_arch of FullAdder_260 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_259 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_259;

architecture SYN_full_adder_arch of FullAdder_259 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_258 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_258;

architecture SYN_full_adder_arch of FullAdder_258 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_257 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_257;

architecture SYN_full_adder_arch of FullAdder_257 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_256 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_256;

architecture SYN_full_adder_arch of FullAdder_256 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_255 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_255;

architecture SYN_full_adder_arch of FullAdder_255 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_254 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_254;

architecture SYN_full_adder_arch of FullAdder_254 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_253 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_253;

architecture SYN_full_adder_arch of FullAdder_253 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_252 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_252;

architecture SYN_full_adder_arch of FullAdder_252 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_251 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_251;

architecture SYN_full_adder_arch of FullAdder_251 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_250 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_250;

architecture SYN_full_adder_arch of FullAdder_250 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_249 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_249;

architecture SYN_full_adder_arch of FullAdder_249 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_248 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_248;

architecture SYN_full_adder_arch of FullAdder_248 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_247 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_247;

architecture SYN_full_adder_arch of FullAdder_247 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_246 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_246;

architecture SYN_full_adder_arch of FullAdder_246 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_245 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_245;

architecture SYN_full_adder_arch of FullAdder_245 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_244 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_244;

architecture SYN_full_adder_arch of FullAdder_244 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_243 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_243;

architecture SYN_full_adder_arch of FullAdder_243 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_242 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_242;

architecture SYN_full_adder_arch of FullAdder_242 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_241 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_241;

architecture SYN_full_adder_arch of FullAdder_241 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_240 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_240;

architecture SYN_full_adder_arch of FullAdder_240 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_239 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_239;

architecture SYN_full_adder_arch of FullAdder_239 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_238 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_238;

architecture SYN_full_adder_arch of FullAdder_238 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_237 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_237;

architecture SYN_full_adder_arch of FullAdder_237 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_236 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_236;

architecture SYN_full_adder_arch of FullAdder_236 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_235 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_235;

architecture SYN_full_adder_arch of FullAdder_235 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_234 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_234;

architecture SYN_full_adder_arch of FullAdder_234 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_233 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_233;

architecture SYN_full_adder_arch of FullAdder_233 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_232 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_232;

architecture SYN_full_adder_arch of FullAdder_232 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_231 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_231;

architecture SYN_full_adder_arch of FullAdder_231 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_230 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_230;

architecture SYN_full_adder_arch of FullAdder_230 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_229 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_229;

architecture SYN_full_adder_arch of FullAdder_229 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_228 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_228;

architecture SYN_full_adder_arch of FullAdder_228 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_227 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_227;

architecture SYN_full_adder_arch of FullAdder_227 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_226 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_226;

architecture SYN_full_adder_arch of FullAdder_226 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_225 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_225;

architecture SYN_full_adder_arch of FullAdder_225 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_224 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_224;

architecture SYN_full_adder_arch of FullAdder_224 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_223 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_223;

architecture SYN_full_adder_arch of FullAdder_223 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_222 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_222;

architecture SYN_full_adder_arch of FullAdder_222 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_221 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_221;

architecture SYN_full_adder_arch of FullAdder_221 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_220 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_220;

architecture SYN_full_adder_arch of FullAdder_220 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_219 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_219;

architecture SYN_full_adder_arch of FullAdder_219 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_218 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_218;

architecture SYN_full_adder_arch of FullAdder_218 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_217 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_217;

architecture SYN_full_adder_arch of FullAdder_217 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_216 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_216;

architecture SYN_full_adder_arch of FullAdder_216 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_215 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_215;

architecture SYN_full_adder_arch of FullAdder_215 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_214 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_214;

architecture SYN_full_adder_arch of FullAdder_214 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_213 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_213;

architecture SYN_full_adder_arch of FullAdder_213 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_212 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_212;

architecture SYN_full_adder_arch of FullAdder_212 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_211 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_211;

architecture SYN_full_adder_arch of FullAdder_211 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_210 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_210;

architecture SYN_full_adder_arch of FullAdder_210 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_209 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_209;

architecture SYN_full_adder_arch of FullAdder_209 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_208 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_208;

architecture SYN_full_adder_arch of FullAdder_208 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_207 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_207;

architecture SYN_full_adder_arch of FullAdder_207 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_206 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_206;

architecture SYN_full_adder_arch of FullAdder_206 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_205 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_205;

architecture SYN_full_adder_arch of FullAdder_205 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_204 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_204;

architecture SYN_full_adder_arch of FullAdder_204 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_203 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_203;

architecture SYN_full_adder_arch of FullAdder_203 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_202 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_202;

architecture SYN_full_adder_arch of FullAdder_202 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_201 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_201;

architecture SYN_full_adder_arch of FullAdder_201 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_200 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_200;

architecture SYN_full_adder_arch of FullAdder_200 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_199 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_199;

architecture SYN_full_adder_arch of FullAdder_199 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_198 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_198;

architecture SYN_full_adder_arch of FullAdder_198 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_197 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_197;

architecture SYN_full_adder_arch of FullAdder_197 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_196 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_196;

architecture SYN_full_adder_arch of FullAdder_196 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_195 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_195;

architecture SYN_full_adder_arch of FullAdder_195 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_194 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_194;

architecture SYN_full_adder_arch of FullAdder_194 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_193 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_193;

architecture SYN_full_adder_arch of FullAdder_193 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_192 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_192;

architecture SYN_full_adder_arch of FullAdder_192 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_191 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_191;

architecture SYN_full_adder_arch of FullAdder_191 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_190 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_190;

architecture SYN_full_adder_arch of FullAdder_190 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_189 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_189;

architecture SYN_full_adder_arch of FullAdder_189 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_188 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_188;

architecture SYN_full_adder_arch of FullAdder_188 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_187 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_187;

architecture SYN_full_adder_arch of FullAdder_187 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_186 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_186;

architecture SYN_full_adder_arch of FullAdder_186 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_185 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_185;

architecture SYN_full_adder_arch of FullAdder_185 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_184 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_184;

architecture SYN_full_adder_arch of FullAdder_184 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_183 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_183;

architecture SYN_full_adder_arch of FullAdder_183 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_182 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_182;

architecture SYN_full_adder_arch of FullAdder_182 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_181 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_181;

architecture SYN_full_adder_arch of FullAdder_181 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_180 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_180;

architecture SYN_full_adder_arch of FullAdder_180 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_179 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_179;

architecture SYN_full_adder_arch of FullAdder_179 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_178 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_178;

architecture SYN_full_adder_arch of FullAdder_178 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_177 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_177;

architecture SYN_full_adder_arch of FullAdder_177 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_176 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_176;

architecture SYN_full_adder_arch of FullAdder_176 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_175 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_175;

architecture SYN_full_adder_arch of FullAdder_175 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_174 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_174;

architecture SYN_full_adder_arch of FullAdder_174 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_173 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_173;

architecture SYN_full_adder_arch of FullAdder_173 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_172 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_172;

architecture SYN_full_adder_arch of FullAdder_172 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_171 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_171;

architecture SYN_full_adder_arch of FullAdder_171 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_170 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_170;

architecture SYN_full_adder_arch of FullAdder_170 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_169 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_169;

architecture SYN_full_adder_arch of FullAdder_169 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_168 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_168;

architecture SYN_full_adder_arch of FullAdder_168 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_167 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_167;

architecture SYN_full_adder_arch of FullAdder_167 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_166 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_166;

architecture SYN_full_adder_arch of FullAdder_166 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_165 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_165;

architecture SYN_full_adder_arch of FullAdder_165 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_164 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_164;

architecture SYN_full_adder_arch of FullAdder_164 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_163 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_163;

architecture SYN_full_adder_arch of FullAdder_163 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_162 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_162;

architecture SYN_full_adder_arch of FullAdder_162 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_161 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_161;

architecture SYN_full_adder_arch of FullAdder_161 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_160 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_160;

architecture SYN_full_adder_arch of FullAdder_160 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_159 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_159;

architecture SYN_full_adder_arch of FullAdder_159 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_158 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_158;

architecture SYN_full_adder_arch of FullAdder_158 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_157 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_157;

architecture SYN_full_adder_arch of FullAdder_157 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_156 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_156;

architecture SYN_full_adder_arch of FullAdder_156 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_155 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_155;

architecture SYN_full_adder_arch of FullAdder_155 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_154 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_154;

architecture SYN_full_adder_arch of FullAdder_154 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_153 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_153;

architecture SYN_full_adder_arch of FullAdder_153 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_152 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_152;

architecture SYN_full_adder_arch of FullAdder_152 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_151 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_151;

architecture SYN_full_adder_arch of FullAdder_151 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_150 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_150;

architecture SYN_full_adder_arch of FullAdder_150 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_149 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_149;

architecture SYN_full_adder_arch of FullAdder_149 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_148 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_148;

architecture SYN_full_adder_arch of FullAdder_148 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_147 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_147;

architecture SYN_full_adder_arch of FullAdder_147 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_146 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_146;

architecture SYN_full_adder_arch of FullAdder_146 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_145 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_145;

architecture SYN_full_adder_arch of FullAdder_145 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_144 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_144;

architecture SYN_full_adder_arch of FullAdder_144 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_143 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_143;

architecture SYN_full_adder_arch of FullAdder_143 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_142 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_142;

architecture SYN_full_adder_arch of FullAdder_142 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_141 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_141;

architecture SYN_full_adder_arch of FullAdder_141 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_140 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_140;

architecture SYN_full_adder_arch of FullAdder_140 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_139 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_139;

architecture SYN_full_adder_arch of FullAdder_139 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_138 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_138;

architecture SYN_full_adder_arch of FullAdder_138 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_137 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_137;

architecture SYN_full_adder_arch of FullAdder_137 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_136 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_136;

architecture SYN_full_adder_arch of FullAdder_136 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_135 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_135;

architecture SYN_full_adder_arch of FullAdder_135 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_134 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_134;

architecture SYN_full_adder_arch of FullAdder_134 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_133 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_133;

architecture SYN_full_adder_arch of FullAdder_133 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_132 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_132;

architecture SYN_full_adder_arch of FullAdder_132 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_131 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_131;

architecture SYN_full_adder_arch of FullAdder_131 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_130 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_130;

architecture SYN_full_adder_arch of FullAdder_130 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_129 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_129;

architecture SYN_full_adder_arch of FullAdder_129 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_128 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_128;

architecture SYN_full_adder_arch of FullAdder_128 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_127 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_127;

architecture SYN_full_adder_arch of FullAdder_127 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_126 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_126;

architecture SYN_full_adder_arch of FullAdder_126 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_125 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_125;

architecture SYN_full_adder_arch of FullAdder_125 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_124 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_124;

architecture SYN_full_adder_arch of FullAdder_124 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_123 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_123;

architecture SYN_full_adder_arch of FullAdder_123 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_122 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_122;

architecture SYN_full_adder_arch of FullAdder_122 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_121 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_121;

architecture SYN_full_adder_arch of FullAdder_121 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_120 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_120;

architecture SYN_full_adder_arch of FullAdder_120 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_119 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_119;

architecture SYN_full_adder_arch of FullAdder_119 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_118 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_118;

architecture SYN_full_adder_arch of FullAdder_118 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_117 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_117;

architecture SYN_full_adder_arch of FullAdder_117 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_116 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_116;

architecture SYN_full_adder_arch of FullAdder_116 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_115 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_115;

architecture SYN_full_adder_arch of FullAdder_115 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_114 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_114;

architecture SYN_full_adder_arch of FullAdder_114 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_113 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_113;

architecture SYN_full_adder_arch of FullAdder_113 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_112 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_112;

architecture SYN_full_adder_arch of FullAdder_112 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_111 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_111;

architecture SYN_full_adder_arch of FullAdder_111 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_110 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_110;

architecture SYN_full_adder_arch of FullAdder_110 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_109 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_109;

architecture SYN_full_adder_arch of FullAdder_109 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_108 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_108;

architecture SYN_full_adder_arch of FullAdder_108 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_107 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_107;

architecture SYN_full_adder_arch of FullAdder_107 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_106 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_106;

architecture SYN_full_adder_arch of FullAdder_106 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_105 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_105;

architecture SYN_full_adder_arch of FullAdder_105 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_104 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_104;

architecture SYN_full_adder_arch of FullAdder_104 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_103 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_103;

architecture SYN_full_adder_arch of FullAdder_103 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_102 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_102;

architecture SYN_full_adder_arch of FullAdder_102 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_101 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_101;

architecture SYN_full_adder_arch of FullAdder_101 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_100 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_100;

architecture SYN_full_adder_arch of FullAdder_100 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_99 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_99;

architecture SYN_full_adder_arch of FullAdder_99 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_98 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_98;

architecture SYN_full_adder_arch of FullAdder_98 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_97 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_97;

architecture SYN_full_adder_arch of FullAdder_97 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_96 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_96;

architecture SYN_full_adder_arch of FullAdder_96 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_95 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_95;

architecture SYN_full_adder_arch of FullAdder_95 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_94 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_94;

architecture SYN_full_adder_arch of FullAdder_94 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_93 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_93;

architecture SYN_full_adder_arch of FullAdder_93 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_92 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_92;

architecture SYN_full_adder_arch of FullAdder_92 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_91 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_91;

architecture SYN_full_adder_arch of FullAdder_91 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_90 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_90;

architecture SYN_full_adder_arch of FullAdder_90 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_89 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_89;

architecture SYN_full_adder_arch of FullAdder_89 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_88 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_88;

architecture SYN_full_adder_arch of FullAdder_88 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_87 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_87;

architecture SYN_full_adder_arch of FullAdder_87 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_86 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_86;

architecture SYN_full_adder_arch of FullAdder_86 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_85 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_85;

architecture SYN_full_adder_arch of FullAdder_85 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_84 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_84;

architecture SYN_full_adder_arch of FullAdder_84 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_83 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_83;

architecture SYN_full_adder_arch of FullAdder_83 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_82 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_82;

architecture SYN_full_adder_arch of FullAdder_82 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_81 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_81;

architecture SYN_full_adder_arch of FullAdder_81 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_80 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_80;

architecture SYN_full_adder_arch of FullAdder_80 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_79 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_79;

architecture SYN_full_adder_arch of FullAdder_79 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_78 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_78;

architecture SYN_full_adder_arch of FullAdder_78 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_77 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_77;

architecture SYN_full_adder_arch of FullAdder_77 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_76 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_76;

architecture SYN_full_adder_arch of FullAdder_76 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_75 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_75;

architecture SYN_full_adder_arch of FullAdder_75 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_74 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_74;

architecture SYN_full_adder_arch of FullAdder_74 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_73 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_73;

architecture SYN_full_adder_arch of FullAdder_73 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_72 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_72;

architecture SYN_full_adder_arch of FullAdder_72 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_71 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_71;

architecture SYN_full_adder_arch of FullAdder_71 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_70 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_70;

architecture SYN_full_adder_arch of FullAdder_70 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_69 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_69;

architecture SYN_full_adder_arch of FullAdder_69 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_68 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_68;

architecture SYN_full_adder_arch of FullAdder_68 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_67 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_67;

architecture SYN_full_adder_arch of FullAdder_67 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_66 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_66;

architecture SYN_full_adder_arch of FullAdder_66 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_65 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_65;

architecture SYN_full_adder_arch of FullAdder_65 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_64 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_64;

architecture SYN_full_adder_arch of FullAdder_64 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_63 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_63;

architecture SYN_full_adder_arch of FullAdder_63 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_62 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_62;

architecture SYN_full_adder_arch of FullAdder_62 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_61 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_61;

architecture SYN_full_adder_arch of FullAdder_61 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_60 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_60;

architecture SYN_full_adder_arch of FullAdder_60 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_59 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_59;

architecture SYN_full_adder_arch of FullAdder_59 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_58 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_58;

architecture SYN_full_adder_arch of FullAdder_58 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_57 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_57;

architecture SYN_full_adder_arch of FullAdder_57 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_56 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_56;

architecture SYN_full_adder_arch of FullAdder_56 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_55 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_55;

architecture SYN_full_adder_arch of FullAdder_55 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_54 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_54;

architecture SYN_full_adder_arch of FullAdder_54 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_53 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_53;

architecture SYN_full_adder_arch of FullAdder_53 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_52 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_52;

architecture SYN_full_adder_arch of FullAdder_52 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_51 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_51;

architecture SYN_full_adder_arch of FullAdder_51 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_50 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_50;

architecture SYN_full_adder_arch of FullAdder_50 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_49 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_49;

architecture SYN_full_adder_arch of FullAdder_49 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_48 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_48;

architecture SYN_full_adder_arch of FullAdder_48 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_47 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_47;

architecture SYN_full_adder_arch of FullAdder_47 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_46 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_46;

architecture SYN_full_adder_arch of FullAdder_46 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_45 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_45;

architecture SYN_full_adder_arch of FullAdder_45 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_44 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_44;

architecture SYN_full_adder_arch of FullAdder_44 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_43 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_43;

architecture SYN_full_adder_arch of FullAdder_43 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_42 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_42;

architecture SYN_full_adder_arch of FullAdder_42 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_41 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_41;

architecture SYN_full_adder_arch of FullAdder_41 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_40 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_40;

architecture SYN_full_adder_arch of FullAdder_40 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_39 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_39;

architecture SYN_full_adder_arch of FullAdder_39 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_38 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_38;

architecture SYN_full_adder_arch of FullAdder_38 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_37 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_37;

architecture SYN_full_adder_arch of FullAdder_37 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_36 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_36;

architecture SYN_full_adder_arch of FullAdder_36 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_35 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_35;

architecture SYN_full_adder_arch of FullAdder_35 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_34 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_34;

architecture SYN_full_adder_arch of FullAdder_34 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_33 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_33;

architecture SYN_full_adder_arch of FullAdder_33 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_32 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_32;

architecture SYN_full_adder_arch of FullAdder_32 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_31 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_31;

architecture SYN_full_adder_arch of FullAdder_31 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_30 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_30;

architecture SYN_full_adder_arch of FullAdder_30 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_29 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_29;

architecture SYN_full_adder_arch of FullAdder_29 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_28 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_28;

architecture SYN_full_adder_arch of FullAdder_28 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_27 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_27;

architecture SYN_full_adder_arch of FullAdder_27 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_26 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_26;

architecture SYN_full_adder_arch of FullAdder_26 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_25 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_25;

architecture SYN_full_adder_arch of FullAdder_25 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_24 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_24;

architecture SYN_full_adder_arch of FullAdder_24 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_23 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_23;

architecture SYN_full_adder_arch of FullAdder_23 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_22 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_22;

architecture SYN_full_adder_arch of FullAdder_22 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_21 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_21;

architecture SYN_full_adder_arch of FullAdder_21 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_20 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_20;

architecture SYN_full_adder_arch of FullAdder_20 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_19 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_19;

architecture SYN_full_adder_arch of FullAdder_19 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_18 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_18;

architecture SYN_full_adder_arch of FullAdder_18 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_17 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_17;

architecture SYN_full_adder_arch of FullAdder_17 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_16 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_16;

architecture SYN_full_adder_arch of FullAdder_16 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_15 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_15;

architecture SYN_full_adder_arch of FullAdder_15 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_14 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_14;

architecture SYN_full_adder_arch of FullAdder_14 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_13 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_13;

architecture SYN_full_adder_arch of FullAdder_13 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_12 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_12;

architecture SYN_full_adder_arch of FullAdder_12 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_11 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_11;

architecture SYN_full_adder_arch of FullAdder_11 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_10 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_10;

architecture SYN_full_adder_arch of FullAdder_10 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_9 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_9;

architecture SYN_full_adder_arch of FullAdder_9 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_8 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_8;

architecture SYN_full_adder_arch of FullAdder_8 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_7 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_7;

architecture SYN_full_adder_arch of FullAdder_7 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_6 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_6;

architecture SYN_full_adder_arch of FullAdder_6 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_5 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_5;

architecture SYN_full_adder_arch of FullAdder_5 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_4 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_4;

architecture SYN_full_adder_arch of FullAdder_4 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_3 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_3;

architecture SYN_full_adder_arch of FullAdder_3 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_2 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_2;

architecture SYN_full_adder_arch of FullAdder_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_1 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_1;

architecture SYN_full_adder_arch of FullAdder_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_83 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_83;

architecture SYN_mux_arch of Mux_DATA_SIZE4_83 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_82 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_82;

architecture SYN_mux_arch of Mux_DATA_SIZE4_82 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_81 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_81;

architecture SYN_mux_arch of Mux_DATA_SIZE4_81 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_80 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_80;

architecture SYN_mux_arch of Mux_DATA_SIZE4_80 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_79 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_79;

architecture SYN_mux_arch of Mux_DATA_SIZE4_79 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_78 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_78;

architecture SYN_mux_arch of Mux_DATA_SIZE4_78 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_77 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_77;

architecture SYN_mux_arch of Mux_DATA_SIZE4_77 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_76 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_76;

architecture SYN_mux_arch of Mux_DATA_SIZE4_76 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_75 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_75;

architecture SYN_mux_arch of Mux_DATA_SIZE4_75 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_74 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_74;

architecture SYN_mux_arch of Mux_DATA_SIZE4_74 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_73 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_73;

architecture SYN_mux_arch of Mux_DATA_SIZE4_73 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_72 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_72;

architecture SYN_mux_arch of Mux_DATA_SIZE4_72 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_71 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_71;

architecture SYN_mux_arch of Mux_DATA_SIZE4_71 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_70 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_70;

architecture SYN_mux_arch of Mux_DATA_SIZE4_70 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_69 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_69;

architecture SYN_mux_arch of Mux_DATA_SIZE4_69 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_68 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_68;

architecture SYN_mux_arch of Mux_DATA_SIZE4_68 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_67 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_67;

architecture SYN_mux_arch of Mux_DATA_SIZE4_67 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_66 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_66;

architecture SYN_mux_arch of Mux_DATA_SIZE4_66 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_65 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_65;

architecture SYN_mux_arch of Mux_DATA_SIZE4_65 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_64 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_64;

architecture SYN_mux_arch of Mux_DATA_SIZE4_64 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_63 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_63;

architecture SYN_mux_arch of Mux_DATA_SIZE4_63 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_62 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_62;

architecture SYN_mux_arch of Mux_DATA_SIZE4_62 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_61 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_61;

architecture SYN_mux_arch of Mux_DATA_SIZE4_61 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_60 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_60;

architecture SYN_mux_arch of Mux_DATA_SIZE4_60 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_59 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_59;

architecture SYN_mux_arch of Mux_DATA_SIZE4_59 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_58 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_58;

architecture SYN_mux_arch of Mux_DATA_SIZE4_58 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_57 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_57;

architecture SYN_mux_arch of Mux_DATA_SIZE4_57 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_56 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_56;

architecture SYN_mux_arch of Mux_DATA_SIZE4_56 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_55 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_55;

architecture SYN_mux_arch of Mux_DATA_SIZE4_55 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_54 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_54;

architecture SYN_mux_arch of Mux_DATA_SIZE4_54 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_53 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_53;

architecture SYN_mux_arch of Mux_DATA_SIZE4_53 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_52 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_52;

architecture SYN_mux_arch of Mux_DATA_SIZE4_52 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_51 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_51;

architecture SYN_mux_arch of Mux_DATA_SIZE4_51 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_50 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_50;

architecture SYN_mux_arch of Mux_DATA_SIZE4_50 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_49 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_49;

architecture SYN_mux_arch of Mux_DATA_SIZE4_49 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_48 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_48;

architecture SYN_mux_arch of Mux_DATA_SIZE4_48 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_47 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_47;

architecture SYN_mux_arch of Mux_DATA_SIZE4_47 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_46 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_46;

architecture SYN_mux_arch of Mux_DATA_SIZE4_46 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_45 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_45;

architecture SYN_mux_arch of Mux_DATA_SIZE4_45 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_44 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_44;

architecture SYN_mux_arch of Mux_DATA_SIZE4_44 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_43 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_43;

architecture SYN_mux_arch of Mux_DATA_SIZE4_43 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_42 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_42;

architecture SYN_mux_arch of Mux_DATA_SIZE4_42 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_41 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_41;

architecture SYN_mux_arch of Mux_DATA_SIZE4_41 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_40 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_40;

architecture SYN_mux_arch of Mux_DATA_SIZE4_40 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_39 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_39;

architecture SYN_mux_arch of Mux_DATA_SIZE4_39 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_38 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_38;

architecture SYN_mux_arch of Mux_DATA_SIZE4_38 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_37 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_37;

architecture SYN_mux_arch of Mux_DATA_SIZE4_37 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_36 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_36;

architecture SYN_mux_arch of Mux_DATA_SIZE4_36 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_35 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_35;

architecture SYN_mux_arch of Mux_DATA_SIZE4_35 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_34 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_34;

architecture SYN_mux_arch of Mux_DATA_SIZE4_34 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_33 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_33;

architecture SYN_mux_arch of Mux_DATA_SIZE4_33 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_32 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_32;

architecture SYN_mux_arch of Mux_DATA_SIZE4_32 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_31 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_31;

architecture SYN_mux_arch of Mux_DATA_SIZE4_31 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_30 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_30;

architecture SYN_mux_arch of Mux_DATA_SIZE4_30 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_29 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_29;

architecture SYN_mux_arch of Mux_DATA_SIZE4_29 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_28 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_28;

architecture SYN_mux_arch of Mux_DATA_SIZE4_28 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_27 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_27;

architecture SYN_mux_arch of Mux_DATA_SIZE4_27 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_26 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_26;

architecture SYN_mux_arch of Mux_DATA_SIZE4_26 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_25 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_25;

architecture SYN_mux_arch of Mux_DATA_SIZE4_25 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_24 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_24;

architecture SYN_mux_arch of Mux_DATA_SIZE4_24 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_23 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_23;

architecture SYN_mux_arch of Mux_DATA_SIZE4_23 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_22 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_22;

architecture SYN_mux_arch of Mux_DATA_SIZE4_22 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_21 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_21;

architecture SYN_mux_arch of Mux_DATA_SIZE4_21 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_20 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_20;

architecture SYN_mux_arch of Mux_DATA_SIZE4_20 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_19 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_19;

architecture SYN_mux_arch of Mux_DATA_SIZE4_19 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_18 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_18;

architecture SYN_mux_arch of Mux_DATA_SIZE4_18 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_17 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_17;

architecture SYN_mux_arch of Mux_DATA_SIZE4_17 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_16 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_16;

architecture SYN_mux_arch of Mux_DATA_SIZE4_16 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_15 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_15;

architecture SYN_mux_arch of Mux_DATA_SIZE4_15 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_14 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_14;

architecture SYN_mux_arch of Mux_DATA_SIZE4_14 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_13 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_13;

architecture SYN_mux_arch of Mux_DATA_SIZE4_13 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_12 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_12;

architecture SYN_mux_arch of Mux_DATA_SIZE4_12 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_11 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_11;

architecture SYN_mux_arch of Mux_DATA_SIZE4_11 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_10 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_10;

architecture SYN_mux_arch of Mux_DATA_SIZE4_10 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_9 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_9;

architecture SYN_mux_arch of Mux_DATA_SIZE4_9 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_8 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_8;

architecture SYN_mux_arch of Mux_DATA_SIZE4_8 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_7 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_7;

architecture SYN_mux_arch of Mux_DATA_SIZE4_7 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_6 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_6;

architecture SYN_mux_arch of Mux_DATA_SIZE4_6 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_5 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_5;

architecture SYN_mux_arch of Mux_DATA_SIZE4_5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_4 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_4;

architecture SYN_mux_arch of Mux_DATA_SIZE4_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_3 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_3;

architecture SYN_mux_arch of Mux_DATA_SIZE4_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_2 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_2;

architecture SYN_mux_arch of Mux_DATA_SIZE4_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_1 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_1;

architecture SYN_mux_arch of Mux_DATA_SIZE4_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_167 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_167;

architecture SYN_rca_arch of Rca_DATA_SIZE4_167 is

   component FullAdder_665
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_666
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_667
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_668
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_668 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_667 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_666 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_665 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_166 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_166;

architecture SYN_rca_arch of Rca_DATA_SIZE4_166 is

   component FullAdder_661
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_662
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_663
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_664
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_664 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_663 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_662 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_661 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_165 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_165;

architecture SYN_rca_arch of Rca_DATA_SIZE4_165 is

   component FullAdder_657
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_658
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_659
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_660
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_660 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_659 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_658 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_657 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_164 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_164;

architecture SYN_rca_arch of Rca_DATA_SIZE4_164 is

   component FullAdder_653
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_654
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_655
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_656
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_656 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_655 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_654 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_653 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_163 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_163;

architecture SYN_rca_arch of Rca_DATA_SIZE4_163 is

   component FullAdder_649
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_650
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_651
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_652
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_652 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_651 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_650 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_649 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_162 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_162;

architecture SYN_rca_arch of Rca_DATA_SIZE4_162 is

   component FullAdder_645
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_646
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_647
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_648
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_648 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_647 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_646 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_645 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_161 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_161;

architecture SYN_rca_arch of Rca_DATA_SIZE4_161 is

   component FullAdder_641
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_642
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_643
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_644
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_644 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_643 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_642 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_641 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_160 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_160;

architecture SYN_rca_arch of Rca_DATA_SIZE4_160 is

   component FullAdder_637
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_638
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_639
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_640
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_640 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_639 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_638 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_637 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_159 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_159;

architecture SYN_rca_arch of Rca_DATA_SIZE4_159 is

   component FullAdder_633
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_634
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_635
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_636
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_636 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_635 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_634 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_633 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_158 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_158;

architecture SYN_rca_arch of Rca_DATA_SIZE4_158 is

   component FullAdder_629
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_630
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_631
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_632
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_632 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_631 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_630 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_629 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_157 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_157;

architecture SYN_rca_arch of Rca_DATA_SIZE4_157 is

   component FullAdder_625
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_626
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_627
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_628
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_628 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_627 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_626 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_625 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_156 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_156;

architecture SYN_rca_arch of Rca_DATA_SIZE4_156 is

   component FullAdder_621
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_622
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_623
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_624
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_624 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_623 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_622 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_621 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_155 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_155;

architecture SYN_rca_arch of Rca_DATA_SIZE4_155 is

   component FullAdder_617
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_618
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_619
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_620
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_620 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_619 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_618 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_617 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_154 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_154;

architecture SYN_rca_arch of Rca_DATA_SIZE4_154 is

   component FullAdder_613
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_614
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_615
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_616
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_616 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_615 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_614 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_613 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_153 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_153;

architecture SYN_rca_arch of Rca_DATA_SIZE4_153 is

   component FullAdder_609
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_610
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_611
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_612
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_612 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_611 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_610 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_609 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_152 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_152;

architecture SYN_rca_arch of Rca_DATA_SIZE4_152 is

   component FullAdder_605
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_606
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_607
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_608
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_608 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_607 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_606 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_605 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_151 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_151;

architecture SYN_rca_arch of Rca_DATA_SIZE4_151 is

   component FullAdder_601
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_602
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_603
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_604
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_604 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_603 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_602 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_601 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_150 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_150;

architecture SYN_rca_arch of Rca_DATA_SIZE4_150 is

   component FullAdder_597
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_598
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_599
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_600
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_600 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_599 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_598 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_597 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_149 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_149;

architecture SYN_rca_arch of Rca_DATA_SIZE4_149 is

   component FullAdder_593
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_594
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_595
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_596
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_596 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_595 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_594 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_593 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_148 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_148;

architecture SYN_rca_arch of Rca_DATA_SIZE4_148 is

   component FullAdder_589
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_590
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_591
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_592
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_592 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_591 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_590 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_589 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_147 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_147;

architecture SYN_rca_arch of Rca_DATA_SIZE4_147 is

   component FullAdder_585
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_586
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_587
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_588
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_588 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_587 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_586 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_585 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_146 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_146;

architecture SYN_rca_arch of Rca_DATA_SIZE4_146 is

   component FullAdder_581
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_582
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_583
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_584
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_584 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_583 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_582 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_581 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_145 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_145;

architecture SYN_rca_arch of Rca_DATA_SIZE4_145 is

   component FullAdder_577
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_578
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_579
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_580
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_580 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_579 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_578 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_577 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_144 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_144;

architecture SYN_rca_arch of Rca_DATA_SIZE4_144 is

   component FullAdder_573
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_574
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_575
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_576
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_576 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_575 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_574 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_573 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_143 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_143;

architecture SYN_rca_arch of Rca_DATA_SIZE4_143 is

   component FullAdder_569
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_570
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_571
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_572
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_572 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_571 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_570 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_569 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_142 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_142;

architecture SYN_rca_arch of Rca_DATA_SIZE4_142 is

   component FullAdder_565
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_566
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_567
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_568
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_568 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_567 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_566 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_565 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_141 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_141;

architecture SYN_rca_arch of Rca_DATA_SIZE4_141 is

   component FullAdder_561
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_562
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_563
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_564
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_564 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_563 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_562 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_561 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_140 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_140;

architecture SYN_rca_arch of Rca_DATA_SIZE4_140 is

   component FullAdder_557
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_558
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_559
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_560
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_560 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_559 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_558 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_557 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_139 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_139;

architecture SYN_rca_arch of Rca_DATA_SIZE4_139 is

   component FullAdder_553
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_554
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_555
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_556
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_556 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_555 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_554 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_553 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_138 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_138;

architecture SYN_rca_arch of Rca_DATA_SIZE4_138 is

   component FullAdder_549
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_550
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_551
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_552
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_552 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_551 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_550 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_549 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_137 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_137;

architecture SYN_rca_arch of Rca_DATA_SIZE4_137 is

   component FullAdder_545
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_546
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_547
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_548
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_548 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_547 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_546 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_545 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_136 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_136;

architecture SYN_rca_arch of Rca_DATA_SIZE4_136 is

   component FullAdder_541
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_542
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_543
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_544
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_544 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_543 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_542 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_541 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_135 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_135;

architecture SYN_rca_arch of Rca_DATA_SIZE4_135 is

   component FullAdder_537
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_538
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_539
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_540
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_540 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_539 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_538 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_537 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_134 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_134;

architecture SYN_rca_arch of Rca_DATA_SIZE4_134 is

   component FullAdder_533
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_534
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_535
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_536
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_536 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_535 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_534 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_533 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_133 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_133;

architecture SYN_rca_arch of Rca_DATA_SIZE4_133 is

   component FullAdder_529
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_530
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_531
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_532
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_532 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_531 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_530 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_529 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_132 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_132;

architecture SYN_rca_arch of Rca_DATA_SIZE4_132 is

   component FullAdder_525
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_526
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_527
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_528
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_528 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_527 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_526 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_525 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_131 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_131;

architecture SYN_rca_arch of Rca_DATA_SIZE4_131 is

   component FullAdder_521
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_522
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_523
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_524
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_524 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_523 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_522 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_521 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_130 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_130;

architecture SYN_rca_arch of Rca_DATA_SIZE4_130 is

   component FullAdder_517
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_518
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_519
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_520
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_520 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_519 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_518 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_517 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_129 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_129;

architecture SYN_rca_arch of Rca_DATA_SIZE4_129 is

   component FullAdder_513
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_514
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_515
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_516
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_516 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_515 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_514 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_513 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_128 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_128;

architecture SYN_rca_arch of Rca_DATA_SIZE4_128 is

   component FullAdder_509
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_510
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_511
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_512
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_512 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_511 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_510 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_509 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_127 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_127;

architecture SYN_rca_arch of Rca_DATA_SIZE4_127 is

   component FullAdder_505
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_506
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_507
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_508
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_508 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_507 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_506 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_505 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_126 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_126;

architecture SYN_rca_arch of Rca_DATA_SIZE4_126 is

   component FullAdder_501
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_502
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_503
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_504
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_504 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_503 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_502 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_501 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_125 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_125;

architecture SYN_rca_arch of Rca_DATA_SIZE4_125 is

   component FullAdder_497
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_498
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_499
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_500
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_500 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_499 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_498 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_497 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_124 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_124;

architecture SYN_rca_arch of Rca_DATA_SIZE4_124 is

   component FullAdder_493
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_494
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_495
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_496
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_496 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_495 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_494 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_493 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_123 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_123;

architecture SYN_rca_arch of Rca_DATA_SIZE4_123 is

   component FullAdder_489
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_490
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_491
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_492
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_492 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_491 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_490 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_489 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_122 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_122;

architecture SYN_rca_arch of Rca_DATA_SIZE4_122 is

   component FullAdder_485
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_486
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_487
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_488
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_488 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_487 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_486 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_485 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_121 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_121;

architecture SYN_rca_arch of Rca_DATA_SIZE4_121 is

   component FullAdder_481
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_482
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_483
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_484
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_484 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_483 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_482 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_481 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_120 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_120;

architecture SYN_rca_arch of Rca_DATA_SIZE4_120 is

   component FullAdder_477
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_478
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_479
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_480
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_480 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_479 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_478 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_477 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_119 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_119;

architecture SYN_rca_arch of Rca_DATA_SIZE4_119 is

   component FullAdder_473
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_474
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_475
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_476
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_476 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_475 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_474 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_473 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_118 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_118;

architecture SYN_rca_arch of Rca_DATA_SIZE4_118 is

   component FullAdder_469
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_470
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_471
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_472
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_472 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_471 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_470 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_469 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_117 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_117;

architecture SYN_rca_arch of Rca_DATA_SIZE4_117 is

   component FullAdder_465
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_466
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_467
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_468
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_468 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_467 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_466 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_465 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_116 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_116;

architecture SYN_rca_arch of Rca_DATA_SIZE4_116 is

   component FullAdder_461
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_462
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_463
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_464
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_464 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_463 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_462 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_461 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_115 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_115;

architecture SYN_rca_arch of Rca_DATA_SIZE4_115 is

   component FullAdder_457
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_458
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_459
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_460
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_460 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_459 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_458 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_457 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_114 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_114;

architecture SYN_rca_arch of Rca_DATA_SIZE4_114 is

   component FullAdder_453
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_454
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_455
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_456
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_456 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_455 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_454 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_453 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_113 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_113;

architecture SYN_rca_arch of Rca_DATA_SIZE4_113 is

   component FullAdder_449
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_450
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_451
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_452
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_452 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_451 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_450 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_449 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_112 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_112;

architecture SYN_rca_arch of Rca_DATA_SIZE4_112 is

   component FullAdder_445
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_446
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_447
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_448
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_448 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_447 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_446 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_445 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_111 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_111;

architecture SYN_rca_arch of Rca_DATA_SIZE4_111 is

   component FullAdder_441
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_442
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_443
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_444
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_444 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_443 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_442 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_441 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_110 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_110;

architecture SYN_rca_arch of Rca_DATA_SIZE4_110 is

   component FullAdder_437
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_438
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_439
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_440
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_440 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_439 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_438 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_437 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_109 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_109;

architecture SYN_rca_arch of Rca_DATA_SIZE4_109 is

   component FullAdder_433
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_434
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_435
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_436
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_436 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_435 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_434 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_433 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_108 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_108;

architecture SYN_rca_arch of Rca_DATA_SIZE4_108 is

   component FullAdder_429
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_430
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_431
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_432
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_432 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_431 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_430 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_429 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_107 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_107;

architecture SYN_rca_arch of Rca_DATA_SIZE4_107 is

   component FullAdder_425
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_426
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_427
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_428
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_428 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_427 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_426 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_425 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_106 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_106;

architecture SYN_rca_arch of Rca_DATA_SIZE4_106 is

   component FullAdder_421
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_422
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_423
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_424
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_424 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_423 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_422 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_421 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_105 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_105;

architecture SYN_rca_arch of Rca_DATA_SIZE4_105 is

   component FullAdder_417
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_418
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_419
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_420
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_420 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_419 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_418 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_417 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_104 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_104;

architecture SYN_rca_arch of Rca_DATA_SIZE4_104 is

   component FullAdder_413
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_414
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_415
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_416
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_416 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_415 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_414 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_413 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_103 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_103;

architecture SYN_rca_arch of Rca_DATA_SIZE4_103 is

   component FullAdder_409
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_410
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_411
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_412
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_412 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_411 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_410 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_409 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_102 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_102;

architecture SYN_rca_arch of Rca_DATA_SIZE4_102 is

   component FullAdder_405
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_406
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_407
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_408
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_408 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_407 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_406 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_405 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_101 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_101;

architecture SYN_rca_arch of Rca_DATA_SIZE4_101 is

   component FullAdder_401
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_402
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_403
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_404
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_404 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_403 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_402 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_401 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_100 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_100;

architecture SYN_rca_arch of Rca_DATA_SIZE4_100 is

   component FullAdder_397
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_398
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_399
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_400
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_400 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_399 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_398 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_397 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_99 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_99;

architecture SYN_rca_arch of Rca_DATA_SIZE4_99 is

   component FullAdder_393
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_394
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_395
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_396
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_396 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_395 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_394 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_393 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_98 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_98;

architecture SYN_rca_arch of Rca_DATA_SIZE4_98 is

   component FullAdder_389
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_390
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_391
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_392
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_392 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_391 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_390 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_389 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_97 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_97;

architecture SYN_rca_arch of Rca_DATA_SIZE4_97 is

   component FullAdder_385
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_386
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_387
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_388
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_388 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_387 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_386 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_385 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_96 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_96;

architecture SYN_rca_arch of Rca_DATA_SIZE4_96 is

   component FullAdder_381
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_382
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_383
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_384
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_384 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_383 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_382 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_381 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_95 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_95;

architecture SYN_rca_arch of Rca_DATA_SIZE4_95 is

   component FullAdder_377
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_378
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_379
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_380
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_380 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_379 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_378 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_377 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_94 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_94;

architecture SYN_rca_arch of Rca_DATA_SIZE4_94 is

   component FullAdder_373
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_374
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_375
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_376
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_376 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_375 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_374 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_373 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_93 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_93;

architecture SYN_rca_arch of Rca_DATA_SIZE4_93 is

   component FullAdder_369
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_370
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_371
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_372
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_372 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_371 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_370 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_369 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_92 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_92;

architecture SYN_rca_arch of Rca_DATA_SIZE4_92 is

   component FullAdder_365
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_366
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_367
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_368
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_368 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_367 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_366 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_365 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_91 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_91;

architecture SYN_rca_arch of Rca_DATA_SIZE4_91 is

   component FullAdder_361
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_362
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_363
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_364
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_364 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_363 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_362 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_361 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_90 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_90;

architecture SYN_rca_arch of Rca_DATA_SIZE4_90 is

   component FullAdder_357
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_358
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_359
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_360
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_360 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_359 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_358 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_357 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_89 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_89;

architecture SYN_rca_arch of Rca_DATA_SIZE4_89 is

   component FullAdder_353
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_354
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_355
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_356
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_356 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_355 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_354 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_353 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_88 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_88;

architecture SYN_rca_arch of Rca_DATA_SIZE4_88 is

   component FullAdder_349
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_350
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_351
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_352
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_352 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_351 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_350 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_349 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_87 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_87;

architecture SYN_rca_arch of Rca_DATA_SIZE4_87 is

   component FullAdder_345
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_346
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_347
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_348
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_348 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_347 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_346 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_345 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_86 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_86;

architecture SYN_rca_arch of Rca_DATA_SIZE4_86 is

   component FullAdder_341
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_342
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_343
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_344
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_344 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_343 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_342 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_341 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_85 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_85;

architecture SYN_rca_arch of Rca_DATA_SIZE4_85 is

   component FullAdder_337
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_338
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_339
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_340
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_340 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_339 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_338 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_337 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_84 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_84;

architecture SYN_rca_arch of Rca_DATA_SIZE4_84 is

   component FullAdder_333
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_334
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_335
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_336
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_336 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_335 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_334 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_333 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_83 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_83;

architecture SYN_rca_arch of Rca_DATA_SIZE4_83 is

   component FullAdder_329
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_330
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_331
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_332
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_332 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_331 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_330 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_329 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_82 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_82;

architecture SYN_rca_arch of Rca_DATA_SIZE4_82 is

   component FullAdder_325
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_326
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_327
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_328
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_328 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_327 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_326 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_325 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_81 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_81;

architecture SYN_rca_arch of Rca_DATA_SIZE4_81 is

   component FullAdder_321
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_322
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_323
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_324
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_324 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_323 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_322 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_321 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_80 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_80;

architecture SYN_rca_arch of Rca_DATA_SIZE4_80 is

   component FullAdder_317
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_318
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_319
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_320
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_320 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_319 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_318 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_317 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_79 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_79;

architecture SYN_rca_arch of Rca_DATA_SIZE4_79 is

   component FullAdder_313
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_314
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_315
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_316
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_316 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_315 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_314 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_313 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_78 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_78;

architecture SYN_rca_arch of Rca_DATA_SIZE4_78 is

   component FullAdder_309
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_310
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_311
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_312
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_312 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_311 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_310 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_309 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_77 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_77;

architecture SYN_rca_arch of Rca_DATA_SIZE4_77 is

   component FullAdder_305
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_306
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_307
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_308
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_308 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_307 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_306 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_305 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_76 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_76;

architecture SYN_rca_arch of Rca_DATA_SIZE4_76 is

   component FullAdder_301
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_302
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_303
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_304
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_304 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_303 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_302 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_301 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_75 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_75;

architecture SYN_rca_arch of Rca_DATA_SIZE4_75 is

   component FullAdder_297
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_298
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_299
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_300
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_300 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_299 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_298 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_297 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_74 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_74;

architecture SYN_rca_arch of Rca_DATA_SIZE4_74 is

   component FullAdder_293
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_294
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_295
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_296
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_296 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_295 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_294 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_293 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_73 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_73;

architecture SYN_rca_arch of Rca_DATA_SIZE4_73 is

   component FullAdder_289
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_290
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_291
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_292
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_292 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_291 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_290 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_289 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_72 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_72;

architecture SYN_rca_arch of Rca_DATA_SIZE4_72 is

   component FullAdder_285
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_286
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_287
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_288
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_288 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_287 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_286 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_285 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_71 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_71;

architecture SYN_rca_arch of Rca_DATA_SIZE4_71 is

   component FullAdder_281
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_282
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_283
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_284
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_284 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_283 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_282 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_281 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_70 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_70;

architecture SYN_rca_arch of Rca_DATA_SIZE4_70 is

   component FullAdder_277
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_278
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_279
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_280
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_280 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_279 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_278 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_277 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_69 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_69;

architecture SYN_rca_arch of Rca_DATA_SIZE4_69 is

   component FullAdder_273
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_274
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_275
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_276
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_276 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_275 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_274 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_273 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_68 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_68;

architecture SYN_rca_arch of Rca_DATA_SIZE4_68 is

   component FullAdder_269
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_270
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_271
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_272
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_272 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_271 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_270 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_269 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_67 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_67;

architecture SYN_rca_arch of Rca_DATA_SIZE4_67 is

   component FullAdder_265
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_266
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_267
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_268
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_268 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_267 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_266 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_265 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_66 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_66;

architecture SYN_rca_arch of Rca_DATA_SIZE4_66 is

   component FullAdder_261
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_262
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_263
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_264
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_264 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_263 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_262 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_261 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_65 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_65;

architecture SYN_rca_arch of Rca_DATA_SIZE4_65 is

   component FullAdder_257
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_258
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_259
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_260
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_260 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_259 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_258 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_257 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_64 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_64;

architecture SYN_rca_arch of Rca_DATA_SIZE4_64 is

   component FullAdder_253
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_254
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_255
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_256
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_256 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_255 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_254 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_253 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_63 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_63;

architecture SYN_rca_arch of Rca_DATA_SIZE4_63 is

   component FullAdder_249
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_250
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_251
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_252
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_252 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_251 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_250 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_249 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_62 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_62;

architecture SYN_rca_arch of Rca_DATA_SIZE4_62 is

   component FullAdder_245
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_246
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_247
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_248
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_248 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_247 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_246 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_245 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_61 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_61;

architecture SYN_rca_arch of Rca_DATA_SIZE4_61 is

   component FullAdder_241
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_242
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_243
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_244
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_244 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_243 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_242 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_241 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_60 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_60;

architecture SYN_rca_arch of Rca_DATA_SIZE4_60 is

   component FullAdder_237
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_238
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_239
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_240
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_240 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_239 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_238 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_237 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_59 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_59;

architecture SYN_rca_arch of Rca_DATA_SIZE4_59 is

   component FullAdder_233
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_234
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_235
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_236
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_236 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_235 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_234 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_233 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_58 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_58;

architecture SYN_rca_arch of Rca_DATA_SIZE4_58 is

   component FullAdder_229
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_230
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_231
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_232
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_232 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_231 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_230 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_229 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_57 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_57;

architecture SYN_rca_arch of Rca_DATA_SIZE4_57 is

   component FullAdder_225
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_226
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_227
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_228
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_228 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_227 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_226 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_225 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_56 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_56;

architecture SYN_rca_arch of Rca_DATA_SIZE4_56 is

   component FullAdder_221
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_222
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_223
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_224
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_224 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_223 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_222 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_221 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_55 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_55;

architecture SYN_rca_arch of Rca_DATA_SIZE4_55 is

   component FullAdder_217
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_218
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_219
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_220
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_220 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_219 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_218 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_217 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_54 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_54;

architecture SYN_rca_arch of Rca_DATA_SIZE4_54 is

   component FullAdder_213
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_214
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_215
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_216
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_216 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_215 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_214 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_213 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_53 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_53;

architecture SYN_rca_arch of Rca_DATA_SIZE4_53 is

   component FullAdder_209
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_210
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_211
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_212
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_212 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_211 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_210 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_209 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_52 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_52;

architecture SYN_rca_arch of Rca_DATA_SIZE4_52 is

   component FullAdder_205
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_206
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_207
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_208
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_208 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_207 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_206 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_205 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_51 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_51;

architecture SYN_rca_arch of Rca_DATA_SIZE4_51 is

   component FullAdder_201
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_202
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_203
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_204
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_204 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_203 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_202 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_201 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_50 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_50;

architecture SYN_rca_arch of Rca_DATA_SIZE4_50 is

   component FullAdder_197
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_198
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_199
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_200
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_200 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_199 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_198 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_197 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_49 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_49;

architecture SYN_rca_arch of Rca_DATA_SIZE4_49 is

   component FullAdder_193
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_194
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_195
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_196
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_196 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_195 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_194 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_193 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_48 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_48;

architecture SYN_rca_arch of Rca_DATA_SIZE4_48 is

   component FullAdder_189
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_190
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_191
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_192
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_192 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_191 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_190 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_189 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_47 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_47;

architecture SYN_rca_arch of Rca_DATA_SIZE4_47 is

   component FullAdder_185
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_186
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_187
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_188
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_188 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_187 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_186 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_185 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_46 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_46;

architecture SYN_rca_arch of Rca_DATA_SIZE4_46 is

   component FullAdder_181
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_182
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_183
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_184
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_184 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_183 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_182 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_181 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_45 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_45;

architecture SYN_rca_arch of Rca_DATA_SIZE4_45 is

   component FullAdder_177
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_178
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_179
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_180
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_180 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_179 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_178 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_177 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_44 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_44;

architecture SYN_rca_arch of Rca_DATA_SIZE4_44 is

   component FullAdder_173
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_174
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_175
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_176
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_176 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_175 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_174 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_173 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_43 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_43;

architecture SYN_rca_arch of Rca_DATA_SIZE4_43 is

   component FullAdder_169
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_170
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_171
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_172
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_172 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_171 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_170 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_169 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_42 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_42;

architecture SYN_rca_arch of Rca_DATA_SIZE4_42 is

   component FullAdder_165
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_166
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_167
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_168
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_168 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_167 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_166 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_165 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_41 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_41;

architecture SYN_rca_arch of Rca_DATA_SIZE4_41 is

   component FullAdder_161
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_162
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_163
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_164
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_164 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_163 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_162 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_161 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_40 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_40;

architecture SYN_rca_arch of Rca_DATA_SIZE4_40 is

   component FullAdder_157
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_158
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_159
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_160
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_160 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_159 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_158 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_157 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_39 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_39;

architecture SYN_rca_arch of Rca_DATA_SIZE4_39 is

   component FullAdder_153
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_154
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_155
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_156
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_156 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_155 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_154 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_153 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_38 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_38;

architecture SYN_rca_arch of Rca_DATA_SIZE4_38 is

   component FullAdder_149
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_150
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_151
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_152
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_152 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_151 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_150 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_149 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_37 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_37;

architecture SYN_rca_arch of Rca_DATA_SIZE4_37 is

   component FullAdder_145
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_146
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_147
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_148
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_148 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_147 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_146 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_145 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_36 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_36;

architecture SYN_rca_arch of Rca_DATA_SIZE4_36 is

   component FullAdder_141
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_142
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_143
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_144
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_144 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_143 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_142 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_141 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_35 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_35;

architecture SYN_rca_arch of Rca_DATA_SIZE4_35 is

   component FullAdder_137
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_138
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_139
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_140
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_140 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_139 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_138 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_137 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_34 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_34;

architecture SYN_rca_arch of Rca_DATA_SIZE4_34 is

   component FullAdder_133
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_134
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_135
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_136
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_136 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_135 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_134 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_133 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_33 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_33;

architecture SYN_rca_arch of Rca_DATA_SIZE4_33 is

   component FullAdder_129
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_130
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_131
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_132
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_132 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_131 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_130 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_129 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_32 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_32;

architecture SYN_rca_arch of Rca_DATA_SIZE4_32 is

   component FullAdder_125
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_126
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_127
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_128
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_128 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_127 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_126 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_125 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_31 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_31;

architecture SYN_rca_arch of Rca_DATA_SIZE4_31 is

   component FullAdder_121
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_122
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_123
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_124
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_124 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_123 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_122 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_121 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_30 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_30;

architecture SYN_rca_arch of Rca_DATA_SIZE4_30 is

   component FullAdder_117
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_118
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_119
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_120
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_120 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_119 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_118 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_117 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_29 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_29;

architecture SYN_rca_arch of Rca_DATA_SIZE4_29 is

   component FullAdder_113
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_114
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_115
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_116
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_116 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_115 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_114 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_113 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_28 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_28;

architecture SYN_rca_arch of Rca_DATA_SIZE4_28 is

   component FullAdder_109
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_110
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_111
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_112
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_112 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_111 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_110 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_109 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_27 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_27;

architecture SYN_rca_arch of Rca_DATA_SIZE4_27 is

   component FullAdder_105
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_106
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_107
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_108
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_108 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_107 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_106 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_105 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_26 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_26;

architecture SYN_rca_arch of Rca_DATA_SIZE4_26 is

   component FullAdder_101
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_102
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_103
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_104
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_104 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_103 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_102 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_101 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_25 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_25;

architecture SYN_rca_arch of Rca_DATA_SIZE4_25 is

   component FullAdder_97
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_98
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_99
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_100
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_100 port map( ci => ci, a => a(0), b => b(0), s => s(0), 
                           co => carry_1_port);
   FA3_1 : FullAdder_99 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_98 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_97 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_24 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_24;

architecture SYN_rca_arch of Rca_DATA_SIZE4_24 is

   component FullAdder_93
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_94
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_95
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_96
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_96 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_95 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_94 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_93 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_23 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_23;

architecture SYN_rca_arch of Rca_DATA_SIZE4_23 is

   component FullAdder_89
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_90
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_91
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_92
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_92 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_91 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_90 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_89 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_22 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_22;

architecture SYN_rca_arch of Rca_DATA_SIZE4_22 is

   component FullAdder_85
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_86
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_87
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_88
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_88 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_87 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_86 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_85 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_21 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_21;

architecture SYN_rca_arch of Rca_DATA_SIZE4_21 is

   component FullAdder_81
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_82
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_83
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_84
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_84 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_83 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_82 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_81 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_20 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_20;

architecture SYN_rca_arch of Rca_DATA_SIZE4_20 is

   component FullAdder_77
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_78
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_79
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_80
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_80 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_79 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_78 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_77 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_19 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_19;

architecture SYN_rca_arch of Rca_DATA_SIZE4_19 is

   component FullAdder_73
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_74
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_75
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_76
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_76 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_75 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_74 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_73 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_18 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_18;

architecture SYN_rca_arch of Rca_DATA_SIZE4_18 is

   component FullAdder_69
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_70
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_71
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_72
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_72 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_71 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_70 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_69 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_17 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_17;

architecture SYN_rca_arch of Rca_DATA_SIZE4_17 is

   component FullAdder_65
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_66
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_67
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_68
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_68 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_67 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_66 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_65 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_16 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_16;

architecture SYN_rca_arch of Rca_DATA_SIZE4_16 is

   component FullAdder_61
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_62
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_63
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_64
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_64 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_63 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_62 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_61 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_15 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_15;

architecture SYN_rca_arch of Rca_DATA_SIZE4_15 is

   component FullAdder_57
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_58
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_59
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_60
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_60 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_59 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_58 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_57 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_14 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_14;

architecture SYN_rca_arch of Rca_DATA_SIZE4_14 is

   component FullAdder_53
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_54
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_55
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_56
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_56 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_55 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_54 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_53 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_13 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_13;

architecture SYN_rca_arch of Rca_DATA_SIZE4_13 is

   component FullAdder_49
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_50
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_51
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_52
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_52 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_51 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_50 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_49 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_12 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_12;

architecture SYN_rca_arch of Rca_DATA_SIZE4_12 is

   component FullAdder_45
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_46
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_47
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_48
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_48 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_47 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_46 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_45 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_11 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_11;

architecture SYN_rca_arch of Rca_DATA_SIZE4_11 is

   component FullAdder_41
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_42
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_43
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_44
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_44 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_43 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_42 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_41 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_10 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_10;

architecture SYN_rca_arch of Rca_DATA_SIZE4_10 is

   component FullAdder_37
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_38
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_39
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_40
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_40 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_39 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_38 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_37 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_9 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_9;

architecture SYN_rca_arch of Rca_DATA_SIZE4_9 is

   component FullAdder_33
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_34
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_35
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_36
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_36 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_35 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_34 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_33 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_8 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_8;

architecture SYN_rca_arch of Rca_DATA_SIZE4_8 is

   component FullAdder_29
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_30
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_31
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_32
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_32 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_31 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_30 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_29 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_7 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_7;

architecture SYN_rca_arch of Rca_DATA_SIZE4_7 is

   component FullAdder_25
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_26
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_27
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_28
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_28 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_27 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_26 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_25 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_6 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_6;

architecture SYN_rca_arch of Rca_DATA_SIZE4_6 is

   component FullAdder_21
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_22
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_23
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_24
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_24 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_23 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_22 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_21 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_5 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_5;

architecture SYN_rca_arch of Rca_DATA_SIZE4_5 is

   component FullAdder_17
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_18
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_19
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_20
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_20 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_19 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_18 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_17 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_4 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_4;

architecture SYN_rca_arch of Rca_DATA_SIZE4_4 is

   component FullAdder_13
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_14
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_15
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_16
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_16 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_15 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_14 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_13 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_3 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_3;

architecture SYN_rca_arch of Rca_DATA_SIZE4_3 is

   component FullAdder_9
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_10
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_11
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_12
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_12 port map( ci => ci, a => a(0), b => b(0), s => s(0), co
                           => carry_1_port);
   FA3_1 : FullAdder_11 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_10 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_9 port map( ci => carry_3_port, a => a(3), b => b(3), s =>
                           s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_2 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_2;

architecture SYN_rca_arch of Rca_DATA_SIZE4_2 is

   component FullAdder_5
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_6
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_7
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_8
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_8 port map( ci => ci, a => a(0), b => b(0), s => s(0), co 
                           => carry_1_port);
   FA3_1 : FullAdder_7 port map( ci => carry_1_port, a => a(1), b => b(1), s =>
                           s(1), co => carry_2_port);
   FA3_2 : FullAdder_6 port map( ci => carry_2_port, a => a(2), b => b(2), s =>
                           s(2), co => carry_3_port);
   FA3_3 : FullAdder_5 port map( ci => carry_3_port, a => a(3), b => b(3), s =>
                           s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_1 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_1;

architecture SYN_rca_arch of Rca_DATA_SIZE4_1 is

   component FullAdder_1
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_2
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_3
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_4
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_4 port map( ci => ci, a => a(0), b => b(0), s => s(0), co 
                           => carry_1_port);
   FA3_1 : FullAdder_3 port map( ci => carry_1_port, a => a(1), b => b(1), s =>
                           s(1), co => carry_2_port);
   FA3_2 : FullAdder_2 port map( ci => carry_2_port, a => a(2), b => b(2), s =>
                           s(2), co => carry_3_port);
   FA3_3 : FullAdder_1 port map( ci => carry_3_port, a => a(3), b => b(3), s =>
                           s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_83 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_83;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_83 is

   component Mux_DATA_SIZE4_83
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_165
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_166
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_166 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_165 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_83 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_82 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_82;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_82 is

   component Mux_DATA_SIZE4_82
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_163
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_164
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_164 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_163 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_82 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_81 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_81;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_81 is

   component Mux_DATA_SIZE4_81
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_161
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_162
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_162 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_161 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_81 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_80 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_80;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_80 is

   component Mux_DATA_SIZE4_80
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_159
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_160
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_160 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_159 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_80 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_79 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_79;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_79 is

   component Mux_DATA_SIZE4_79
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_157
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_158
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_158 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_157 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_79 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_78 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_78;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_78 is

   component Mux_DATA_SIZE4_78
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_155
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_156
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_156 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_155 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_78 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_77 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_77;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_77 is

   component Mux_DATA_SIZE4_77
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_153
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_154
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_154 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_153 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_77 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_76 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_76;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_76 is

   component Mux_DATA_SIZE4_76
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_151
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_152
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_152 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_151 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_76 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_75 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_75;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_75 is

   component Mux_DATA_SIZE4_75
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_149
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_150
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_150 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_149 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_75 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_74 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_74;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_74 is

   component Mux_DATA_SIZE4_74
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_147
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_148
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_148 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_147 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_74 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_73 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_73;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_73 is

   component Mux_DATA_SIZE4_73
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_145
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_146
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_146 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_145 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_73 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_72 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_72;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_72 is

   component Mux_DATA_SIZE4_72
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_143
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_144
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_144 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_143 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_72 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_71 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_71;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_71 is

   component Mux_DATA_SIZE4_71
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_141
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_142
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_142 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_141 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_71 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_70 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_70;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_70 is

   component Mux_DATA_SIZE4_70
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_139
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_140
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_140 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_139 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_70 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_69 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_69;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_69 is

   component Mux_DATA_SIZE4_69
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_137
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_138
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_138 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_137 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_69 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_68 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_68;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_68 is

   component Mux_DATA_SIZE4_68
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_135
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_136
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_136 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_135 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_68 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_67 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_67;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_67 is

   component Mux_DATA_SIZE4_67
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_133
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_134
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_134 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_133 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_67 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_66 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_66;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_66 is

   component Mux_DATA_SIZE4_66
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_131
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_132
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_132 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_131 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_66 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_65 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_65;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_65 is

   component Mux_DATA_SIZE4_65
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_129
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_130
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_130 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_129 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_65 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_64 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_64;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_64 is

   component Mux_DATA_SIZE4_64
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_127
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_128
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_128 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_127 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_64 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_63 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_63;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_63 is

   component Mux_DATA_SIZE4_63
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_125
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_126
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_126 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_125 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_63 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_62 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_62;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_62 is

   component Mux_DATA_SIZE4_62
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_123
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_124
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_124 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_123 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_62 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_61 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_61;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_61 is

   component Mux_DATA_SIZE4_61
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_121
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_122
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_122 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_121 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_61 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_60 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_60;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_60 is

   component Mux_DATA_SIZE4_60
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_119
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_120
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_120 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_119 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_60 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_59 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_59;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_59 is

   component Mux_DATA_SIZE4_59
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_117
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_118
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_118 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_117 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_59 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_58 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_58;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_58 is

   component Mux_DATA_SIZE4_58
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_115
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_116
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_116 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_115 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_58 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_57 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_57;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_57 is

   component Mux_DATA_SIZE4_57
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_113
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_114
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_114 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_113 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_57 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_56 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_56;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_56 is

   component Mux_DATA_SIZE4_56
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_111
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_112
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_112 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_111 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_56 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_55 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_55;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_55 is

   component Mux_DATA_SIZE4_55
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_109
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_110
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_110 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_109 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_55 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_54 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_54;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_54 is

   component Mux_DATA_SIZE4_54
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_107
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_108
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_108 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_107 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_54 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_53 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_53;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_53 is

   component Mux_DATA_SIZE4_53
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_105
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_106
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_106 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_105 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_53 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_52 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_52;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_52 is

   component Mux_DATA_SIZE4_52
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_103
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_104
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_104 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_103 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_52 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_51 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_51;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_51 is

   component Mux_DATA_SIZE4_51
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_101
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_102
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_102 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_101 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_51 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_50 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_50;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_50 is

   component Mux_DATA_SIZE4_50
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_99
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_100
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_100 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_99 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_50 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_49 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_49;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_49 is

   component Mux_DATA_SIZE4_49
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_97
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_98
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_98 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_97 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_49 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_48 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_48;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_48 is

   component Mux_DATA_SIZE4_48
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_95
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_96
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_96 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_95 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_48 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_47 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_47;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_47 is

   component Mux_DATA_SIZE4_47
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_93
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_94
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_94 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_93 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_47 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_46 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_46;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_46 is

   component Mux_DATA_SIZE4_46
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_91
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_92
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_92 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_91 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_46 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_45 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_45;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_45 is

   component Mux_DATA_SIZE4_45
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_89
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_90
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_90 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_89 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_45 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_44 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_44;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_44 is

   component Mux_DATA_SIZE4_44
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_87
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_88
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_88 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_87 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_44 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_43 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_43;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_43 is

   component Mux_DATA_SIZE4_43
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_85
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_86
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_86 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_85 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_43 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_42 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_42;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_42 is

   component Mux_DATA_SIZE4_42
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_83
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_84
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_84 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_83 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_42 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_41 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_41;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_41 is

   component Mux_DATA_SIZE4_41
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_81
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_82
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_82 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_81 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_41 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_40 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_40;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_40 is

   component Mux_DATA_SIZE4_40
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_79
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_80
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_80 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_79 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_40 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_39 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_39;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_39 is

   component Mux_DATA_SIZE4_39
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_77
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_78
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_78 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_77 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_39 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_38 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_38;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_38 is

   component Mux_DATA_SIZE4_38
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_75
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_76
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_76 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_75 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_38 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_37 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_37;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_37 is

   component Mux_DATA_SIZE4_37
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_73
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_74
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_74 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_73 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_37 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_36 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_36;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_36 is

   component Mux_DATA_SIZE4_36
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_71
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_72
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_72 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_71 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_36 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_35 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_35;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_35 is

   component Mux_DATA_SIZE4_35
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_69
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_70
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_70 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_69 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_35 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_34 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_34;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_34 is

   component Mux_DATA_SIZE4_34
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_67
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_68
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_68 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_67 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_34 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_33 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_33;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_33 is

   component Mux_DATA_SIZE4_33
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_65
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_66
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_66 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_65 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_33 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_32 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_32;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_32 is

   component Mux_DATA_SIZE4_32
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_63
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_64
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_64 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_63 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_32 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_31 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_31;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_31 is

   component Mux_DATA_SIZE4_31
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_61
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_62
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_62 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_61 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_31 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_30 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_30;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_30 is

   component Mux_DATA_SIZE4_30
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_59
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_60
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_60 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_59 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_30 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_29 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_29;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_29 is

   component Mux_DATA_SIZE4_29
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_57
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_58
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_58 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_57 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_29 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_28 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_28;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_28 is

   component Mux_DATA_SIZE4_28
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_55
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_56
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_56 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_55 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_28 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_27 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_27;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_27 is

   component Mux_DATA_SIZE4_27
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_53
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_54
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_54 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_53 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_27 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_26 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_26;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_26 is

   component Mux_DATA_SIZE4_26
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_51
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_52
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_52 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_51 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_26 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_25 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_25;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_25 is

   component Mux_DATA_SIZE4_25
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_49
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_50
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_50 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_49 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_25 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_24 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_24;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_24 is

   component Mux_DATA_SIZE4_24
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_47
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_48
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_48 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_47 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_24 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_23 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_23;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_23 is

   component Mux_DATA_SIZE4_23
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_45
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_46
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_46 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_45 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_23 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_22 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_22;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_22 is

   component Mux_DATA_SIZE4_22
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_43
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_44
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_44 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_43 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_22 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_21 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_21;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_21 is

   component Mux_DATA_SIZE4_21
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_41
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_42
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_42 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_41 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_21 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_20 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_20;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_20 is

   component Mux_DATA_SIZE4_20
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_39
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_40
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_40 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_39 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_20 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_19 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_19;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_19 is

   component Mux_DATA_SIZE4_19
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_37
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_38
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_38 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_37 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_19 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_18 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_18;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_18 is

   component Mux_DATA_SIZE4_18
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_35
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_36
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_36 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_35 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_18 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_17 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_17;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_17 is

   component Mux_DATA_SIZE4_17
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_33
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_34
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_34 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_33 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_17 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_16 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_16;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_16 is

   component Mux_DATA_SIZE4_16
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_31
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_32
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_32 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_31 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_16 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_15 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_15;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_15 is

   component Mux_DATA_SIZE4_15
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_29
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_30
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_30 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_29 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_15 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_14 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_14;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_14 is

   component Mux_DATA_SIZE4_14
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_27
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_28
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_28 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_27 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_14 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_13 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_13;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_13 is

   component Mux_DATA_SIZE4_13
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_25
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_26
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_26 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_25 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_13 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_12 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_12;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_12 is

   component Mux_DATA_SIZE4_12
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_23
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_24
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_24 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_23 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_12 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_11 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_11;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_11 is

   component Mux_DATA_SIZE4_11
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_21
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_22
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_22 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_21 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_11 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_10 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_10;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_10 is

   component Mux_DATA_SIZE4_10
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_19
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_20
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_20 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_19 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_10 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_9 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_9;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_9 is

   component Mux_DATA_SIZE4_9
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_17
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_18
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_18 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_17 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_9 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_8 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_8;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_8 is

   component Mux_DATA_SIZE4_8
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_15
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_16
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_16 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_15 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_8 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_7 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_7;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_7 is

   component Mux_DATA_SIZE4_7
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_13
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_14
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_14 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_13 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_7 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_6 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_6;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_6 is

   component Mux_DATA_SIZE4_6
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_11
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_12
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_12 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_11 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_6 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_5 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_5;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_5 is

   component Mux_DATA_SIZE4_5
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_9
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_10
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_10 port map( ci => X_Logic0_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_9 port map( ci => X_Logic1_port, a(3) => a(3), a(2) =>
                           a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2)
                           => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_5 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_4 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_4;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_4 is

   component Mux_DATA_SIZE4_4
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_7
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_8
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_8 port map( ci => X_Logic0_port, a(3) => a(3), a(2) =>
                           a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2)
                           => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_7 port map( ci => X_Logic1_port, a(3) => a(3), a(2) =>
                           a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2)
                           => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_4 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_3 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_3;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_3 is

   component Mux_DATA_SIZE4_3
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_5
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_6
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_6 port map( ci => X_Logic0_port, a(3) => a(3), a(2) =>
                           a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2)
                           => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_5 port map( ci => X_Logic1_port, a(3) => a(3), a(2) =>
                           a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2)
                           => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_3 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_2 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_2;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_2 is

   component Mux_DATA_SIZE4_2
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_3
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_4
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_4 port map( ci => X_Logic0_port, a(3) => a(3), a(2) =>
                           a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2)
                           => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_3 port map( ci => X_Logic1_port, a(3) => a(3), a(2) =>
                           a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2)
                           => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_2 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_1 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_1;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_1 is

   component Mux_DATA_SIZE4_1
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_1
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_2
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_2 port map( ci => X_Logic0_port, a(3) => a(3), a(2) =>
                           a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2)
                           => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_1 port map( ci => X_Logic1_port, a(3) => a(3), a(2) =>
                           a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2)
                           => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_1 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderSumGenerator_DATA_SIZE32_SPARSITY4_7 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic_vector 
         (7 downto 0);  sum : out std_logic_vector (31 downto 0));

end AdderSumGenerator_DATA_SIZE32_SPARSITY4_7;

architecture SYN_adder_sum_generator_arch of 
   AdderSumGenerator_DATA_SIZE32_SPARSITY4_7 is

   component AdderCarrySelect_DATA_SIZE4_69
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_70
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_71
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_72
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_73
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_74
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_75
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_76
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;

begin
   
   ACSi_0 : AdderCarrySelect_DATA_SIZE4_76 port map( a(3) => a(3), a(2) => a(2)
                           , a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), sel => cin(0), 
                           sum(3) => sum(3), sum(2) => sum(2), sum(1) => sum(1)
                           , sum(0) => sum(0));
   ACSi_1 : AdderCarrySelect_DATA_SIZE4_75 port map( a(3) => a(7), a(2) => a(6)
                           , a(1) => a(5), a(0) => a(4), b(3) => b(7), b(2) => 
                           b(6), b(1) => b(5), b(0) => b(4), sel => cin(1), 
                           sum(3) => sum(7), sum(2) => sum(6), sum(1) => sum(5)
                           , sum(0) => sum(4));
   ACSi_2 : AdderCarrySelect_DATA_SIZE4_74 port map( a(3) => a(11), a(2) => 
                           a(10), a(1) => a(9), a(0) => a(8), b(3) => b(11), 
                           b(2) => b(10), b(1) => b(9), b(0) => b(8), sel => 
                           cin(2), sum(3) => sum(11), sum(2) => sum(10), sum(1)
                           => sum(9), sum(0) => sum(8));
   ACSi_3 : AdderCarrySelect_DATA_SIZE4_73 port map( a(3) => a(15), a(2) => 
                           a(14), a(1) => a(13), a(0) => a(12), b(3) => b(15), 
                           b(2) => b(14), b(1) => b(13), b(0) => b(12), sel => 
                           cin(3), sum(3) => sum(15), sum(2) => sum(14), sum(1)
                           => sum(13), sum(0) => sum(12));
   ACSi_4 : AdderCarrySelect_DATA_SIZE4_72 port map( a(3) => a(19), a(2) => 
                           a(18), a(1) => a(17), a(0) => a(16), b(3) => b(19), 
                           b(2) => b(18), b(1) => b(17), b(0) => b(16), sel => 
                           cin(4), sum(3) => sum(19), sum(2) => sum(18), sum(1)
                           => sum(17), sum(0) => sum(16));
   ACSi_5 : AdderCarrySelect_DATA_SIZE4_71 port map( a(3) => a(23), a(2) => 
                           a(22), a(1) => a(21), a(0) => a(20), b(3) => b(23), 
                           b(2) => b(22), b(1) => b(21), b(0) => b(20), sel => 
                           cin(5), sum(3) => sum(23), sum(2) => sum(22), sum(1)
                           => sum(21), sum(0) => sum(20));
   ACSi_6 : AdderCarrySelect_DATA_SIZE4_70 port map( a(3) => a(27), a(2) => 
                           a(26), a(1) => a(25), a(0) => a(24), b(3) => b(27), 
                           b(2) => b(26), b(1) => b(25), b(0) => b(24), sel => 
                           cin(6), sum(3) => sum(27), sum(2) => sum(26), sum(1)
                           => sum(25), sum(0) => sum(24));
   ACSi_7 : AdderCarrySelect_DATA_SIZE4_69 port map( a(3) => a(31), a(2) => 
                           a(30), a(1) => a(29), a(0) => a(28), b(3) => b(31), 
                           b(2) => b(30), b(1) => b(29), b(0) => b(28), sel => 
                           cin(7), sum(3) => sum(31), sum(2) => sum(30), sum(1)
                           => sum(29), sum(0) => sum(28));

end SYN_adder_sum_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderSumGenerator_DATA_SIZE32_SPARSITY4_6 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic_vector 
         (7 downto 0);  sum : out std_logic_vector (31 downto 0));

end AdderSumGenerator_DATA_SIZE32_SPARSITY4_6;

architecture SYN_adder_sum_generator_arch of 
   AdderSumGenerator_DATA_SIZE32_SPARSITY4_6 is

   component AdderCarrySelect_DATA_SIZE4_61
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_62
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_63
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_64
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_65
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_66
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_67
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_68
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;

begin
   
   ACSi_0 : AdderCarrySelect_DATA_SIZE4_68 port map( a(3) => a(3), a(2) => a(2)
                           , a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), sel => cin(0), 
                           sum(3) => sum(3), sum(2) => sum(2), sum(1) => sum(1)
                           , sum(0) => sum(0));
   ACSi_1 : AdderCarrySelect_DATA_SIZE4_67 port map( a(3) => a(7), a(2) => a(6)
                           , a(1) => a(5), a(0) => a(4), b(3) => b(7), b(2) => 
                           b(6), b(1) => b(5), b(0) => b(4), sel => cin(1), 
                           sum(3) => sum(7), sum(2) => sum(6), sum(1) => sum(5)
                           , sum(0) => sum(4));
   ACSi_2 : AdderCarrySelect_DATA_SIZE4_66 port map( a(3) => a(11), a(2) => 
                           a(10), a(1) => a(9), a(0) => a(8), b(3) => b(11), 
                           b(2) => b(10), b(1) => b(9), b(0) => b(8), sel => 
                           cin(2), sum(3) => sum(11), sum(2) => sum(10), sum(1)
                           => sum(9), sum(0) => sum(8));
   ACSi_3 : AdderCarrySelect_DATA_SIZE4_65 port map( a(3) => a(15), a(2) => 
                           a(14), a(1) => a(13), a(0) => a(12), b(3) => b(15), 
                           b(2) => b(14), b(1) => b(13), b(0) => b(12), sel => 
                           cin(3), sum(3) => sum(15), sum(2) => sum(14), sum(1)
                           => sum(13), sum(0) => sum(12));
   ACSi_4 : AdderCarrySelect_DATA_SIZE4_64 port map( a(3) => a(19), a(2) => 
                           a(18), a(1) => a(17), a(0) => a(16), b(3) => b(19), 
                           b(2) => b(18), b(1) => b(17), b(0) => b(16), sel => 
                           cin(4), sum(3) => sum(19), sum(2) => sum(18), sum(1)
                           => sum(17), sum(0) => sum(16));
   ACSi_5 : AdderCarrySelect_DATA_SIZE4_63 port map( a(3) => a(23), a(2) => 
                           a(22), a(1) => a(21), a(0) => a(20), b(3) => b(23), 
                           b(2) => b(22), b(1) => b(21), b(0) => b(20), sel => 
                           cin(5), sum(3) => sum(23), sum(2) => sum(22), sum(1)
                           => sum(21), sum(0) => sum(20));
   ACSi_6 : AdderCarrySelect_DATA_SIZE4_62 port map( a(3) => a(27), a(2) => 
                           a(26), a(1) => a(25), a(0) => a(24), b(3) => b(27), 
                           b(2) => b(26), b(1) => b(25), b(0) => b(24), sel => 
                           cin(6), sum(3) => sum(27), sum(2) => sum(26), sum(1)
                           => sum(25), sum(0) => sum(24));
   ACSi_7 : AdderCarrySelect_DATA_SIZE4_61 port map( a(3) => a(31), a(2) => 
                           a(30), a(1) => a(29), a(0) => a(28), b(3) => b(31), 
                           b(2) => b(30), b(1) => b(29), b(0) => b(28), sel => 
                           cin(7), sum(3) => sum(31), sum(2) => sum(30), sum(1)
                           => sum(29), sum(0) => sum(28));

end SYN_adder_sum_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderSumGenerator_DATA_SIZE32_SPARSITY4_5 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic_vector 
         (7 downto 0);  sum : out std_logic_vector (31 downto 0));

end AdderSumGenerator_DATA_SIZE32_SPARSITY4_5;

architecture SYN_adder_sum_generator_arch of 
   AdderSumGenerator_DATA_SIZE32_SPARSITY4_5 is

   component AdderCarrySelect_DATA_SIZE4_49
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_50
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_51
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_52
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_53
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_54
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_55
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_56
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;

begin
   
   ACSi_0 : AdderCarrySelect_DATA_SIZE4_56 port map( a(3) => a(3), a(2) => a(2)
                           , a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), sel => cin(0), 
                           sum(3) => sum(3), sum(2) => sum(2), sum(1) => sum(1)
                           , sum(0) => sum(0));
   ACSi_1 : AdderCarrySelect_DATA_SIZE4_55 port map( a(3) => a(7), a(2) => a(6)
                           , a(1) => a(5), a(0) => a(4), b(3) => b(7), b(2) => 
                           b(6), b(1) => b(5), b(0) => b(4), sel => cin(1), 
                           sum(3) => sum(7), sum(2) => sum(6), sum(1) => sum(5)
                           , sum(0) => sum(4));
   ACSi_2 : AdderCarrySelect_DATA_SIZE4_54 port map( a(3) => a(11), a(2) => 
                           a(10), a(1) => a(9), a(0) => a(8), b(3) => b(11), 
                           b(2) => b(10), b(1) => b(9), b(0) => b(8), sel => 
                           cin(2), sum(3) => sum(11), sum(2) => sum(10), sum(1)
                           => sum(9), sum(0) => sum(8));
   ACSi_3 : AdderCarrySelect_DATA_SIZE4_53 port map( a(3) => a(15), a(2) => 
                           a(14), a(1) => a(13), a(0) => a(12), b(3) => b(15), 
                           b(2) => b(14), b(1) => b(13), b(0) => b(12), sel => 
                           cin(3), sum(3) => sum(15), sum(2) => sum(14), sum(1)
                           => sum(13), sum(0) => sum(12));
   ACSi_4 : AdderCarrySelect_DATA_SIZE4_52 port map( a(3) => a(19), a(2) => 
                           a(18), a(1) => a(17), a(0) => a(16), b(3) => b(19), 
                           b(2) => b(18), b(1) => b(17), b(0) => b(16), sel => 
                           cin(4), sum(3) => sum(19), sum(2) => sum(18), sum(1)
                           => sum(17), sum(0) => sum(16));
   ACSi_5 : AdderCarrySelect_DATA_SIZE4_51 port map( a(3) => a(23), a(2) => 
                           a(22), a(1) => a(21), a(0) => a(20), b(3) => b(23), 
                           b(2) => b(22), b(1) => b(21), b(0) => b(20), sel => 
                           cin(5), sum(3) => sum(23), sum(2) => sum(22), sum(1)
                           => sum(21), sum(0) => sum(20));
   ACSi_6 : AdderCarrySelect_DATA_SIZE4_50 port map( a(3) => a(27), a(2) => 
                           a(26), a(1) => a(25), a(0) => a(24), b(3) => b(27), 
                           b(2) => b(26), b(1) => b(25), b(0) => b(24), sel => 
                           cin(6), sum(3) => sum(27), sum(2) => sum(26), sum(1)
                           => sum(25), sum(0) => sum(24));
   ACSi_7 : AdderCarrySelect_DATA_SIZE4_49 port map( a(3) => a(31), a(2) => 
                           a(30), a(1) => a(29), a(0) => a(28), b(3) => b(31), 
                           b(2) => b(30), b(1) => b(29), b(0) => b(28), sel => 
                           cin(7), sum(3) => sum(31), sum(2) => sum(30), sum(1)
                           => sum(29), sum(0) => sum(28));

end SYN_adder_sum_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderSumGenerator_DATA_SIZE32_SPARSITY4_4 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic_vector 
         (7 downto 0);  sum : out std_logic_vector (31 downto 0));

end AdderSumGenerator_DATA_SIZE32_SPARSITY4_4;

architecture SYN_adder_sum_generator_arch of 
   AdderSumGenerator_DATA_SIZE32_SPARSITY4_4 is

   component AdderCarrySelect_DATA_SIZE4_41
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_42
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_43
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_44
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_45
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_46
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_47
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_48
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;

begin
   
   ACSi_0 : AdderCarrySelect_DATA_SIZE4_48 port map( a(3) => a(3), a(2) => a(2)
                           , a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), sel => cin(0), 
                           sum(3) => sum(3), sum(2) => sum(2), sum(1) => sum(1)
                           , sum(0) => sum(0));
   ACSi_1 : AdderCarrySelect_DATA_SIZE4_47 port map( a(3) => a(7), a(2) => a(6)
                           , a(1) => a(5), a(0) => a(4), b(3) => b(7), b(2) => 
                           b(6), b(1) => b(5), b(0) => b(4), sel => cin(1), 
                           sum(3) => sum(7), sum(2) => sum(6), sum(1) => sum(5)
                           , sum(0) => sum(4));
   ACSi_2 : AdderCarrySelect_DATA_SIZE4_46 port map( a(3) => a(11), a(2) => 
                           a(10), a(1) => a(9), a(0) => a(8), b(3) => b(11), 
                           b(2) => b(10), b(1) => b(9), b(0) => b(8), sel => 
                           cin(2), sum(3) => sum(11), sum(2) => sum(10), sum(1)
                           => sum(9), sum(0) => sum(8));
   ACSi_3 : AdderCarrySelect_DATA_SIZE4_45 port map( a(3) => a(15), a(2) => 
                           a(14), a(1) => a(13), a(0) => a(12), b(3) => b(15), 
                           b(2) => b(14), b(1) => b(13), b(0) => b(12), sel => 
                           cin(3), sum(3) => sum(15), sum(2) => sum(14), sum(1)
                           => sum(13), sum(0) => sum(12));
   ACSi_4 : AdderCarrySelect_DATA_SIZE4_44 port map( a(3) => a(19), a(2) => 
                           a(18), a(1) => a(17), a(0) => a(16), b(3) => b(19), 
                           b(2) => b(18), b(1) => b(17), b(0) => b(16), sel => 
                           cin(4), sum(3) => sum(19), sum(2) => sum(18), sum(1)
                           => sum(17), sum(0) => sum(16));
   ACSi_5 : AdderCarrySelect_DATA_SIZE4_43 port map( a(3) => a(23), a(2) => 
                           a(22), a(1) => a(21), a(0) => a(20), b(3) => b(23), 
                           b(2) => b(22), b(1) => b(21), b(0) => b(20), sel => 
                           cin(5), sum(3) => sum(23), sum(2) => sum(22), sum(1)
                           => sum(21), sum(0) => sum(20));
   ACSi_6 : AdderCarrySelect_DATA_SIZE4_42 port map( a(3) => a(27), a(2) => 
                           a(26), a(1) => a(25), a(0) => a(24), b(3) => b(27), 
                           b(2) => b(26), b(1) => b(25), b(0) => b(24), sel => 
                           cin(6), sum(3) => sum(27), sum(2) => sum(26), sum(1)
                           => sum(25), sum(0) => sum(24));
   ACSi_7 : AdderCarrySelect_DATA_SIZE4_41 port map( a(3) => a(31), a(2) => 
                           a(30), a(1) => a(29), a(0) => a(28), b(3) => b(31), 
                           b(2) => b(30), b(1) => b(29), b(0) => b(28), sel => 
                           cin(7), sum(3) => sum(31), sum(2) => sum(30), sum(1)
                           => sum(29), sum(0) => sum(28));

end SYN_adder_sum_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderSumGenerator_DATA_SIZE32_SPARSITY4_3 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic_vector 
         (7 downto 0);  sum : out std_logic_vector (31 downto 0));

end AdderSumGenerator_DATA_SIZE32_SPARSITY4_3;

architecture SYN_adder_sum_generator_arch of 
   AdderSumGenerator_DATA_SIZE32_SPARSITY4_3 is

   component AdderCarrySelect_DATA_SIZE4_33
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_34
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_35
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_36
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_37
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_38
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_39
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_40
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;

begin
   
   ACSi_0 : AdderCarrySelect_DATA_SIZE4_40 port map( a(3) => a(3), a(2) => a(2)
                           , a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), sel => cin(0), 
                           sum(3) => sum(3), sum(2) => sum(2), sum(1) => sum(1)
                           , sum(0) => sum(0));
   ACSi_1 : AdderCarrySelect_DATA_SIZE4_39 port map( a(3) => a(7), a(2) => a(6)
                           , a(1) => a(5), a(0) => a(4), b(3) => b(7), b(2) => 
                           b(6), b(1) => b(5), b(0) => b(4), sel => cin(1), 
                           sum(3) => sum(7), sum(2) => sum(6), sum(1) => sum(5)
                           , sum(0) => sum(4));
   ACSi_2 : AdderCarrySelect_DATA_SIZE4_38 port map( a(3) => a(11), a(2) => 
                           a(10), a(1) => a(9), a(0) => a(8), b(3) => b(11), 
                           b(2) => b(10), b(1) => b(9), b(0) => b(8), sel => 
                           cin(2), sum(3) => sum(11), sum(2) => sum(10), sum(1)
                           => sum(9), sum(0) => sum(8));
   ACSi_3 : AdderCarrySelect_DATA_SIZE4_37 port map( a(3) => a(15), a(2) => 
                           a(14), a(1) => a(13), a(0) => a(12), b(3) => b(15), 
                           b(2) => b(14), b(1) => b(13), b(0) => b(12), sel => 
                           cin(3), sum(3) => sum(15), sum(2) => sum(14), sum(1)
                           => sum(13), sum(0) => sum(12));
   ACSi_4 : AdderCarrySelect_DATA_SIZE4_36 port map( a(3) => a(19), a(2) => 
                           a(18), a(1) => a(17), a(0) => a(16), b(3) => b(19), 
                           b(2) => b(18), b(1) => b(17), b(0) => b(16), sel => 
                           cin(4), sum(3) => sum(19), sum(2) => sum(18), sum(1)
                           => sum(17), sum(0) => sum(16));
   ACSi_5 : AdderCarrySelect_DATA_SIZE4_35 port map( a(3) => a(23), a(2) => 
                           a(22), a(1) => a(21), a(0) => a(20), b(3) => b(23), 
                           b(2) => b(22), b(1) => b(21), b(0) => b(20), sel => 
                           cin(5), sum(3) => sum(23), sum(2) => sum(22), sum(1)
                           => sum(21), sum(0) => sum(20));
   ACSi_6 : AdderCarrySelect_DATA_SIZE4_34 port map( a(3) => a(27), a(2) => 
                           a(26), a(1) => a(25), a(0) => a(24), b(3) => b(27), 
                           b(2) => b(26), b(1) => b(25), b(0) => b(24), sel => 
                           cin(6), sum(3) => sum(27), sum(2) => sum(26), sum(1)
                           => sum(25), sum(0) => sum(24));
   ACSi_7 : AdderCarrySelect_DATA_SIZE4_33 port map( a(3) => a(31), a(2) => 
                           a(30), a(1) => a(29), a(0) => a(28), b(3) => b(31), 
                           b(2) => b(30), b(1) => b(29), b(0) => b(28), sel => 
                           cin(7), sum(3) => sum(31), sum(2) => sum(30), sum(1)
                           => sum(29), sum(0) => sum(28));

end SYN_adder_sum_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderSumGenerator_DATA_SIZE32_SPARSITY4_2 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic_vector 
         (7 downto 0);  sum : out std_logic_vector (31 downto 0));

end AdderSumGenerator_DATA_SIZE32_SPARSITY4_2;

architecture SYN_adder_sum_generator_arch of 
   AdderSumGenerator_DATA_SIZE32_SPARSITY4_2 is

   component AdderCarrySelect_DATA_SIZE4_9
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_10
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_11
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_12
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_13
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_14
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_15
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_16
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;

begin
   
   ACSi_0 : AdderCarrySelect_DATA_SIZE4_16 port map( a(3) => a(3), a(2) => a(2)
                           , a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), sel => cin(0), 
                           sum(3) => sum(3), sum(2) => sum(2), sum(1) => sum(1)
                           , sum(0) => sum(0));
   ACSi_1 : AdderCarrySelect_DATA_SIZE4_15 port map( a(3) => a(7), a(2) => a(6)
                           , a(1) => a(5), a(0) => a(4), b(3) => b(7), b(2) => 
                           b(6), b(1) => b(5), b(0) => b(4), sel => cin(1), 
                           sum(3) => sum(7), sum(2) => sum(6), sum(1) => sum(5)
                           , sum(0) => sum(4));
   ACSi_2 : AdderCarrySelect_DATA_SIZE4_14 port map( a(3) => a(11), a(2) => 
                           a(10), a(1) => a(9), a(0) => a(8), b(3) => b(11), 
                           b(2) => b(10), b(1) => b(9), b(0) => b(8), sel => 
                           cin(2), sum(3) => sum(11), sum(2) => sum(10), sum(1)
                           => sum(9), sum(0) => sum(8));
   ACSi_3 : AdderCarrySelect_DATA_SIZE4_13 port map( a(3) => a(15), a(2) => 
                           a(14), a(1) => a(13), a(0) => a(12), b(3) => b(15), 
                           b(2) => b(14), b(1) => b(13), b(0) => b(12), sel => 
                           cin(3), sum(3) => sum(15), sum(2) => sum(14), sum(1)
                           => sum(13), sum(0) => sum(12));
   ACSi_4 : AdderCarrySelect_DATA_SIZE4_12 port map( a(3) => a(19), a(2) => 
                           a(18), a(1) => a(17), a(0) => a(16), b(3) => b(19), 
                           b(2) => b(18), b(1) => b(17), b(0) => b(16), sel => 
                           cin(4), sum(3) => sum(19), sum(2) => sum(18), sum(1)
                           => sum(17), sum(0) => sum(16));
   ACSi_5 : AdderCarrySelect_DATA_SIZE4_11 port map( a(3) => a(23), a(2) => 
                           a(22), a(1) => a(21), a(0) => a(20), b(3) => b(23), 
                           b(2) => b(22), b(1) => b(21), b(0) => b(20), sel => 
                           cin(5), sum(3) => sum(23), sum(2) => sum(22), sum(1)
                           => sum(21), sum(0) => sum(20));
   ACSi_6 : AdderCarrySelect_DATA_SIZE4_10 port map( a(3) => a(27), a(2) => 
                           a(26), a(1) => a(25), a(0) => a(24), b(3) => b(27), 
                           b(2) => b(26), b(1) => b(25), b(0) => b(24), sel => 
                           cin(6), sum(3) => sum(27), sum(2) => sum(26), sum(1)
                           => sum(25), sum(0) => sum(24));
   ACSi_7 : AdderCarrySelect_DATA_SIZE4_9 port map( a(3) => a(31), a(2) => 
                           a(30), a(1) => a(29), a(0) => a(28), b(3) => b(31), 
                           b(2) => b(30), b(1) => b(29), b(0) => b(28), sel => 
                           cin(7), sum(3) => sum(31), sum(2) => sum(30), sum(1)
                           => sum(29), sum(0) => sum(28));

end SYN_adder_sum_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderSumGenerator_DATA_SIZE32_SPARSITY4_1 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic_vector 
         (7 downto 0);  sum : out std_logic_vector (31 downto 0));

end AdderSumGenerator_DATA_SIZE32_SPARSITY4_1;

architecture SYN_adder_sum_generator_arch of 
   AdderSumGenerator_DATA_SIZE32_SPARSITY4_1 is

   component AdderCarrySelect_DATA_SIZE4_1
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_2
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_3
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_4
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_5
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_6
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_7
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_8
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;

begin
   
   ACSi_0 : AdderCarrySelect_DATA_SIZE4_8 port map( a(3) => a(3), a(2) => a(2),
                           a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), sel => cin(0), 
                           sum(3) => sum(3), sum(2) => sum(2), sum(1) => sum(1)
                           , sum(0) => sum(0));
   ACSi_1 : AdderCarrySelect_DATA_SIZE4_7 port map( a(3) => a(7), a(2) => a(6),
                           a(1) => a(5), a(0) => a(4), b(3) => b(7), b(2) => 
                           b(6), b(1) => b(5), b(0) => b(4), sel => cin(1), 
                           sum(3) => sum(7), sum(2) => sum(6), sum(1) => sum(5)
                           , sum(0) => sum(4));
   ACSi_2 : AdderCarrySelect_DATA_SIZE4_6 port map( a(3) => a(11), a(2) => 
                           a(10), a(1) => a(9), a(0) => a(8), b(3) => b(11), 
                           b(2) => b(10), b(1) => b(9), b(0) => b(8), sel => 
                           cin(2), sum(3) => sum(11), sum(2) => sum(10), sum(1)
                           => sum(9), sum(0) => sum(8));
   ACSi_3 : AdderCarrySelect_DATA_SIZE4_5 port map( a(3) => a(15), a(2) => 
                           a(14), a(1) => a(13), a(0) => a(12), b(3) => b(15), 
                           b(2) => b(14), b(1) => b(13), b(0) => b(12), sel => 
                           cin(3), sum(3) => sum(15), sum(2) => sum(14), sum(1)
                           => sum(13), sum(0) => sum(12));
   ACSi_4 : AdderCarrySelect_DATA_SIZE4_4 port map( a(3) => a(19), a(2) => 
                           a(18), a(1) => a(17), a(0) => a(16), b(3) => b(19), 
                           b(2) => b(18), b(1) => b(17), b(0) => b(16), sel => 
                           cin(4), sum(3) => sum(19), sum(2) => sum(18), sum(1)
                           => sum(17), sum(0) => sum(16));
   ACSi_5 : AdderCarrySelect_DATA_SIZE4_3 port map( a(3) => a(23), a(2) => 
                           a(22), a(1) => a(21), a(0) => a(20), b(3) => b(23), 
                           b(2) => b(22), b(1) => b(21), b(0) => b(20), sel => 
                           cin(5), sum(3) => sum(23), sum(2) => sum(22), sum(1)
                           => sum(21), sum(0) => sum(20));
   ACSi_6 : AdderCarrySelect_DATA_SIZE4_2 port map( a(3) => a(27), a(2) => 
                           a(26), a(1) => a(25), a(0) => a(24), b(3) => b(27), 
                           b(2) => b(26), b(1) => b(25), b(0) => b(24), sel => 
                           cin(6), sum(3) => sum(27), sum(2) => sum(26), sum(1)
                           => sum(25), sum(0) => sum(24));
   ACSi_7 : AdderCarrySelect_DATA_SIZE4_1 port map( a(3) => a(31), a(2) => 
                           a(30), a(1) => a(29), a(0) => a(28), b(3) => b(31), 
                           b(2) => b(30), b(1) => b(29), b(0) => b(28), sel => 
                           cin(7), sum(3) => sum(31), sum(2) => sum(30), sum(1)
                           => sum(29), sum(0) => sum(28));

end SYN_adder_sum_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4CarryGenerator_DATA_SIZE32_SPARSITY4_7 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  cout :
         out std_logic_vector (7 downto 0));

end P4CarryGenerator_DATA_SIZE32_SPARSITY4_7;

architecture SYN_p4_carry_generator_arch of 
   P4CarryGenerator_DATA_SIZE32_SPARSITY4_7 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal cout_7_port, cout_6_port, cout_5_port, cout_4_port, cout_3_port, 
      cout_2_port, cout_1_port, cout_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9
      , n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, 
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101 : std_logic;

begin
   cout <= ( cout_7_port, cout_6_port, cout_5_port, cout_4_port, cout_3_port, 
      cout_2_port, cout_1_port, cout_0_port );
   
   U1 : OAI22_X1 port map( A1 => n1, A2 => n2, B1 => n3, B2 => n4, ZN => 
                           cout_7_port);
   U2 : AOI22_X1 port map( A1 => b(30), A2 => n5, B1 => a(30), B2 => n6, ZN => 
                           n4);
   U3 : OR2_X1 port map( A1 => n6, A2 => a(30), ZN => n5);
   U4 : OAI21_X1 port map( B1 => n7, B2 => n8, A => n9, ZN => n6);
   U5 : OAI21_X1 port map( B1 => b(29), B2 => a(29), A => n10, ZN => n9);
   U6 : INV_X1 port map( A => n11, ZN => n10);
   U7 : AOI21_X1 port map( B1 => cout_6_port, B2 => a(28), A => n12, ZN => n11)
                           ;
   U8 : INV_X1 port map( A => n13, ZN => n12);
   U9 : OAI21_X1 port map( B1 => a(28), B2 => cout_6_port, A => b(28), ZN => 
                           n13);
   U10 : INV_X1 port map( A => b(29), ZN => n8);
   U11 : INV_X1 port map( A => a(29), ZN => n7);
   U12 : NOR2_X1 port map( A1 => b(31), A2 => a(31), ZN => n3);
   U13 : INV_X1 port map( A => b(31), ZN => n2);
   U14 : INV_X1 port map( A => a(31), ZN => n1);
   U15 : OAI21_X1 port map( B1 => n14, B2 => n15, A => n16, ZN => cout_6_port);
   U16 : OAI21_X1 port map( B1 => a(27), B2 => n17, A => b(27), ZN => n16);
   U17 : INV_X1 port map( A => n14, ZN => n17);
   U18 : INV_X1 port map( A => a(27), ZN => n15);
   U19 : AOI21_X1 port map( B1 => a(26), B2 => b(26), A => n18, ZN => n14);
   U20 : INV_X1 port map( A => n19, ZN => n18);
   U21 : OAI22_X1 port map( A1 => n20, A2 => n21, B1 => a(26), B2 => b(26), ZN 
                           => n19);
   U22 : NOR2_X1 port map( A1 => n22, A2 => n23, ZN => n21);
   U23 : AOI22_X1 port map( A1 => n22, A2 => n23, B1 => n24, B2 => n25, ZN => 
                           n20);
   U24 : OAI21_X1 port map( B1 => a(24), B2 => cout_5_port, A => b(24), ZN => 
                           n25);
   U25 : NAND2_X1 port map( A1 => a(24), A2 => cout_5_port, ZN => n24);
   U26 : INV_X1 port map( A => b(25), ZN => n23);
   U27 : INV_X1 port map( A => a(25), ZN => n22);
   U28 : OAI22_X1 port map( A1 => n26, A2 => n27, B1 => n28, B2 => n29, ZN => 
                           cout_5_port);
   U29 : AOI22_X1 port map( A1 => b(22), A2 => n30, B1 => a(22), B2 => n31, ZN 
                           => n29);
   U30 : OR2_X1 port map( A1 => n31, A2 => a(22), ZN => n30);
   U31 : OAI21_X1 port map( B1 => n32, B2 => n33, A => n34, ZN => n31);
   U32 : OAI21_X1 port map( B1 => b(21), B2 => a(21), A => n35, ZN => n34);
   U33 : OAI21_X1 port map( B1 => n36, B2 => n37, A => n38, ZN => n35);
   U34 : OAI21_X1 port map( B1 => a(20), B2 => cout_4_port, A => b(20), ZN => 
                           n38);
   U35 : INV_X1 port map( A => a(20), ZN => n37);
   U36 : INV_X1 port map( A => cout_4_port, ZN => n36);
   U37 : INV_X1 port map( A => b(21), ZN => n33);
   U38 : INV_X1 port map( A => a(21), ZN => n32);
   U39 : NOR2_X1 port map( A1 => b(23), A2 => a(23), ZN => n28);
   U40 : INV_X1 port map( A => b(23), ZN => n27);
   U41 : INV_X1 port map( A => a(23), ZN => n26);
   U42 : OAI211_X1 port map( C1 => n39, C2 => n40, A => n41, B => n42, ZN => 
                           cout_4_port);
   U43 : OAI211_X1 port map( C1 => b(19), C2 => a(19), A => cout_3_port, B => 
                           n43, ZN => n42);
   U44 : AOI221_X1 port map( B1 => n44, B2 => n45, C1 => n46, C2 => n47, A => 
                           n48, ZN => n43);
   U45 : OAI21_X1 port map( B1 => n49, B2 => a(19), A => b(19), ZN => n41);
   U46 : INV_X1 port map( A => a(19), ZN => n40);
   U47 : INV_X1 port map( A => n49, ZN => n39);
   U48 : AOI21_X1 port map( B1 => n44, B2 => n50, A => n51, ZN => n49);
   U49 : INV_X1 port map( A => n52, ZN => n51);
   U50 : OAI21_X1 port map( B1 => n50, B2 => n44, A => n45, ZN => n52);
   U51 : INV_X1 port map( A => b(18), ZN => n45);
   U52 : AOI21_X1 port map( B1 => a(17), B2 => b(17), A => n53, ZN => n50);
   U53 : NOR3_X1 port map( A1 => n46, A2 => n48, A3 => n47, ZN => n53);
   U54 : INV_X1 port map( A => b(16), ZN => n47);
   U55 : NOR2_X1 port map( A1 => b(17), A2 => a(17), ZN => n48);
   U56 : INV_X1 port map( A => a(16), ZN => n46);
   U57 : INV_X1 port map( A => a(18), ZN => n44);
   U58 : INV_X1 port map( A => n54, ZN => cout_3_port);
   U59 : OAI22_X1 port map( A1 => a(15), A2 => n55, B1 => b(15), B2 => n56, ZN 
                           => n54);
   U60 : AND2_X1 port map( A1 => n55, A2 => a(15), ZN => n56);
   U61 : INV_X1 port map( A => n57, ZN => n55);
   U62 : OAI22_X1 port map( A1 => a(14), A2 => n58, B1 => b(14), B2 => n59, ZN 
                           => n57);
   U63 : AND2_X1 port map( A1 => n58, A2 => a(14), ZN => n59);
   U64 : OAI21_X1 port map( B1 => n60, B2 => n61, A => n62, ZN => n58);
   U65 : OAI21_X1 port map( B1 => b(13), B2 => a(13), A => n63, ZN => n62);
   U66 : INV_X1 port map( A => n64, ZN => n63);
   U67 : AOI21_X1 port map( B1 => cout_2_port, B2 => a(12), A => n65, ZN => n64
                           );
   U68 : INV_X1 port map( A => n66, ZN => n65);
   U69 : OAI21_X1 port map( B1 => a(12), B2 => cout_2_port, A => b(12), ZN => 
                           n66);
   U70 : INV_X1 port map( A => b(13), ZN => n61);
   U71 : INV_X1 port map( A => a(13), ZN => n60);
   U72 : OAI21_X1 port map( B1 => n67, B2 => n68, A => n69, ZN => cout_2_port);
   U73 : OAI21_X1 port map( B1 => a(11), B2 => n70, A => b(11), ZN => n69);
   U74 : INV_X1 port map( A => n67, ZN => n70);
   U75 : INV_X1 port map( A => a(11), ZN => n68);
   U76 : AOI21_X1 port map( B1 => a(10), B2 => b(10), A => n71, ZN => n67);
   U77 : INV_X1 port map( A => n72, ZN => n71);
   U78 : OAI22_X1 port map( A1 => n73, A2 => n74, B1 => a(10), B2 => b(10), ZN 
                           => n72);
   U79 : NOR2_X1 port map( A1 => n75, A2 => n76, ZN => n74);
   U80 : AOI22_X1 port map( A1 => n75, A2 => n76, B1 => n77, B2 => n78, ZN => 
                           n73);
   U81 : OAI21_X1 port map( B1 => a(8), B2 => cout_1_port, A => b(8), ZN => n78
                           );
   U82 : NAND2_X1 port map( A1 => a(8), A2 => cout_1_port, ZN => n77);
   U83 : INV_X1 port map( A => b(9), ZN => n76);
   U84 : INV_X1 port map( A => a(9), ZN => n75);
   U85 : OAI21_X1 port map( B1 => n79, B2 => n80, A => n81, ZN => cout_1_port);
   U86 : OAI21_X1 port map( B1 => b(7), B2 => a(7), A => n82, ZN => n81);
   U87 : OAI21_X1 port map( B1 => n83, B2 => n84, A => n85, ZN => n82);
   U88 : OAI21_X1 port map( B1 => a(6), B2 => n86, A => b(6), ZN => n85);
   U89 : INV_X1 port map( A => n83, ZN => n86);
   U90 : INV_X1 port map( A => a(6), ZN => n84);
   U91 : AOI22_X1 port map( A1 => a(5), A2 => b(5), B1 => n87, B2 => n88, ZN =>
                           n83);
   U92 : INV_X1 port map( A => n89, ZN => n88);
   U93 : AOI22_X1 port map( A1 => b(4), A2 => n90, B1 => a(4), B2 => 
                           cout_0_port, ZN => n89);
   U94 : OR2_X1 port map( A1 => a(4), A2 => cout_0_port, ZN => n90);
   U95 : OR2_X1 port map( A1 => b(5), A2 => a(5), ZN => n87);
   U96 : INV_X1 port map( A => b(7), ZN => n80);
   U97 : INV_X1 port map( A => a(7), ZN => n79);
   U98 : INV_X1 port map( A => n91, ZN => cout_0_port);
   U99 : OAI22_X1 port map( A1 => a(3), A2 => n92, B1 => b(3), B2 => n93, ZN =>
                           n91);
   U100 : AND2_X1 port map( A1 => n92, A2 => a(3), ZN => n93);
   U101 : INV_X1 port map( A => n94, ZN => n92);
   U102 : OAI22_X1 port map( A1 => a(2), A2 => n95, B1 => b(2), B2 => n96, ZN 
                           => n94);
   U103 : AND2_X1 port map( A1 => n95, A2 => a(2), ZN => n96);
   U104 : INV_X1 port map( A => n97, ZN => n95);
   U105 : AOI22_X1 port map( A1 => a(1), A2 => b(1), B1 => n98, B2 => n99, ZN 
                           => n97);
   U106 : INV_X1 port map( A => n100, ZN => n99);
   U107 : AOI22_X1 port map( A1 => cin, A2 => n101, B1 => b(0), B2 => a(0), ZN 
                           => n100);
   U108 : OR2_X1 port map( A1 => b(0), A2 => a(0), ZN => n101);
   U109 : OR2_X1 port map( A1 => b(1), A2 => a(1), ZN => n98);

end SYN_p4_carry_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4CarryGenerator_DATA_SIZE32_SPARSITY4_6 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  cout :
         out std_logic_vector (7 downto 0));

end P4CarryGenerator_DATA_SIZE32_SPARSITY4_6;

architecture SYN_p4_carry_generator_arch of 
   P4CarryGenerator_DATA_SIZE32_SPARSITY4_6 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal cout_7_port, cout_6_port, cout_5_port, cout_4_port, cout_3_port, 
      cout_2_port, cout_1_port, cout_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9
      , n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, 
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101 : std_logic;

begin
   cout <= ( cout_7_port, cout_6_port, cout_5_port, cout_4_port, cout_3_port, 
      cout_2_port, cout_1_port, cout_0_port );
   
   U1 : OAI22_X1 port map( A1 => n1, A2 => n2, B1 => n3, B2 => n4, ZN => 
                           cout_7_port);
   U2 : AOI22_X1 port map( A1 => b(30), A2 => n5, B1 => a(30), B2 => n6, ZN => 
                           n4);
   U3 : OR2_X1 port map( A1 => n6, A2 => a(30), ZN => n5);
   U4 : OAI21_X1 port map( B1 => n7, B2 => n8, A => n9, ZN => n6);
   U5 : OAI21_X1 port map( B1 => b(29), B2 => a(29), A => n10, ZN => n9);
   U6 : INV_X1 port map( A => n11, ZN => n10);
   U7 : AOI21_X1 port map( B1 => cout_6_port, B2 => a(28), A => n12, ZN => n11)
                           ;
   U8 : INV_X1 port map( A => n13, ZN => n12);
   U9 : OAI21_X1 port map( B1 => a(28), B2 => cout_6_port, A => b(28), ZN => 
                           n13);
   U10 : INV_X1 port map( A => b(29), ZN => n8);
   U11 : INV_X1 port map( A => a(29), ZN => n7);
   U12 : NOR2_X1 port map( A1 => b(31), A2 => a(31), ZN => n3);
   U13 : INV_X1 port map( A => b(31), ZN => n2);
   U14 : INV_X1 port map( A => a(31), ZN => n1);
   U15 : OAI21_X1 port map( B1 => n14, B2 => n15, A => n16, ZN => cout_6_port);
   U16 : OAI21_X1 port map( B1 => a(27), B2 => n17, A => b(27), ZN => n16);
   U17 : INV_X1 port map( A => n14, ZN => n17);
   U18 : INV_X1 port map( A => a(27), ZN => n15);
   U19 : AOI21_X1 port map( B1 => a(26), B2 => b(26), A => n18, ZN => n14);
   U20 : INV_X1 port map( A => n19, ZN => n18);
   U21 : OAI22_X1 port map( A1 => n20, A2 => n21, B1 => a(26), B2 => b(26), ZN 
                           => n19);
   U22 : NOR2_X1 port map( A1 => n22, A2 => n23, ZN => n21);
   U23 : AOI22_X1 port map( A1 => n22, A2 => n23, B1 => n24, B2 => n25, ZN => 
                           n20);
   U24 : OAI21_X1 port map( B1 => a(24), B2 => cout_5_port, A => b(24), ZN => 
                           n25);
   U25 : NAND2_X1 port map( A1 => a(24), A2 => cout_5_port, ZN => n24);
   U26 : INV_X1 port map( A => b(25), ZN => n23);
   U27 : INV_X1 port map( A => a(25), ZN => n22);
   U28 : OAI22_X1 port map( A1 => n26, A2 => n27, B1 => n28, B2 => n29, ZN => 
                           cout_5_port);
   U29 : AOI22_X1 port map( A1 => b(22), A2 => n30, B1 => a(22), B2 => n31, ZN 
                           => n29);
   U30 : OR2_X1 port map( A1 => n31, A2 => a(22), ZN => n30);
   U31 : OAI21_X1 port map( B1 => n32, B2 => n33, A => n34, ZN => n31);
   U32 : OAI21_X1 port map( B1 => b(21), B2 => a(21), A => n35, ZN => n34);
   U33 : OAI21_X1 port map( B1 => n36, B2 => n37, A => n38, ZN => n35);
   U34 : OAI21_X1 port map( B1 => a(20), B2 => cout_4_port, A => b(20), ZN => 
                           n38);
   U35 : INV_X1 port map( A => a(20), ZN => n37);
   U36 : INV_X1 port map( A => cout_4_port, ZN => n36);
   U37 : INV_X1 port map( A => b(21), ZN => n33);
   U38 : INV_X1 port map( A => a(21), ZN => n32);
   U39 : NOR2_X1 port map( A1 => b(23), A2 => a(23), ZN => n28);
   U40 : INV_X1 port map( A => b(23), ZN => n27);
   U41 : INV_X1 port map( A => a(23), ZN => n26);
   U42 : OAI211_X1 port map( C1 => n39, C2 => n40, A => n41, B => n42, ZN => 
                           cout_4_port);
   U43 : OAI211_X1 port map( C1 => b(19), C2 => a(19), A => cout_3_port, B => 
                           n43, ZN => n42);
   U44 : AOI221_X1 port map( B1 => n44, B2 => n45, C1 => n46, C2 => n47, A => 
                           n48, ZN => n43);
   U45 : OAI21_X1 port map( B1 => n49, B2 => a(19), A => b(19), ZN => n41);
   U46 : INV_X1 port map( A => a(19), ZN => n40);
   U47 : INV_X1 port map( A => n49, ZN => n39);
   U48 : AOI21_X1 port map( B1 => n44, B2 => n50, A => n51, ZN => n49);
   U49 : INV_X1 port map( A => n52, ZN => n51);
   U50 : OAI21_X1 port map( B1 => n50, B2 => n44, A => n45, ZN => n52);
   U51 : INV_X1 port map( A => b(18), ZN => n45);
   U52 : AOI21_X1 port map( B1 => a(17), B2 => b(17), A => n53, ZN => n50);
   U53 : NOR3_X1 port map( A1 => n46, A2 => n48, A3 => n47, ZN => n53);
   U54 : INV_X1 port map( A => b(16), ZN => n47);
   U55 : NOR2_X1 port map( A1 => b(17), A2 => a(17), ZN => n48);
   U56 : INV_X1 port map( A => a(16), ZN => n46);
   U57 : INV_X1 port map( A => a(18), ZN => n44);
   U58 : INV_X1 port map( A => n54, ZN => cout_3_port);
   U59 : OAI22_X1 port map( A1 => a(15), A2 => n55, B1 => b(15), B2 => n56, ZN 
                           => n54);
   U60 : AND2_X1 port map( A1 => n55, A2 => a(15), ZN => n56);
   U61 : INV_X1 port map( A => n57, ZN => n55);
   U62 : OAI22_X1 port map( A1 => a(14), A2 => n58, B1 => b(14), B2 => n59, ZN 
                           => n57);
   U63 : AND2_X1 port map( A1 => n58, A2 => a(14), ZN => n59);
   U64 : OAI21_X1 port map( B1 => n60, B2 => n61, A => n62, ZN => n58);
   U65 : OAI21_X1 port map( B1 => b(13), B2 => a(13), A => n63, ZN => n62);
   U66 : INV_X1 port map( A => n64, ZN => n63);
   U67 : AOI21_X1 port map( B1 => cout_2_port, B2 => a(12), A => n65, ZN => n64
                           );
   U68 : INV_X1 port map( A => n66, ZN => n65);
   U69 : OAI21_X1 port map( B1 => a(12), B2 => cout_2_port, A => b(12), ZN => 
                           n66);
   U70 : INV_X1 port map( A => b(13), ZN => n61);
   U71 : INV_X1 port map( A => a(13), ZN => n60);
   U72 : OAI21_X1 port map( B1 => n67, B2 => n68, A => n69, ZN => cout_2_port);
   U73 : OAI21_X1 port map( B1 => a(11), B2 => n70, A => b(11), ZN => n69);
   U74 : INV_X1 port map( A => n67, ZN => n70);
   U75 : INV_X1 port map( A => a(11), ZN => n68);
   U76 : AOI21_X1 port map( B1 => a(10), B2 => b(10), A => n71, ZN => n67);
   U77 : INV_X1 port map( A => n72, ZN => n71);
   U78 : OAI22_X1 port map( A1 => n73, A2 => n74, B1 => a(10), B2 => b(10), ZN 
                           => n72);
   U79 : NOR2_X1 port map( A1 => n75, A2 => n76, ZN => n74);
   U80 : AOI22_X1 port map( A1 => n75, A2 => n76, B1 => n77, B2 => n78, ZN => 
                           n73);
   U81 : OAI21_X1 port map( B1 => a(8), B2 => cout_1_port, A => b(8), ZN => n78
                           );
   U82 : NAND2_X1 port map( A1 => a(8), A2 => cout_1_port, ZN => n77);
   U83 : INV_X1 port map( A => b(9), ZN => n76);
   U84 : INV_X1 port map( A => a(9), ZN => n75);
   U85 : OAI21_X1 port map( B1 => n79, B2 => n80, A => n81, ZN => cout_1_port);
   U86 : OAI21_X1 port map( B1 => b(7), B2 => a(7), A => n82, ZN => n81);
   U87 : OAI21_X1 port map( B1 => n83, B2 => n84, A => n85, ZN => n82);
   U88 : OAI21_X1 port map( B1 => a(6), B2 => n86, A => b(6), ZN => n85);
   U89 : INV_X1 port map( A => n83, ZN => n86);
   U90 : INV_X1 port map( A => a(6), ZN => n84);
   U91 : AOI22_X1 port map( A1 => a(5), A2 => b(5), B1 => n87, B2 => n88, ZN =>
                           n83);
   U92 : INV_X1 port map( A => n89, ZN => n88);
   U93 : AOI22_X1 port map( A1 => b(4), A2 => n90, B1 => a(4), B2 => 
                           cout_0_port, ZN => n89);
   U94 : OR2_X1 port map( A1 => a(4), A2 => cout_0_port, ZN => n90);
   U95 : OR2_X1 port map( A1 => b(5), A2 => a(5), ZN => n87);
   U96 : INV_X1 port map( A => b(7), ZN => n80);
   U97 : INV_X1 port map( A => a(7), ZN => n79);
   U98 : INV_X1 port map( A => n91, ZN => cout_0_port);
   U99 : OAI22_X1 port map( A1 => a(3), A2 => n92, B1 => b(3), B2 => n93, ZN =>
                           n91);
   U100 : AND2_X1 port map( A1 => n92, A2 => a(3), ZN => n93);
   U101 : INV_X1 port map( A => n94, ZN => n92);
   U102 : OAI22_X1 port map( A1 => a(2), A2 => n95, B1 => b(2), B2 => n96, ZN 
                           => n94);
   U103 : AND2_X1 port map( A1 => n95, A2 => a(2), ZN => n96);
   U104 : INV_X1 port map( A => n97, ZN => n95);
   U105 : AOI22_X1 port map( A1 => a(1), A2 => b(1), B1 => n98, B2 => n99, ZN 
                           => n97);
   U106 : INV_X1 port map( A => n100, ZN => n99);
   U107 : AOI22_X1 port map( A1 => cin, A2 => n101, B1 => b(0), B2 => a(0), ZN 
                           => n100);
   U108 : OR2_X1 port map( A1 => b(0), A2 => a(0), ZN => n101);
   U109 : OR2_X1 port map( A1 => b(1), A2 => a(1), ZN => n98);

end SYN_p4_carry_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4CarryGenerator_DATA_SIZE32_SPARSITY4_5 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  cout :
         out std_logic_vector (7 downto 0));

end P4CarryGenerator_DATA_SIZE32_SPARSITY4_5;

architecture SYN_p4_carry_generator_arch of 
   P4CarryGenerator_DATA_SIZE32_SPARSITY4_5 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal cout_7_port, cout_6_port, cout_5_port, cout_4_port, cout_3_port, 
      cout_2_port, cout_1_port, cout_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9
      , n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, 
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101 : std_logic;

begin
   cout <= ( cout_7_port, cout_6_port, cout_5_port, cout_4_port, cout_3_port, 
      cout_2_port, cout_1_port, cout_0_port );
   
   U1 : OAI22_X1 port map( A1 => n1, A2 => n2, B1 => n3, B2 => n4, ZN => 
                           cout_7_port);
   U2 : AOI22_X1 port map( A1 => b(30), A2 => n5, B1 => a(30), B2 => n6, ZN => 
                           n4);
   U3 : OR2_X1 port map( A1 => n6, A2 => a(30), ZN => n5);
   U4 : OAI21_X1 port map( B1 => n7, B2 => n8, A => n9, ZN => n6);
   U5 : OAI21_X1 port map( B1 => b(29), B2 => a(29), A => n10, ZN => n9);
   U6 : INV_X1 port map( A => n11, ZN => n10);
   U7 : AOI21_X1 port map( B1 => cout_6_port, B2 => a(28), A => n12, ZN => n11)
                           ;
   U8 : INV_X1 port map( A => n13, ZN => n12);
   U9 : OAI21_X1 port map( B1 => a(28), B2 => cout_6_port, A => b(28), ZN => 
                           n13);
   U10 : INV_X1 port map( A => b(29), ZN => n8);
   U11 : INV_X1 port map( A => a(29), ZN => n7);
   U12 : NOR2_X1 port map( A1 => b(31), A2 => a(31), ZN => n3);
   U13 : INV_X1 port map( A => b(31), ZN => n2);
   U14 : INV_X1 port map( A => a(31), ZN => n1);
   U15 : OAI21_X1 port map( B1 => n14, B2 => n15, A => n16, ZN => cout_6_port);
   U16 : OAI21_X1 port map( B1 => a(27), B2 => n17, A => b(27), ZN => n16);
   U17 : INV_X1 port map( A => n14, ZN => n17);
   U18 : INV_X1 port map( A => a(27), ZN => n15);
   U19 : AOI21_X1 port map( B1 => a(26), B2 => b(26), A => n18, ZN => n14);
   U20 : INV_X1 port map( A => n19, ZN => n18);
   U21 : OAI22_X1 port map( A1 => n20, A2 => n21, B1 => a(26), B2 => b(26), ZN 
                           => n19);
   U22 : NOR2_X1 port map( A1 => n22, A2 => n23, ZN => n21);
   U23 : AOI22_X1 port map( A1 => n22, A2 => n23, B1 => n24, B2 => n25, ZN => 
                           n20);
   U24 : OAI21_X1 port map( B1 => a(24), B2 => cout_5_port, A => b(24), ZN => 
                           n25);
   U25 : NAND2_X1 port map( A1 => a(24), A2 => cout_5_port, ZN => n24);
   U26 : INV_X1 port map( A => b(25), ZN => n23);
   U27 : INV_X1 port map( A => a(25), ZN => n22);
   U28 : OAI22_X1 port map( A1 => n26, A2 => n27, B1 => n28, B2 => n29, ZN => 
                           cout_5_port);
   U29 : AOI22_X1 port map( A1 => b(22), A2 => n30, B1 => a(22), B2 => n31, ZN 
                           => n29);
   U30 : OR2_X1 port map( A1 => n31, A2 => a(22), ZN => n30);
   U31 : OAI21_X1 port map( B1 => n32, B2 => n33, A => n34, ZN => n31);
   U32 : OAI21_X1 port map( B1 => b(21), B2 => a(21), A => n35, ZN => n34);
   U33 : OAI21_X1 port map( B1 => n36, B2 => n37, A => n38, ZN => n35);
   U34 : OAI21_X1 port map( B1 => a(20), B2 => cout_4_port, A => b(20), ZN => 
                           n38);
   U35 : INV_X1 port map( A => a(20), ZN => n37);
   U36 : INV_X1 port map( A => cout_4_port, ZN => n36);
   U37 : INV_X1 port map( A => b(21), ZN => n33);
   U38 : INV_X1 port map( A => a(21), ZN => n32);
   U39 : NOR2_X1 port map( A1 => b(23), A2 => a(23), ZN => n28);
   U40 : INV_X1 port map( A => b(23), ZN => n27);
   U41 : INV_X1 port map( A => a(23), ZN => n26);
   U42 : OAI211_X1 port map( C1 => n39, C2 => n40, A => n41, B => n42, ZN => 
                           cout_4_port);
   U43 : OAI211_X1 port map( C1 => b(19), C2 => a(19), A => cout_3_port, B => 
                           n43, ZN => n42);
   U44 : AOI221_X1 port map( B1 => n44, B2 => n45, C1 => n46, C2 => n47, A => 
                           n48, ZN => n43);
   U45 : OAI21_X1 port map( B1 => n49, B2 => a(19), A => b(19), ZN => n41);
   U46 : INV_X1 port map( A => a(19), ZN => n40);
   U47 : INV_X1 port map( A => n49, ZN => n39);
   U48 : AOI21_X1 port map( B1 => n44, B2 => n50, A => n51, ZN => n49);
   U49 : INV_X1 port map( A => n52, ZN => n51);
   U50 : OAI21_X1 port map( B1 => n50, B2 => n44, A => n45, ZN => n52);
   U51 : INV_X1 port map( A => b(18), ZN => n45);
   U52 : AOI21_X1 port map( B1 => a(17), B2 => b(17), A => n53, ZN => n50);
   U53 : NOR3_X1 port map( A1 => n46, A2 => n48, A3 => n47, ZN => n53);
   U54 : INV_X1 port map( A => b(16), ZN => n47);
   U55 : NOR2_X1 port map( A1 => b(17), A2 => a(17), ZN => n48);
   U56 : INV_X1 port map( A => a(16), ZN => n46);
   U57 : INV_X1 port map( A => a(18), ZN => n44);
   U58 : INV_X1 port map( A => n54, ZN => cout_3_port);
   U59 : OAI22_X1 port map( A1 => a(15), A2 => n55, B1 => b(15), B2 => n56, ZN 
                           => n54);
   U60 : AND2_X1 port map( A1 => n55, A2 => a(15), ZN => n56);
   U61 : INV_X1 port map( A => n57, ZN => n55);
   U62 : OAI22_X1 port map( A1 => a(14), A2 => n58, B1 => b(14), B2 => n59, ZN 
                           => n57);
   U63 : AND2_X1 port map( A1 => n58, A2 => a(14), ZN => n59);
   U64 : OAI21_X1 port map( B1 => n60, B2 => n61, A => n62, ZN => n58);
   U65 : OAI21_X1 port map( B1 => b(13), B2 => a(13), A => n63, ZN => n62);
   U66 : INV_X1 port map( A => n64, ZN => n63);
   U67 : AOI21_X1 port map( B1 => cout_2_port, B2 => a(12), A => n65, ZN => n64
                           );
   U68 : INV_X1 port map( A => n66, ZN => n65);
   U69 : OAI21_X1 port map( B1 => a(12), B2 => cout_2_port, A => b(12), ZN => 
                           n66);
   U70 : INV_X1 port map( A => b(13), ZN => n61);
   U71 : INV_X1 port map( A => a(13), ZN => n60);
   U72 : OAI21_X1 port map( B1 => n67, B2 => n68, A => n69, ZN => cout_2_port);
   U73 : OAI21_X1 port map( B1 => a(11), B2 => n70, A => b(11), ZN => n69);
   U74 : INV_X1 port map( A => n67, ZN => n70);
   U75 : INV_X1 port map( A => a(11), ZN => n68);
   U76 : AOI21_X1 port map( B1 => a(10), B2 => b(10), A => n71, ZN => n67);
   U77 : INV_X1 port map( A => n72, ZN => n71);
   U78 : OAI22_X1 port map( A1 => n73, A2 => n74, B1 => a(10), B2 => b(10), ZN 
                           => n72);
   U79 : NOR2_X1 port map( A1 => n75, A2 => n76, ZN => n74);
   U80 : AOI22_X1 port map( A1 => n75, A2 => n76, B1 => n77, B2 => n78, ZN => 
                           n73);
   U81 : OAI21_X1 port map( B1 => a(8), B2 => cout_1_port, A => b(8), ZN => n78
                           );
   U82 : NAND2_X1 port map( A1 => a(8), A2 => cout_1_port, ZN => n77);
   U83 : INV_X1 port map( A => b(9), ZN => n76);
   U84 : INV_X1 port map( A => a(9), ZN => n75);
   U85 : OAI21_X1 port map( B1 => n79, B2 => n80, A => n81, ZN => cout_1_port);
   U86 : OAI21_X1 port map( B1 => b(7), B2 => a(7), A => n82, ZN => n81);
   U87 : OAI21_X1 port map( B1 => n83, B2 => n84, A => n85, ZN => n82);
   U88 : OAI21_X1 port map( B1 => a(6), B2 => n86, A => b(6), ZN => n85);
   U89 : INV_X1 port map( A => n83, ZN => n86);
   U90 : INV_X1 port map( A => a(6), ZN => n84);
   U91 : AOI22_X1 port map( A1 => a(5), A2 => b(5), B1 => n87, B2 => n88, ZN =>
                           n83);
   U92 : INV_X1 port map( A => n89, ZN => n88);
   U93 : AOI22_X1 port map( A1 => b(4), A2 => n90, B1 => a(4), B2 => 
                           cout_0_port, ZN => n89);
   U94 : OR2_X1 port map( A1 => a(4), A2 => cout_0_port, ZN => n90);
   U95 : OR2_X1 port map( A1 => b(5), A2 => a(5), ZN => n87);
   U96 : INV_X1 port map( A => b(7), ZN => n80);
   U97 : INV_X1 port map( A => a(7), ZN => n79);
   U98 : INV_X1 port map( A => n91, ZN => cout_0_port);
   U99 : OAI22_X1 port map( A1 => a(3), A2 => n92, B1 => b(3), B2 => n93, ZN =>
                           n91);
   U100 : AND2_X1 port map( A1 => n92, A2 => a(3), ZN => n93);
   U101 : INV_X1 port map( A => n94, ZN => n92);
   U102 : OAI22_X1 port map( A1 => a(2), A2 => n95, B1 => b(2), B2 => n96, ZN 
                           => n94);
   U103 : AND2_X1 port map( A1 => n95, A2 => a(2), ZN => n96);
   U104 : INV_X1 port map( A => n97, ZN => n95);
   U105 : AOI22_X1 port map( A1 => a(1), A2 => b(1), B1 => n98, B2 => n99, ZN 
                           => n97);
   U106 : INV_X1 port map( A => n100, ZN => n99);
   U107 : AOI22_X1 port map( A1 => cin, A2 => n101, B1 => b(0), B2 => a(0), ZN 
                           => n100);
   U108 : OR2_X1 port map( A1 => b(0), A2 => a(0), ZN => n101);
   U109 : OR2_X1 port map( A1 => b(1), A2 => a(1), ZN => n98);

end SYN_p4_carry_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4CarryGenerator_DATA_SIZE32_SPARSITY4_4 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  cout :
         out std_logic_vector (7 downto 0));

end P4CarryGenerator_DATA_SIZE32_SPARSITY4_4;

architecture SYN_p4_carry_generator_arch of 
   P4CarryGenerator_DATA_SIZE32_SPARSITY4_4 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal cout_7_port, cout_6_port, cout_5_port, cout_4_port, cout_3_port, 
      cout_2_port, cout_1_port, cout_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9
      , n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, 
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101 : std_logic;

begin
   cout <= ( cout_7_port, cout_6_port, cout_5_port, cout_4_port, cout_3_port, 
      cout_2_port, cout_1_port, cout_0_port );
   
   U1 : OAI22_X1 port map( A1 => n1, A2 => n2, B1 => n3, B2 => n4, ZN => 
                           cout_7_port);
   U2 : AOI22_X1 port map( A1 => b(30), A2 => n5, B1 => a(30), B2 => n6, ZN => 
                           n4);
   U3 : OR2_X1 port map( A1 => n6, A2 => a(30), ZN => n5);
   U4 : OAI21_X1 port map( B1 => n7, B2 => n8, A => n9, ZN => n6);
   U5 : OAI21_X1 port map( B1 => b(29), B2 => a(29), A => n10, ZN => n9);
   U6 : INV_X1 port map( A => n11, ZN => n10);
   U7 : AOI21_X1 port map( B1 => cout_6_port, B2 => a(28), A => n12, ZN => n11)
                           ;
   U8 : INV_X1 port map( A => n13, ZN => n12);
   U9 : OAI21_X1 port map( B1 => a(28), B2 => cout_6_port, A => b(28), ZN => 
                           n13);
   U10 : INV_X1 port map( A => b(29), ZN => n8);
   U11 : INV_X1 port map( A => a(29), ZN => n7);
   U12 : NOR2_X1 port map( A1 => b(31), A2 => a(31), ZN => n3);
   U13 : INV_X1 port map( A => b(31), ZN => n2);
   U14 : INV_X1 port map( A => a(31), ZN => n1);
   U15 : OAI21_X1 port map( B1 => n14, B2 => n15, A => n16, ZN => cout_6_port);
   U16 : OAI21_X1 port map( B1 => a(27), B2 => n17, A => b(27), ZN => n16);
   U17 : INV_X1 port map( A => n14, ZN => n17);
   U18 : INV_X1 port map( A => a(27), ZN => n15);
   U19 : AOI21_X1 port map( B1 => a(26), B2 => b(26), A => n18, ZN => n14);
   U20 : INV_X1 port map( A => n19, ZN => n18);
   U21 : OAI22_X1 port map( A1 => n20, A2 => n21, B1 => a(26), B2 => b(26), ZN 
                           => n19);
   U22 : NOR2_X1 port map( A1 => n22, A2 => n23, ZN => n21);
   U23 : AOI22_X1 port map( A1 => n22, A2 => n23, B1 => n24, B2 => n25, ZN => 
                           n20);
   U24 : OAI21_X1 port map( B1 => a(24), B2 => cout_5_port, A => b(24), ZN => 
                           n25);
   U25 : NAND2_X1 port map( A1 => a(24), A2 => cout_5_port, ZN => n24);
   U26 : INV_X1 port map( A => b(25), ZN => n23);
   U27 : INV_X1 port map( A => a(25), ZN => n22);
   U28 : OAI22_X1 port map( A1 => n26, A2 => n27, B1 => n28, B2 => n29, ZN => 
                           cout_5_port);
   U29 : AOI22_X1 port map( A1 => b(22), A2 => n30, B1 => a(22), B2 => n31, ZN 
                           => n29);
   U30 : OR2_X1 port map( A1 => n31, A2 => a(22), ZN => n30);
   U31 : OAI21_X1 port map( B1 => n32, B2 => n33, A => n34, ZN => n31);
   U32 : OAI21_X1 port map( B1 => b(21), B2 => a(21), A => n35, ZN => n34);
   U33 : OAI21_X1 port map( B1 => n36, B2 => n37, A => n38, ZN => n35);
   U34 : OAI21_X1 port map( B1 => a(20), B2 => cout_4_port, A => b(20), ZN => 
                           n38);
   U35 : INV_X1 port map( A => a(20), ZN => n37);
   U36 : INV_X1 port map( A => cout_4_port, ZN => n36);
   U37 : INV_X1 port map( A => b(21), ZN => n33);
   U38 : INV_X1 port map( A => a(21), ZN => n32);
   U39 : NOR2_X1 port map( A1 => b(23), A2 => a(23), ZN => n28);
   U40 : INV_X1 port map( A => b(23), ZN => n27);
   U41 : INV_X1 port map( A => a(23), ZN => n26);
   U42 : OAI211_X1 port map( C1 => n39, C2 => n40, A => n41, B => n42, ZN => 
                           cout_4_port);
   U43 : OAI211_X1 port map( C1 => b(19), C2 => a(19), A => cout_3_port, B => 
                           n43, ZN => n42);
   U44 : AOI221_X1 port map( B1 => n44, B2 => n45, C1 => n46, C2 => n47, A => 
                           n48, ZN => n43);
   U45 : OAI21_X1 port map( B1 => n49, B2 => a(19), A => b(19), ZN => n41);
   U46 : INV_X1 port map( A => a(19), ZN => n40);
   U47 : INV_X1 port map( A => n49, ZN => n39);
   U48 : AOI21_X1 port map( B1 => n44, B2 => n50, A => n51, ZN => n49);
   U49 : INV_X1 port map( A => n52, ZN => n51);
   U50 : OAI21_X1 port map( B1 => n50, B2 => n44, A => n45, ZN => n52);
   U51 : INV_X1 port map( A => b(18), ZN => n45);
   U52 : AOI21_X1 port map( B1 => a(17), B2 => b(17), A => n53, ZN => n50);
   U53 : NOR3_X1 port map( A1 => n46, A2 => n48, A3 => n47, ZN => n53);
   U54 : INV_X1 port map( A => b(16), ZN => n47);
   U55 : NOR2_X1 port map( A1 => b(17), A2 => a(17), ZN => n48);
   U56 : INV_X1 port map( A => a(16), ZN => n46);
   U57 : INV_X1 port map( A => a(18), ZN => n44);
   U58 : INV_X1 port map( A => n54, ZN => cout_3_port);
   U59 : OAI22_X1 port map( A1 => a(15), A2 => n55, B1 => b(15), B2 => n56, ZN 
                           => n54);
   U60 : AND2_X1 port map( A1 => n55, A2 => a(15), ZN => n56);
   U61 : INV_X1 port map( A => n57, ZN => n55);
   U62 : OAI22_X1 port map( A1 => a(14), A2 => n58, B1 => b(14), B2 => n59, ZN 
                           => n57);
   U63 : AND2_X1 port map( A1 => n58, A2 => a(14), ZN => n59);
   U64 : OAI21_X1 port map( B1 => n60, B2 => n61, A => n62, ZN => n58);
   U65 : OAI21_X1 port map( B1 => b(13), B2 => a(13), A => n63, ZN => n62);
   U66 : INV_X1 port map( A => n64, ZN => n63);
   U67 : AOI21_X1 port map( B1 => cout_2_port, B2 => a(12), A => n65, ZN => n64
                           );
   U68 : INV_X1 port map( A => n66, ZN => n65);
   U69 : OAI21_X1 port map( B1 => a(12), B2 => cout_2_port, A => b(12), ZN => 
                           n66);
   U70 : INV_X1 port map( A => b(13), ZN => n61);
   U71 : INV_X1 port map( A => a(13), ZN => n60);
   U72 : OAI21_X1 port map( B1 => n67, B2 => n68, A => n69, ZN => cout_2_port);
   U73 : OAI21_X1 port map( B1 => a(11), B2 => n70, A => b(11), ZN => n69);
   U74 : INV_X1 port map( A => n67, ZN => n70);
   U75 : INV_X1 port map( A => a(11), ZN => n68);
   U76 : AOI21_X1 port map( B1 => a(10), B2 => b(10), A => n71, ZN => n67);
   U77 : INV_X1 port map( A => n72, ZN => n71);
   U78 : OAI22_X1 port map( A1 => n73, A2 => n74, B1 => a(10), B2 => b(10), ZN 
                           => n72);
   U79 : NOR2_X1 port map( A1 => n75, A2 => n76, ZN => n74);
   U80 : AOI22_X1 port map( A1 => n75, A2 => n76, B1 => n77, B2 => n78, ZN => 
                           n73);
   U81 : OAI21_X1 port map( B1 => a(8), B2 => cout_1_port, A => b(8), ZN => n78
                           );
   U82 : NAND2_X1 port map( A1 => a(8), A2 => cout_1_port, ZN => n77);
   U83 : INV_X1 port map( A => b(9), ZN => n76);
   U84 : INV_X1 port map( A => a(9), ZN => n75);
   U85 : OAI21_X1 port map( B1 => n79, B2 => n80, A => n81, ZN => cout_1_port);
   U86 : OAI21_X1 port map( B1 => b(7), B2 => a(7), A => n82, ZN => n81);
   U87 : OAI21_X1 port map( B1 => n83, B2 => n84, A => n85, ZN => n82);
   U88 : OAI21_X1 port map( B1 => a(6), B2 => n86, A => b(6), ZN => n85);
   U89 : INV_X1 port map( A => n83, ZN => n86);
   U90 : INV_X1 port map( A => a(6), ZN => n84);
   U91 : AOI22_X1 port map( A1 => a(5), A2 => b(5), B1 => n87, B2 => n88, ZN =>
                           n83);
   U92 : INV_X1 port map( A => n89, ZN => n88);
   U93 : AOI22_X1 port map( A1 => b(4), A2 => n90, B1 => a(4), B2 => 
                           cout_0_port, ZN => n89);
   U94 : OR2_X1 port map( A1 => a(4), A2 => cout_0_port, ZN => n90);
   U95 : OR2_X1 port map( A1 => b(5), A2 => a(5), ZN => n87);
   U96 : INV_X1 port map( A => b(7), ZN => n80);
   U97 : INV_X1 port map( A => a(7), ZN => n79);
   U98 : INV_X1 port map( A => n91, ZN => cout_0_port);
   U99 : OAI22_X1 port map( A1 => a(3), A2 => n92, B1 => b(3), B2 => n93, ZN =>
                           n91);
   U100 : AND2_X1 port map( A1 => n92, A2 => a(3), ZN => n93);
   U101 : INV_X1 port map( A => n94, ZN => n92);
   U102 : OAI22_X1 port map( A1 => a(2), A2 => n95, B1 => b(2), B2 => n96, ZN 
                           => n94);
   U103 : AND2_X1 port map( A1 => n95, A2 => a(2), ZN => n96);
   U104 : INV_X1 port map( A => n97, ZN => n95);
   U105 : AOI22_X1 port map( A1 => a(1), A2 => b(1), B1 => n98, B2 => n99, ZN 
                           => n97);
   U106 : INV_X1 port map( A => n100, ZN => n99);
   U107 : AOI22_X1 port map( A1 => cin, A2 => n101, B1 => b(0), B2 => a(0), ZN 
                           => n100);
   U108 : OR2_X1 port map( A1 => b(0), A2 => a(0), ZN => n101);
   U109 : OR2_X1 port map( A1 => b(1), A2 => a(1), ZN => n98);

end SYN_p4_carry_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4CarryGenerator_DATA_SIZE32_SPARSITY4_3 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  cout :
         out std_logic_vector (7 downto 0));

end P4CarryGenerator_DATA_SIZE32_SPARSITY4_3;

architecture SYN_p4_carry_generator_arch of 
   P4CarryGenerator_DATA_SIZE32_SPARSITY4_3 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal cout_7_port, cout_6_port, cout_5_port, cout_4_port, cout_3_port, 
      cout_2_port, cout_1_port, cout_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9
      , n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, 
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101 : std_logic;

begin
   cout <= ( cout_7_port, cout_6_port, cout_5_port, cout_4_port, cout_3_port, 
      cout_2_port, cout_1_port, cout_0_port );
   
   U1 : OAI22_X1 port map( A1 => n1, A2 => n2, B1 => n3, B2 => n4, ZN => 
                           cout_7_port);
   U2 : AOI22_X1 port map( A1 => b(30), A2 => n5, B1 => a(30), B2 => n6, ZN => 
                           n4);
   U3 : OR2_X1 port map( A1 => n6, A2 => a(30), ZN => n5);
   U4 : OAI21_X1 port map( B1 => n7, B2 => n8, A => n9, ZN => n6);
   U5 : OAI21_X1 port map( B1 => b(29), B2 => a(29), A => n10, ZN => n9);
   U6 : INV_X1 port map( A => n11, ZN => n10);
   U7 : AOI21_X1 port map( B1 => cout_6_port, B2 => a(28), A => n12, ZN => n11)
                           ;
   U8 : INV_X1 port map( A => n13, ZN => n12);
   U9 : OAI21_X1 port map( B1 => a(28), B2 => cout_6_port, A => b(28), ZN => 
                           n13);
   U10 : INV_X1 port map( A => b(29), ZN => n8);
   U11 : INV_X1 port map( A => a(29), ZN => n7);
   U12 : NOR2_X1 port map( A1 => b(31), A2 => a(31), ZN => n3);
   U13 : INV_X1 port map( A => b(31), ZN => n2);
   U14 : INV_X1 port map( A => a(31), ZN => n1);
   U15 : OAI21_X1 port map( B1 => n14, B2 => n15, A => n16, ZN => cout_6_port);
   U16 : OAI21_X1 port map( B1 => a(27), B2 => n17, A => b(27), ZN => n16);
   U17 : INV_X1 port map( A => n14, ZN => n17);
   U18 : INV_X1 port map( A => a(27), ZN => n15);
   U19 : AOI21_X1 port map( B1 => a(26), B2 => b(26), A => n18, ZN => n14);
   U20 : INV_X1 port map( A => n19, ZN => n18);
   U21 : OAI22_X1 port map( A1 => n20, A2 => n21, B1 => a(26), B2 => b(26), ZN 
                           => n19);
   U22 : NOR2_X1 port map( A1 => n22, A2 => n23, ZN => n21);
   U23 : AOI22_X1 port map( A1 => n22, A2 => n23, B1 => n24, B2 => n25, ZN => 
                           n20);
   U24 : OAI21_X1 port map( B1 => a(24), B2 => cout_5_port, A => b(24), ZN => 
                           n25);
   U25 : NAND2_X1 port map( A1 => a(24), A2 => cout_5_port, ZN => n24);
   U26 : INV_X1 port map( A => b(25), ZN => n23);
   U27 : INV_X1 port map( A => a(25), ZN => n22);
   U28 : OAI22_X1 port map( A1 => n26, A2 => n27, B1 => n28, B2 => n29, ZN => 
                           cout_5_port);
   U29 : AOI22_X1 port map( A1 => b(22), A2 => n30, B1 => a(22), B2 => n31, ZN 
                           => n29);
   U30 : OR2_X1 port map( A1 => n31, A2 => a(22), ZN => n30);
   U31 : OAI21_X1 port map( B1 => n32, B2 => n33, A => n34, ZN => n31);
   U32 : OAI21_X1 port map( B1 => b(21), B2 => a(21), A => n35, ZN => n34);
   U33 : OAI21_X1 port map( B1 => n36, B2 => n37, A => n38, ZN => n35);
   U34 : OAI21_X1 port map( B1 => a(20), B2 => cout_4_port, A => b(20), ZN => 
                           n38);
   U35 : INV_X1 port map( A => a(20), ZN => n37);
   U36 : INV_X1 port map( A => cout_4_port, ZN => n36);
   U37 : INV_X1 port map( A => b(21), ZN => n33);
   U38 : INV_X1 port map( A => a(21), ZN => n32);
   U39 : NOR2_X1 port map( A1 => b(23), A2 => a(23), ZN => n28);
   U40 : INV_X1 port map( A => b(23), ZN => n27);
   U41 : INV_X1 port map( A => a(23), ZN => n26);
   U42 : OAI211_X1 port map( C1 => n39, C2 => n40, A => n41, B => n42, ZN => 
                           cout_4_port);
   U43 : OAI211_X1 port map( C1 => b(19), C2 => a(19), A => cout_3_port, B => 
                           n43, ZN => n42);
   U44 : AOI221_X1 port map( B1 => n44, B2 => n45, C1 => n46, C2 => n47, A => 
                           n48, ZN => n43);
   U45 : OAI21_X1 port map( B1 => n49, B2 => a(19), A => b(19), ZN => n41);
   U46 : INV_X1 port map( A => a(19), ZN => n40);
   U47 : INV_X1 port map( A => n49, ZN => n39);
   U48 : AOI21_X1 port map( B1 => n44, B2 => n50, A => n51, ZN => n49);
   U49 : INV_X1 port map( A => n52, ZN => n51);
   U50 : OAI21_X1 port map( B1 => n50, B2 => n44, A => n45, ZN => n52);
   U51 : INV_X1 port map( A => b(18), ZN => n45);
   U52 : AOI21_X1 port map( B1 => a(17), B2 => b(17), A => n53, ZN => n50);
   U53 : NOR3_X1 port map( A1 => n46, A2 => n48, A3 => n47, ZN => n53);
   U54 : INV_X1 port map( A => b(16), ZN => n47);
   U55 : NOR2_X1 port map( A1 => b(17), A2 => a(17), ZN => n48);
   U56 : INV_X1 port map( A => a(16), ZN => n46);
   U57 : INV_X1 port map( A => a(18), ZN => n44);
   U58 : INV_X1 port map( A => n54, ZN => cout_3_port);
   U59 : OAI22_X1 port map( A1 => a(15), A2 => n55, B1 => b(15), B2 => n56, ZN 
                           => n54);
   U60 : AND2_X1 port map( A1 => n55, A2 => a(15), ZN => n56);
   U61 : INV_X1 port map( A => n57, ZN => n55);
   U62 : OAI22_X1 port map( A1 => a(14), A2 => n58, B1 => b(14), B2 => n59, ZN 
                           => n57);
   U63 : AND2_X1 port map( A1 => n58, A2 => a(14), ZN => n59);
   U64 : OAI21_X1 port map( B1 => n60, B2 => n61, A => n62, ZN => n58);
   U65 : OAI21_X1 port map( B1 => b(13), B2 => a(13), A => n63, ZN => n62);
   U66 : INV_X1 port map( A => n64, ZN => n63);
   U67 : AOI21_X1 port map( B1 => cout_2_port, B2 => a(12), A => n65, ZN => n64
                           );
   U68 : INV_X1 port map( A => n66, ZN => n65);
   U69 : OAI21_X1 port map( B1 => a(12), B2 => cout_2_port, A => b(12), ZN => 
                           n66);
   U70 : INV_X1 port map( A => b(13), ZN => n61);
   U71 : INV_X1 port map( A => a(13), ZN => n60);
   U72 : OAI21_X1 port map( B1 => n67, B2 => n68, A => n69, ZN => cout_2_port);
   U73 : OAI21_X1 port map( B1 => a(11), B2 => n70, A => b(11), ZN => n69);
   U74 : INV_X1 port map( A => n67, ZN => n70);
   U75 : INV_X1 port map( A => a(11), ZN => n68);
   U76 : AOI21_X1 port map( B1 => a(10), B2 => b(10), A => n71, ZN => n67);
   U77 : INV_X1 port map( A => n72, ZN => n71);
   U78 : OAI22_X1 port map( A1 => n73, A2 => n74, B1 => a(10), B2 => b(10), ZN 
                           => n72);
   U79 : NOR2_X1 port map( A1 => n75, A2 => n76, ZN => n74);
   U80 : AOI22_X1 port map( A1 => n75, A2 => n76, B1 => n77, B2 => n78, ZN => 
                           n73);
   U81 : OAI21_X1 port map( B1 => a(8), B2 => cout_1_port, A => b(8), ZN => n78
                           );
   U82 : NAND2_X1 port map( A1 => a(8), A2 => cout_1_port, ZN => n77);
   U83 : INV_X1 port map( A => b(9), ZN => n76);
   U84 : INV_X1 port map( A => a(9), ZN => n75);
   U85 : OAI21_X1 port map( B1 => n79, B2 => n80, A => n81, ZN => cout_1_port);
   U86 : OAI21_X1 port map( B1 => b(7), B2 => a(7), A => n82, ZN => n81);
   U87 : OAI21_X1 port map( B1 => n83, B2 => n84, A => n85, ZN => n82);
   U88 : OAI21_X1 port map( B1 => a(6), B2 => n86, A => b(6), ZN => n85);
   U89 : INV_X1 port map( A => n83, ZN => n86);
   U90 : INV_X1 port map( A => a(6), ZN => n84);
   U91 : AOI22_X1 port map( A1 => a(5), A2 => b(5), B1 => n87, B2 => n88, ZN =>
                           n83);
   U92 : INV_X1 port map( A => n89, ZN => n88);
   U93 : AOI22_X1 port map( A1 => b(4), A2 => n90, B1 => a(4), B2 => 
                           cout_0_port, ZN => n89);
   U94 : OR2_X1 port map( A1 => a(4), A2 => cout_0_port, ZN => n90);
   U95 : OR2_X1 port map( A1 => b(5), A2 => a(5), ZN => n87);
   U96 : INV_X1 port map( A => b(7), ZN => n80);
   U97 : INV_X1 port map( A => a(7), ZN => n79);
   U98 : INV_X1 port map( A => n91, ZN => cout_0_port);
   U99 : OAI22_X1 port map( A1 => a(3), A2 => n92, B1 => b(3), B2 => n93, ZN =>
                           n91);
   U100 : AND2_X1 port map( A1 => n92, A2 => a(3), ZN => n93);
   U101 : INV_X1 port map( A => n94, ZN => n92);
   U102 : OAI22_X1 port map( A1 => a(2), A2 => n95, B1 => b(2), B2 => n96, ZN 
                           => n94);
   U103 : AND2_X1 port map( A1 => n95, A2 => a(2), ZN => n96);
   U104 : INV_X1 port map( A => n97, ZN => n95);
   U105 : AOI22_X1 port map( A1 => a(1), A2 => b(1), B1 => n98, B2 => n99, ZN 
                           => n97);
   U106 : INV_X1 port map( A => n100, ZN => n99);
   U107 : AOI22_X1 port map( A1 => cin, A2 => n101, B1 => b(0), B2 => a(0), ZN 
                           => n100);
   U108 : OR2_X1 port map( A1 => b(0), A2 => a(0), ZN => n101);
   U109 : OR2_X1 port map( A1 => b(1), A2 => a(1), ZN => n98);

end SYN_p4_carry_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4CarryGenerator_DATA_SIZE32_SPARSITY4_2 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  cout :
         out std_logic_vector (7 downto 0));

end P4CarryGenerator_DATA_SIZE32_SPARSITY4_2;

architecture SYN_p4_carry_generator_arch of 
   P4CarryGenerator_DATA_SIZE32_SPARSITY4_2 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal cout_7_port, cout_6_port, cout_5_port, cout_4_port, cout_3_port, 
      cout_2_port, cout_1_port, cout_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9
      , n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, 
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101 : std_logic;

begin
   cout <= ( cout_7_port, cout_6_port, cout_5_port, cout_4_port, cout_3_port, 
      cout_2_port, cout_1_port, cout_0_port );
   
   U1 : OAI22_X1 port map( A1 => n1, A2 => n2, B1 => n3, B2 => n4, ZN => 
                           cout_7_port);
   U2 : AOI22_X1 port map( A1 => b(30), A2 => n5, B1 => a(30), B2 => n6, ZN => 
                           n4);
   U3 : OR2_X1 port map( A1 => n6, A2 => a(30), ZN => n5);
   U4 : OAI21_X1 port map( B1 => n7, B2 => n8, A => n9, ZN => n6);
   U5 : OAI21_X1 port map( B1 => b(29), B2 => a(29), A => n10, ZN => n9);
   U6 : INV_X1 port map( A => n11, ZN => n10);
   U7 : AOI21_X1 port map( B1 => cout_6_port, B2 => a(28), A => n12, ZN => n11)
                           ;
   U8 : INV_X1 port map( A => n13, ZN => n12);
   U9 : OAI21_X1 port map( B1 => a(28), B2 => cout_6_port, A => b(28), ZN => 
                           n13);
   U10 : INV_X1 port map( A => b(29), ZN => n8);
   U11 : INV_X1 port map( A => a(29), ZN => n7);
   U12 : NOR2_X1 port map( A1 => b(31), A2 => a(31), ZN => n3);
   U13 : INV_X1 port map( A => b(31), ZN => n2);
   U14 : INV_X1 port map( A => a(31), ZN => n1);
   U15 : OAI21_X1 port map( B1 => n14, B2 => n15, A => n16, ZN => cout_6_port);
   U16 : OAI21_X1 port map( B1 => a(27), B2 => n17, A => b(27), ZN => n16);
   U17 : INV_X1 port map( A => n14, ZN => n17);
   U18 : INV_X1 port map( A => a(27), ZN => n15);
   U19 : AOI21_X1 port map( B1 => a(26), B2 => b(26), A => n18, ZN => n14);
   U20 : INV_X1 port map( A => n19, ZN => n18);
   U21 : OAI22_X1 port map( A1 => n20, A2 => n21, B1 => a(26), B2 => b(26), ZN 
                           => n19);
   U22 : NOR2_X1 port map( A1 => n22, A2 => n23, ZN => n21);
   U23 : AOI22_X1 port map( A1 => n22, A2 => n23, B1 => n24, B2 => n25, ZN => 
                           n20);
   U24 : OAI21_X1 port map( B1 => a(24), B2 => cout_5_port, A => b(24), ZN => 
                           n25);
   U25 : NAND2_X1 port map( A1 => a(24), A2 => cout_5_port, ZN => n24);
   U26 : INV_X1 port map( A => b(25), ZN => n23);
   U27 : INV_X1 port map( A => a(25), ZN => n22);
   U28 : OAI22_X1 port map( A1 => n26, A2 => n27, B1 => n28, B2 => n29, ZN => 
                           cout_5_port);
   U29 : AOI22_X1 port map( A1 => b(22), A2 => n30, B1 => a(22), B2 => n31, ZN 
                           => n29);
   U30 : OR2_X1 port map( A1 => n31, A2 => a(22), ZN => n30);
   U31 : OAI21_X1 port map( B1 => n32, B2 => n33, A => n34, ZN => n31);
   U32 : OAI21_X1 port map( B1 => b(21), B2 => a(21), A => n35, ZN => n34);
   U33 : OAI21_X1 port map( B1 => n36, B2 => n37, A => n38, ZN => n35);
   U34 : OAI21_X1 port map( B1 => a(20), B2 => cout_4_port, A => b(20), ZN => 
                           n38);
   U35 : INV_X1 port map( A => a(20), ZN => n37);
   U36 : INV_X1 port map( A => cout_4_port, ZN => n36);
   U37 : INV_X1 port map( A => b(21), ZN => n33);
   U38 : INV_X1 port map( A => a(21), ZN => n32);
   U39 : NOR2_X1 port map( A1 => b(23), A2 => a(23), ZN => n28);
   U40 : INV_X1 port map( A => b(23), ZN => n27);
   U41 : INV_X1 port map( A => a(23), ZN => n26);
   U42 : OAI211_X1 port map( C1 => n39, C2 => n40, A => n41, B => n42, ZN => 
                           cout_4_port);
   U43 : OAI211_X1 port map( C1 => b(19), C2 => a(19), A => cout_3_port, B => 
                           n43, ZN => n42);
   U44 : AOI221_X1 port map( B1 => n44, B2 => n45, C1 => n46, C2 => n47, A => 
                           n48, ZN => n43);
   U45 : OAI21_X1 port map( B1 => n49, B2 => a(19), A => b(19), ZN => n41);
   U46 : INV_X1 port map( A => a(19), ZN => n40);
   U47 : INV_X1 port map( A => n49, ZN => n39);
   U48 : AOI21_X1 port map( B1 => n44, B2 => n50, A => n51, ZN => n49);
   U49 : INV_X1 port map( A => n52, ZN => n51);
   U50 : OAI21_X1 port map( B1 => n50, B2 => n44, A => n45, ZN => n52);
   U51 : INV_X1 port map( A => b(18), ZN => n45);
   U52 : AOI21_X1 port map( B1 => a(17), B2 => b(17), A => n53, ZN => n50);
   U53 : NOR3_X1 port map( A1 => n46, A2 => n48, A3 => n47, ZN => n53);
   U54 : INV_X1 port map( A => b(16), ZN => n47);
   U55 : NOR2_X1 port map( A1 => b(17), A2 => a(17), ZN => n48);
   U56 : INV_X1 port map( A => a(16), ZN => n46);
   U57 : INV_X1 port map( A => a(18), ZN => n44);
   U58 : INV_X1 port map( A => n54, ZN => cout_3_port);
   U59 : OAI22_X1 port map( A1 => a(15), A2 => n55, B1 => b(15), B2 => n56, ZN 
                           => n54);
   U60 : AND2_X1 port map( A1 => n55, A2 => a(15), ZN => n56);
   U61 : INV_X1 port map( A => n57, ZN => n55);
   U62 : OAI22_X1 port map( A1 => a(14), A2 => n58, B1 => b(14), B2 => n59, ZN 
                           => n57);
   U63 : AND2_X1 port map( A1 => n58, A2 => a(14), ZN => n59);
   U64 : OAI21_X1 port map( B1 => n60, B2 => n61, A => n62, ZN => n58);
   U65 : OAI21_X1 port map( B1 => b(13), B2 => a(13), A => n63, ZN => n62);
   U66 : INV_X1 port map( A => n64, ZN => n63);
   U67 : AOI21_X1 port map( B1 => cout_2_port, B2 => a(12), A => n65, ZN => n64
                           );
   U68 : INV_X1 port map( A => n66, ZN => n65);
   U69 : OAI21_X1 port map( B1 => a(12), B2 => cout_2_port, A => b(12), ZN => 
                           n66);
   U70 : INV_X1 port map( A => b(13), ZN => n61);
   U71 : INV_X1 port map( A => a(13), ZN => n60);
   U72 : OAI21_X1 port map( B1 => n67, B2 => n68, A => n69, ZN => cout_2_port);
   U73 : OAI21_X1 port map( B1 => a(11), B2 => n70, A => b(11), ZN => n69);
   U74 : INV_X1 port map( A => n67, ZN => n70);
   U75 : INV_X1 port map( A => a(11), ZN => n68);
   U76 : AOI21_X1 port map( B1 => a(10), B2 => b(10), A => n71, ZN => n67);
   U77 : INV_X1 port map( A => n72, ZN => n71);
   U78 : OAI22_X1 port map( A1 => n73, A2 => n74, B1 => a(10), B2 => b(10), ZN 
                           => n72);
   U79 : NOR2_X1 port map( A1 => n75, A2 => n76, ZN => n74);
   U80 : AOI22_X1 port map( A1 => n75, A2 => n76, B1 => n77, B2 => n78, ZN => 
                           n73);
   U81 : OAI21_X1 port map( B1 => a(8), B2 => cout_1_port, A => b(8), ZN => n78
                           );
   U82 : NAND2_X1 port map( A1 => a(8), A2 => cout_1_port, ZN => n77);
   U83 : INV_X1 port map( A => b(9), ZN => n76);
   U84 : INV_X1 port map( A => a(9), ZN => n75);
   U85 : OAI21_X1 port map( B1 => n79, B2 => n80, A => n81, ZN => cout_1_port);
   U86 : OAI21_X1 port map( B1 => b(7), B2 => a(7), A => n82, ZN => n81);
   U87 : OAI21_X1 port map( B1 => n83, B2 => n84, A => n85, ZN => n82);
   U88 : OAI21_X1 port map( B1 => a(6), B2 => n86, A => b(6), ZN => n85);
   U89 : INV_X1 port map( A => n83, ZN => n86);
   U90 : INV_X1 port map( A => a(6), ZN => n84);
   U91 : AOI22_X1 port map( A1 => a(5), A2 => b(5), B1 => n87, B2 => n88, ZN =>
                           n83);
   U92 : INV_X1 port map( A => n89, ZN => n88);
   U93 : AOI22_X1 port map( A1 => b(4), A2 => n90, B1 => a(4), B2 => 
                           cout_0_port, ZN => n89);
   U94 : OR2_X1 port map( A1 => a(4), A2 => cout_0_port, ZN => n90);
   U95 : OR2_X1 port map( A1 => b(5), A2 => a(5), ZN => n87);
   U96 : INV_X1 port map( A => b(7), ZN => n80);
   U97 : INV_X1 port map( A => a(7), ZN => n79);
   U98 : INV_X1 port map( A => n91, ZN => cout_0_port);
   U99 : OAI22_X1 port map( A1 => a(3), A2 => n92, B1 => b(3), B2 => n93, ZN =>
                           n91);
   U100 : AND2_X1 port map( A1 => n92, A2 => a(3), ZN => n93);
   U101 : INV_X1 port map( A => n94, ZN => n92);
   U102 : OAI22_X1 port map( A1 => a(2), A2 => n95, B1 => b(2), B2 => n96, ZN 
                           => n94);
   U103 : AND2_X1 port map( A1 => n95, A2 => a(2), ZN => n96);
   U104 : INV_X1 port map( A => n97, ZN => n95);
   U105 : AOI22_X1 port map( A1 => a(1), A2 => b(1), B1 => n98, B2 => n99, ZN 
                           => n97);
   U106 : INV_X1 port map( A => n100, ZN => n99);
   U107 : AOI22_X1 port map( A1 => cin, A2 => n101, B1 => b(0), B2 => a(0), ZN 
                           => n100);
   U108 : OR2_X1 port map( A1 => b(0), A2 => a(0), ZN => n101);
   U109 : OR2_X1 port map( A1 => b(1), A2 => a(1), ZN => n98);

end SYN_p4_carry_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4CarryGenerator_DATA_SIZE32_SPARSITY4_1 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  cout :
         out std_logic_vector (7 downto 0));

end P4CarryGenerator_DATA_SIZE32_SPARSITY4_1;

architecture SYN_p4_carry_generator_arch of 
   P4CarryGenerator_DATA_SIZE32_SPARSITY4_1 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal cout_7_port, cout_6_port, cout_5_port, cout_4_port, cout_3_port, 
      cout_2_port, cout_1_port, cout_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9
      , n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, 
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101 : std_logic;

begin
   cout <= ( cout_7_port, cout_6_port, cout_5_port, cout_4_port, cout_3_port, 
      cout_2_port, cout_1_port, cout_0_port );
   
   U1 : OAI22_X1 port map( A1 => n1, A2 => n2, B1 => n3, B2 => n4, ZN => 
                           cout_7_port);
   U2 : AOI22_X1 port map( A1 => b(30), A2 => n5, B1 => a(30), B2 => n6, ZN => 
                           n4);
   U3 : OR2_X1 port map( A1 => n6, A2 => a(30), ZN => n5);
   U4 : OAI21_X1 port map( B1 => n7, B2 => n8, A => n9, ZN => n6);
   U5 : OAI21_X1 port map( B1 => b(29), B2 => a(29), A => n10, ZN => n9);
   U6 : INV_X1 port map( A => n11, ZN => n10);
   U7 : AOI21_X1 port map( B1 => cout_6_port, B2 => a(28), A => n12, ZN => n11)
                           ;
   U8 : INV_X1 port map( A => n13, ZN => n12);
   U9 : OAI21_X1 port map( B1 => a(28), B2 => cout_6_port, A => b(28), ZN => 
                           n13);
   U10 : INV_X1 port map( A => b(29), ZN => n8);
   U11 : INV_X1 port map( A => a(29), ZN => n7);
   U12 : NOR2_X1 port map( A1 => b(31), A2 => a(31), ZN => n3);
   U13 : INV_X1 port map( A => b(31), ZN => n2);
   U14 : INV_X1 port map( A => a(31), ZN => n1);
   U15 : OAI21_X1 port map( B1 => n14, B2 => n15, A => n16, ZN => cout_6_port);
   U16 : OAI21_X1 port map( B1 => a(27), B2 => n17, A => b(27), ZN => n16);
   U17 : INV_X1 port map( A => n14, ZN => n17);
   U18 : INV_X1 port map( A => a(27), ZN => n15);
   U19 : AOI21_X1 port map( B1 => a(26), B2 => b(26), A => n18, ZN => n14);
   U20 : INV_X1 port map( A => n19, ZN => n18);
   U21 : OAI22_X1 port map( A1 => n20, A2 => n21, B1 => a(26), B2 => b(26), ZN 
                           => n19);
   U22 : NOR2_X1 port map( A1 => n22, A2 => n23, ZN => n21);
   U23 : AOI22_X1 port map( A1 => n22, A2 => n23, B1 => n24, B2 => n25, ZN => 
                           n20);
   U24 : OAI21_X1 port map( B1 => a(24), B2 => cout_5_port, A => b(24), ZN => 
                           n25);
   U25 : NAND2_X1 port map( A1 => a(24), A2 => cout_5_port, ZN => n24);
   U26 : INV_X1 port map( A => b(25), ZN => n23);
   U27 : INV_X1 port map( A => a(25), ZN => n22);
   U28 : OAI22_X1 port map( A1 => n26, A2 => n27, B1 => n28, B2 => n29, ZN => 
                           cout_5_port);
   U29 : AOI22_X1 port map( A1 => b(22), A2 => n30, B1 => a(22), B2 => n31, ZN 
                           => n29);
   U30 : OR2_X1 port map( A1 => n31, A2 => a(22), ZN => n30);
   U31 : OAI21_X1 port map( B1 => n32, B2 => n33, A => n34, ZN => n31);
   U32 : OAI21_X1 port map( B1 => b(21), B2 => a(21), A => n35, ZN => n34);
   U33 : OAI21_X1 port map( B1 => n36, B2 => n37, A => n38, ZN => n35);
   U34 : OAI21_X1 port map( B1 => a(20), B2 => cout_4_port, A => b(20), ZN => 
                           n38);
   U35 : INV_X1 port map( A => a(20), ZN => n37);
   U36 : INV_X1 port map( A => cout_4_port, ZN => n36);
   U37 : INV_X1 port map( A => b(21), ZN => n33);
   U38 : INV_X1 port map( A => a(21), ZN => n32);
   U39 : NOR2_X1 port map( A1 => b(23), A2 => a(23), ZN => n28);
   U40 : INV_X1 port map( A => b(23), ZN => n27);
   U41 : INV_X1 port map( A => a(23), ZN => n26);
   U42 : OAI211_X1 port map( C1 => n39, C2 => n40, A => n41, B => n42, ZN => 
                           cout_4_port);
   U43 : OAI211_X1 port map( C1 => b(19), C2 => a(19), A => cout_3_port, B => 
                           n43, ZN => n42);
   U44 : AOI221_X1 port map( B1 => n44, B2 => n45, C1 => n46, C2 => n47, A => 
                           n48, ZN => n43);
   U45 : OAI21_X1 port map( B1 => n49, B2 => a(19), A => b(19), ZN => n41);
   U46 : INV_X1 port map( A => a(19), ZN => n40);
   U47 : INV_X1 port map( A => n49, ZN => n39);
   U48 : AOI21_X1 port map( B1 => n44, B2 => n50, A => n51, ZN => n49);
   U49 : INV_X1 port map( A => n52, ZN => n51);
   U50 : OAI21_X1 port map( B1 => n50, B2 => n44, A => n45, ZN => n52);
   U51 : INV_X1 port map( A => b(18), ZN => n45);
   U52 : AOI21_X1 port map( B1 => a(17), B2 => b(17), A => n53, ZN => n50);
   U53 : NOR3_X1 port map( A1 => n46, A2 => n48, A3 => n47, ZN => n53);
   U54 : INV_X1 port map( A => b(16), ZN => n47);
   U55 : NOR2_X1 port map( A1 => b(17), A2 => a(17), ZN => n48);
   U56 : INV_X1 port map( A => a(16), ZN => n46);
   U57 : INV_X1 port map( A => a(18), ZN => n44);
   U58 : INV_X1 port map( A => n54, ZN => cout_3_port);
   U59 : OAI22_X1 port map( A1 => a(15), A2 => n55, B1 => b(15), B2 => n56, ZN 
                           => n54);
   U60 : AND2_X1 port map( A1 => n55, A2 => a(15), ZN => n56);
   U61 : INV_X1 port map( A => n57, ZN => n55);
   U62 : OAI22_X1 port map( A1 => a(14), A2 => n58, B1 => b(14), B2 => n59, ZN 
                           => n57);
   U63 : AND2_X1 port map( A1 => n58, A2 => a(14), ZN => n59);
   U64 : OAI21_X1 port map( B1 => n60, B2 => n61, A => n62, ZN => n58);
   U65 : OAI21_X1 port map( B1 => b(13), B2 => a(13), A => n63, ZN => n62);
   U66 : INV_X1 port map( A => n64, ZN => n63);
   U67 : AOI21_X1 port map( B1 => cout_2_port, B2 => a(12), A => n65, ZN => n64
                           );
   U68 : INV_X1 port map( A => n66, ZN => n65);
   U69 : OAI21_X1 port map( B1 => a(12), B2 => cout_2_port, A => b(12), ZN => 
                           n66);
   U70 : INV_X1 port map( A => b(13), ZN => n61);
   U71 : INV_X1 port map( A => a(13), ZN => n60);
   U72 : OAI21_X1 port map( B1 => n67, B2 => n68, A => n69, ZN => cout_2_port);
   U73 : OAI21_X1 port map( B1 => a(11), B2 => n70, A => b(11), ZN => n69);
   U74 : INV_X1 port map( A => n67, ZN => n70);
   U75 : INV_X1 port map( A => a(11), ZN => n68);
   U76 : AOI21_X1 port map( B1 => a(10), B2 => b(10), A => n71, ZN => n67);
   U77 : INV_X1 port map( A => n72, ZN => n71);
   U78 : OAI22_X1 port map( A1 => n73, A2 => n74, B1 => a(10), B2 => b(10), ZN 
                           => n72);
   U79 : NOR2_X1 port map( A1 => n75, A2 => n76, ZN => n74);
   U80 : AOI22_X1 port map( A1 => n75, A2 => n76, B1 => n77, B2 => n78, ZN => 
                           n73);
   U81 : OAI21_X1 port map( B1 => a(8), B2 => cout_1_port, A => b(8), ZN => n78
                           );
   U82 : NAND2_X1 port map( A1 => a(8), A2 => cout_1_port, ZN => n77);
   U83 : INV_X1 port map( A => b(9), ZN => n76);
   U84 : INV_X1 port map( A => a(9), ZN => n75);
   U85 : OAI21_X1 port map( B1 => n79, B2 => n80, A => n81, ZN => cout_1_port);
   U86 : OAI21_X1 port map( B1 => b(7), B2 => a(7), A => n82, ZN => n81);
   U87 : OAI21_X1 port map( B1 => n83, B2 => n84, A => n85, ZN => n82);
   U88 : OAI21_X1 port map( B1 => a(6), B2 => n86, A => b(6), ZN => n85);
   U89 : INV_X1 port map( A => n83, ZN => n86);
   U90 : INV_X1 port map( A => a(6), ZN => n84);
   U91 : AOI22_X1 port map( A1 => a(5), A2 => b(5), B1 => n87, B2 => n88, ZN =>
                           n83);
   U92 : INV_X1 port map( A => n89, ZN => n88);
   U93 : AOI22_X1 port map( A1 => b(4), A2 => n90, B1 => a(4), B2 => 
                           cout_0_port, ZN => n89);
   U94 : OR2_X1 port map( A1 => a(4), A2 => cout_0_port, ZN => n90);
   U95 : OR2_X1 port map( A1 => b(5), A2 => a(5), ZN => n87);
   U96 : INV_X1 port map( A => b(7), ZN => n80);
   U97 : INV_X1 port map( A => a(7), ZN => n79);
   U98 : INV_X1 port map( A => n91, ZN => cout_0_port);
   U99 : OAI22_X1 port map( A1 => a(3), A2 => n92, B1 => b(3), B2 => n93, ZN =>
                           n91);
   U100 : AND2_X1 port map( A1 => n92, A2 => a(3), ZN => n93);
   U101 : INV_X1 port map( A => n94, ZN => n92);
   U102 : OAI22_X1 port map( A1 => a(2), A2 => n95, B1 => b(2), B2 => n96, ZN 
                           => n94);
   U103 : AND2_X1 port map( A1 => n95, A2 => a(2), ZN => n96);
   U104 : INV_X1 port map( A => n97, ZN => n95);
   U105 : AOI22_X1 port map( A1 => a(1), A2 => b(1), B1 => n98, B2 => n99, ZN 
                           => n97);
   U106 : INV_X1 port map( A => n100, ZN => n99);
   U107 : AOI22_X1 port map( A1 => cin, A2 => n101, B1 => b(0), B2 => a(0), ZN 
                           => n100);
   U108 : OR2_X1 port map( A1 => b(0), A2 => a(0), ZN => n101);
   U109 : OR2_X1 port map( A1 => b(1), A2 => a(1), ZN => n98);

end SYN_p4_carry_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AddSub_DATA_SIZE32_3 is

   port( as : in std_logic;  a, b : in std_logic_vector (31 downto 0);  re : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end AddSub_DATA_SIZE32_3;

architecture SYN_add_sub_arch of AddSub_DATA_SIZE32_3 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component Adder_DATA_SIZE32_3
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;
   
   signal b_new_31_port, b_new_30_port, b_new_29_port, b_new_28_port, 
      b_new_27_port, b_new_26_port, b_new_25_port, b_new_24_port, b_new_23_port
      , b_new_22_port, b_new_21_port, b_new_20_port, b_new_19_port, 
      b_new_18_port, b_new_17_port, b_new_16_port, b_new_15_port, b_new_14_port
      , b_new_13_port, b_new_12_port, b_new_11_port, b_new_10_port, 
      b_new_9_port, b_new_8_port, b_new_7_port, b_new_6_port, b_new_5_port, 
      b_new_4_port, b_new_3_port, b_new_2_port, b_new_1_port, b_new_0_port : 
      std_logic;

begin
   
   ADDER0 : Adder_DATA_SIZE32_3 port map( cin => as, a(31) => a(31), a(30) => 
                           a(30), a(29) => a(29), a(28) => a(28), a(27) => 
                           a(27), a(26) => a(26), a(25) => a(25), a(24) => 
                           a(24), a(23) => a(23), a(22) => a(22), a(21) => 
                           a(21), a(20) => a(20), a(19) => a(19), a(18) => 
                           a(18), a(17) => a(17), a(16) => a(16), a(15) => 
                           a(15), a(14) => a(14), a(13) => a(13), a(12) => 
                           a(12), a(11) => a(11), a(10) => a(10), a(9) => a(9),
                           a(8) => a(8), a(7) => a(7), a(6) => a(6), a(5) => 
                           a(5), a(4) => a(4), a(3) => a(3), a(2) => a(2), a(1)
                           => a(1), a(0) => a(0), b(31) => b_new_31_port, b(30)
                           => b_new_30_port, b(29) => b_new_29_port, b(28) => 
                           b_new_28_port, b(27) => b_new_27_port, b(26) => 
                           b_new_26_port, b(25) => b_new_25_port, b(24) => 
                           b_new_24_port, b(23) => b_new_23_port, b(22) => 
                           b_new_22_port, b(21) => b_new_21_port, b(20) => 
                           b_new_20_port, b(19) => b_new_19_port, b(18) => 
                           b_new_18_port, b(17) => b_new_17_port, b(16) => 
                           b_new_16_port, b(15) => b_new_15_port, b(14) => 
                           b_new_14_port, b(13) => b_new_13_port, b(12) => 
                           b_new_12_port, b(11) => b_new_11_port, b(10) => 
                           b_new_10_port, b(9) => b_new_9_port, b(8) => 
                           b_new_8_port, b(7) => b_new_7_port, b(6) => 
                           b_new_6_port, b(5) => b_new_5_port, b(4) => 
                           b_new_4_port, b(3) => b_new_3_port, b(2) => 
                           b_new_2_port, b(1) => b_new_1_port, b(0) => 
                           b_new_0_port, s(31) => re(31), s(30) => re(30), 
                           s(29) => re(29), s(28) => re(28), s(27) => re(27), 
                           s(26) => re(26), s(25) => re(25), s(24) => re(24), 
                           s(23) => re(23), s(22) => re(22), s(21) => re(21), 
                           s(20) => re(20), s(19) => re(19), s(18) => re(18), 
                           s(17) => re(17), s(16) => re(16), s(15) => re(15), 
                           s(14) => re(14), s(13) => re(13), s(12) => re(12), 
                           s(11) => re(11), s(10) => re(10), s(9) => re(9), 
                           s(8) => re(8), s(7) => re(7), s(6) => re(6), s(5) =>
                           re(5), s(4) => re(4), s(3) => re(3), s(2) => re(2), 
                           s(1) => re(1), s(0) => re(0), cout => cout);
   U1 : XOR2_X1 port map( A => b(9), B => as, Z => b_new_9_port);
   U2 : XOR2_X1 port map( A => b(8), B => as, Z => b_new_8_port);
   U3 : XOR2_X1 port map( A => b(7), B => as, Z => b_new_7_port);
   U4 : XOR2_X1 port map( A => b(6), B => as, Z => b_new_6_port);
   U5 : XOR2_X1 port map( A => b(5), B => as, Z => b_new_5_port);
   U6 : XOR2_X1 port map( A => b(4), B => as, Z => b_new_4_port);
   U7 : XOR2_X1 port map( A => b(3), B => as, Z => b_new_3_port);
   U8 : XOR2_X1 port map( A => b(31), B => as, Z => b_new_31_port);
   U9 : XOR2_X1 port map( A => b(30), B => as, Z => b_new_30_port);
   U10 : XOR2_X1 port map( A => b(2), B => as, Z => b_new_2_port);
   U11 : XOR2_X1 port map( A => b(29), B => as, Z => b_new_29_port);
   U12 : XOR2_X1 port map( A => b(28), B => as, Z => b_new_28_port);
   U13 : XOR2_X1 port map( A => b(27), B => as, Z => b_new_27_port);
   U14 : XOR2_X1 port map( A => b(26), B => as, Z => b_new_26_port);
   U15 : XOR2_X1 port map( A => b(25), B => as, Z => b_new_25_port);
   U16 : XOR2_X1 port map( A => b(24), B => as, Z => b_new_24_port);
   U17 : XOR2_X1 port map( A => b(23), B => as, Z => b_new_23_port);
   U18 : XOR2_X1 port map( A => b(22), B => as, Z => b_new_22_port);
   U19 : XOR2_X1 port map( A => b(21), B => as, Z => b_new_21_port);
   U20 : XOR2_X1 port map( A => b(20), B => as, Z => b_new_20_port);
   U21 : XOR2_X1 port map( A => b(1), B => as, Z => b_new_1_port);
   U22 : XOR2_X1 port map( A => b(19), B => as, Z => b_new_19_port);
   U23 : XOR2_X1 port map( A => b(18), B => as, Z => b_new_18_port);
   U24 : XOR2_X1 port map( A => b(17), B => as, Z => b_new_17_port);
   U25 : XOR2_X1 port map( A => b(16), B => as, Z => b_new_16_port);
   U26 : XOR2_X1 port map( A => b(15), B => as, Z => b_new_15_port);
   U27 : XOR2_X1 port map( A => b(14), B => as, Z => b_new_14_port);
   U28 : XOR2_X1 port map( A => b(13), B => as, Z => b_new_13_port);
   U29 : XOR2_X1 port map( A => b(12), B => as, Z => b_new_12_port);
   U30 : XOR2_X1 port map( A => b(11), B => as, Z => b_new_11_port);
   U31 : XOR2_X1 port map( A => b(10), B => as, Z => b_new_10_port);
   U32 : XOR2_X1 port map( A => b(0), B => as, Z => b_new_0_port);

end SYN_add_sub_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AddSub_DATA_SIZE32_2 is

   port( as : in std_logic;  a, b : in std_logic_vector (31 downto 0);  re : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end AddSub_DATA_SIZE32_2;

architecture SYN_add_sub_arch of AddSub_DATA_SIZE32_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component Adder_DATA_SIZE32_2
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;
   
   signal b_new_31_port, b_new_30_port, b_new_29_port, b_new_28_port, 
      b_new_27_port, b_new_26_port, b_new_25_port, b_new_24_port, b_new_23_port
      , b_new_22_port, b_new_21_port, b_new_20_port, b_new_19_port, 
      b_new_18_port, b_new_17_port, b_new_16_port, b_new_15_port, b_new_14_port
      , b_new_13_port, b_new_12_port, b_new_11_port, b_new_10_port, 
      b_new_9_port, b_new_8_port, b_new_7_port, b_new_6_port, b_new_5_port, 
      b_new_4_port, b_new_3_port, b_new_2_port, b_new_1_port, b_new_0_port : 
      std_logic;

begin
   
   ADDER0 : Adder_DATA_SIZE32_2 port map( cin => as, a(31) => a(31), a(30) => 
                           a(30), a(29) => a(29), a(28) => a(28), a(27) => 
                           a(27), a(26) => a(26), a(25) => a(25), a(24) => 
                           a(24), a(23) => a(23), a(22) => a(22), a(21) => 
                           a(21), a(20) => a(20), a(19) => a(19), a(18) => 
                           a(18), a(17) => a(17), a(16) => a(16), a(15) => 
                           a(15), a(14) => a(14), a(13) => a(13), a(12) => 
                           a(12), a(11) => a(11), a(10) => a(10), a(9) => a(9),
                           a(8) => a(8), a(7) => a(7), a(6) => a(6), a(5) => 
                           a(5), a(4) => a(4), a(3) => a(3), a(2) => a(2), a(1)
                           => a(1), a(0) => a(0), b(31) => b_new_31_port, b(30)
                           => b_new_30_port, b(29) => b_new_29_port, b(28) => 
                           b_new_28_port, b(27) => b_new_27_port, b(26) => 
                           b_new_26_port, b(25) => b_new_25_port, b(24) => 
                           b_new_24_port, b(23) => b_new_23_port, b(22) => 
                           b_new_22_port, b(21) => b_new_21_port, b(20) => 
                           b_new_20_port, b(19) => b_new_19_port, b(18) => 
                           b_new_18_port, b(17) => b_new_17_port, b(16) => 
                           b_new_16_port, b(15) => b_new_15_port, b(14) => 
                           b_new_14_port, b(13) => b_new_13_port, b(12) => 
                           b_new_12_port, b(11) => b_new_11_port, b(10) => 
                           b_new_10_port, b(9) => b_new_9_port, b(8) => 
                           b_new_8_port, b(7) => b_new_7_port, b(6) => 
                           b_new_6_port, b(5) => b_new_5_port, b(4) => 
                           b_new_4_port, b(3) => b_new_3_port, b(2) => 
                           b_new_2_port, b(1) => b_new_1_port, b(0) => 
                           b_new_0_port, s(31) => re(31), s(30) => re(30), 
                           s(29) => re(29), s(28) => re(28), s(27) => re(27), 
                           s(26) => re(26), s(25) => re(25), s(24) => re(24), 
                           s(23) => re(23), s(22) => re(22), s(21) => re(21), 
                           s(20) => re(20), s(19) => re(19), s(18) => re(18), 
                           s(17) => re(17), s(16) => re(16), s(15) => re(15), 
                           s(14) => re(14), s(13) => re(13), s(12) => re(12), 
                           s(11) => re(11), s(10) => re(10), s(9) => re(9), 
                           s(8) => re(8), s(7) => re(7), s(6) => re(6), s(5) =>
                           re(5), s(4) => re(4), s(3) => re(3), s(2) => re(2), 
                           s(1) => re(1), s(0) => re(0), cout => cout);
   U1 : XOR2_X1 port map( A => b(9), B => as, Z => b_new_9_port);
   U2 : XOR2_X1 port map( A => b(8), B => as, Z => b_new_8_port);
   U3 : XOR2_X1 port map( A => b(7), B => as, Z => b_new_7_port);
   U4 : XOR2_X1 port map( A => b(6), B => as, Z => b_new_6_port);
   U5 : XOR2_X1 port map( A => b(5), B => as, Z => b_new_5_port);
   U6 : XOR2_X1 port map( A => b(4), B => as, Z => b_new_4_port);
   U7 : XOR2_X1 port map( A => b(3), B => as, Z => b_new_3_port);
   U8 : XOR2_X1 port map( A => b(31), B => as, Z => b_new_31_port);
   U9 : XOR2_X1 port map( A => b(30), B => as, Z => b_new_30_port);
   U10 : XOR2_X1 port map( A => b(2), B => as, Z => b_new_2_port);
   U11 : XOR2_X1 port map( A => b(29), B => as, Z => b_new_29_port);
   U12 : XOR2_X1 port map( A => b(28), B => as, Z => b_new_28_port);
   U13 : XOR2_X1 port map( A => b(27), B => as, Z => b_new_27_port);
   U14 : XOR2_X1 port map( A => b(26), B => as, Z => b_new_26_port);
   U15 : XOR2_X1 port map( A => b(25), B => as, Z => b_new_25_port);
   U16 : XOR2_X1 port map( A => b(24), B => as, Z => b_new_24_port);
   U17 : XOR2_X1 port map( A => b(23), B => as, Z => b_new_23_port);
   U18 : XOR2_X1 port map( A => b(22), B => as, Z => b_new_22_port);
   U19 : XOR2_X1 port map( A => b(21), B => as, Z => b_new_21_port);
   U20 : XOR2_X1 port map( A => b(20), B => as, Z => b_new_20_port);
   U21 : XOR2_X1 port map( A => b(1), B => as, Z => b_new_1_port);
   U22 : XOR2_X1 port map( A => b(19), B => as, Z => b_new_19_port);
   U23 : XOR2_X1 port map( A => b(18), B => as, Z => b_new_18_port);
   U24 : XOR2_X1 port map( A => b(17), B => as, Z => b_new_17_port);
   U25 : XOR2_X1 port map( A => b(16), B => as, Z => b_new_16_port);
   U26 : XOR2_X1 port map( A => b(15), B => as, Z => b_new_15_port);
   U27 : XOR2_X1 port map( A => b(14), B => as, Z => b_new_14_port);
   U28 : XOR2_X1 port map( A => b(13), B => as, Z => b_new_13_port);
   U29 : XOR2_X1 port map( A => b(12), B => as, Z => b_new_12_port);
   U30 : XOR2_X1 port map( A => b(11), B => as, Z => b_new_11_port);
   U31 : XOR2_X1 port map( A => b(10), B => as, Z => b_new_10_port);
   U32 : XOR2_X1 port map( A => b(0), B => as, Z => b_new_0_port);

end SYN_add_sub_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AddSub_DATA_SIZE32_1 is

   port( as : in std_logic;  a, b : in std_logic_vector (31 downto 0);  re : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end AddSub_DATA_SIZE32_1;

architecture SYN_add_sub_arch of AddSub_DATA_SIZE32_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component Adder_DATA_SIZE32_1
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;
   
   signal b_new_31_port, b_new_30_port, b_new_29_port, b_new_28_port, 
      b_new_27_port, b_new_26_port, b_new_25_port, b_new_24_port, b_new_23_port
      , b_new_22_port, b_new_21_port, b_new_20_port, b_new_19_port, 
      b_new_18_port, b_new_17_port, b_new_16_port, b_new_15_port, b_new_14_port
      , b_new_13_port, b_new_12_port, b_new_11_port, b_new_10_port, 
      b_new_9_port, b_new_8_port, b_new_7_port, b_new_6_port, b_new_5_port, 
      b_new_4_port, b_new_3_port, b_new_2_port, b_new_1_port, b_new_0_port : 
      std_logic;

begin
   
   ADDER0 : Adder_DATA_SIZE32_1 port map( cin => as, a(31) => a(31), a(30) => 
                           a(30), a(29) => a(29), a(28) => a(28), a(27) => 
                           a(27), a(26) => a(26), a(25) => a(25), a(24) => 
                           a(24), a(23) => a(23), a(22) => a(22), a(21) => 
                           a(21), a(20) => a(20), a(19) => a(19), a(18) => 
                           a(18), a(17) => a(17), a(16) => a(16), a(15) => 
                           a(15), a(14) => a(14), a(13) => a(13), a(12) => 
                           a(12), a(11) => a(11), a(10) => a(10), a(9) => a(9),
                           a(8) => a(8), a(7) => a(7), a(6) => a(6), a(5) => 
                           a(5), a(4) => a(4), a(3) => a(3), a(2) => a(2), a(1)
                           => a(1), a(0) => a(0), b(31) => b_new_31_port, b(30)
                           => b_new_30_port, b(29) => b_new_29_port, b(28) => 
                           b_new_28_port, b(27) => b_new_27_port, b(26) => 
                           b_new_26_port, b(25) => b_new_25_port, b(24) => 
                           b_new_24_port, b(23) => b_new_23_port, b(22) => 
                           b_new_22_port, b(21) => b_new_21_port, b(20) => 
                           b_new_20_port, b(19) => b_new_19_port, b(18) => 
                           b_new_18_port, b(17) => b_new_17_port, b(16) => 
                           b_new_16_port, b(15) => b_new_15_port, b(14) => 
                           b_new_14_port, b(13) => b_new_13_port, b(12) => 
                           b_new_12_port, b(11) => b_new_11_port, b(10) => 
                           b_new_10_port, b(9) => b_new_9_port, b(8) => 
                           b_new_8_port, b(7) => b_new_7_port, b(6) => 
                           b_new_6_port, b(5) => b_new_5_port, b(4) => 
                           b_new_4_port, b(3) => b_new_3_port, b(2) => 
                           b_new_2_port, b(1) => b_new_1_port, b(0) => 
                           b_new_0_port, s(31) => re(31), s(30) => re(30), 
                           s(29) => re(29), s(28) => re(28), s(27) => re(27), 
                           s(26) => re(26), s(25) => re(25), s(24) => re(24), 
                           s(23) => re(23), s(22) => re(22), s(21) => re(21), 
                           s(20) => re(20), s(19) => re(19), s(18) => re(18), 
                           s(17) => re(17), s(16) => re(16), s(15) => re(15), 
                           s(14) => re(14), s(13) => re(13), s(12) => re(12), 
                           s(11) => re(11), s(10) => re(10), s(9) => re(9), 
                           s(8) => re(8), s(7) => re(7), s(6) => re(6), s(5) =>
                           re(5), s(4) => re(4), s(3) => re(3), s(2) => re(2), 
                           s(1) => re(1), s(0) => re(0), cout => cout);
   U1 : XOR2_X1 port map( A => b(9), B => as, Z => b_new_9_port);
   U2 : XOR2_X1 port map( A => b(8), B => as, Z => b_new_8_port);
   U3 : XOR2_X1 port map( A => b(7), B => as, Z => b_new_7_port);
   U4 : XOR2_X1 port map( A => b(6), B => as, Z => b_new_6_port);
   U5 : XOR2_X1 port map( A => b(5), B => as, Z => b_new_5_port);
   U6 : XOR2_X1 port map( A => b(4), B => as, Z => b_new_4_port);
   U7 : XOR2_X1 port map( A => b(3), B => as, Z => b_new_3_port);
   U8 : XOR2_X1 port map( A => b(31), B => as, Z => b_new_31_port);
   U9 : XOR2_X1 port map( A => b(30), B => as, Z => b_new_30_port);
   U10 : XOR2_X1 port map( A => b(2), B => as, Z => b_new_2_port);
   U11 : XOR2_X1 port map( A => b(29), B => as, Z => b_new_29_port);
   U12 : XOR2_X1 port map( A => b(28), B => as, Z => b_new_28_port);
   U13 : XOR2_X1 port map( A => b(27), B => as, Z => b_new_27_port);
   U14 : XOR2_X1 port map( A => b(26), B => as, Z => b_new_26_port);
   U15 : XOR2_X1 port map( A => b(25), B => as, Z => b_new_25_port);
   U16 : XOR2_X1 port map( A => b(24), B => as, Z => b_new_24_port);
   U17 : XOR2_X1 port map( A => b(23), B => as, Z => b_new_23_port);
   U18 : XOR2_X1 port map( A => b(22), B => as, Z => b_new_22_port);
   U19 : XOR2_X1 port map( A => b(21), B => as, Z => b_new_21_port);
   U20 : XOR2_X1 port map( A => b(20), B => as, Z => b_new_20_port);
   U21 : XOR2_X1 port map( A => b(1), B => as, Z => b_new_1_port);
   U22 : XOR2_X1 port map( A => b(19), B => as, Z => b_new_19_port);
   U23 : XOR2_X1 port map( A => b(18), B => as, Z => b_new_18_port);
   U24 : XOR2_X1 port map( A => b(17), B => as, Z => b_new_17_port);
   U25 : XOR2_X1 port map( A => b(16), B => as, Z => b_new_16_port);
   U26 : XOR2_X1 port map( A => b(15), B => as, Z => b_new_15_port);
   U27 : XOR2_X1 port map( A => b(14), B => as, Z => b_new_14_port);
   U28 : XOR2_X1 port map( A => b(13), B => as, Z => b_new_13_port);
   U29 : XOR2_X1 port map( A => b(12), B => as, Z => b_new_12_port);
   U30 : XOR2_X1 port map( A => b(11), B => as, Z => b_new_11_port);
   U31 : XOR2_X1 port map( A => b(10), B => as, Z => b_new_10_port);
   U32 : XOR2_X1 port map( A => b(0), B => as, Z => b_new_0_port);

end SYN_add_sub_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4Adder_DATA_SIZE32_SPARSITY4_7 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end P4Adder_DATA_SIZE32_SPARSITY4_7;

architecture SYN_p4_adder_arch of P4Adder_DATA_SIZE32_SPARSITY4_7 is

   component AdderSumGenerator_DATA_SIZE32_SPARSITY4_7
      port( a, b : in std_logic_vector (31 downto 0);  cin : in 
            std_logic_vector (7 downto 0);  sum : out std_logic_vector (31 
            downto 0));
   end component;
   
   component P4CarryGenerator_DATA_SIZE32_SPARSITY4_7
      port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  
            cout : out std_logic_vector (7 downto 0));
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, carry_1_port : std_logic;

begin
   
   CG0 : P4CarryGenerator_DATA_SIZE32_SPARSITY4_7 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), cin => cin, 
                           cout(7) => cout, cout(6) => carry_7_port, cout(5) =>
                           carry_6_port, cout(4) => carry_5_port, cout(3) => 
                           carry_4_port, cout(2) => carry_3_port, cout(1) => 
                           carry_2_port, cout(0) => carry_1_port);
   SG0 : AdderSumGenerator_DATA_SIZE32_SPARSITY4_7 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), cin(7) => 
                           carry_7_port, cin(6) => carry_6_port, cin(5) => 
                           carry_5_port, cin(4) => carry_4_port, cin(3) => 
                           carry_3_port, cin(2) => carry_2_port, cin(1) => 
                           carry_1_port, cin(0) => cin, sum(31) => s(31), 
                           sum(30) => s(30), sum(29) => s(29), sum(28) => s(28)
                           , sum(27) => s(27), sum(26) => s(26), sum(25) => 
                           s(25), sum(24) => s(24), sum(23) => s(23), sum(22) 
                           => s(22), sum(21) => s(21), sum(20) => s(20), 
                           sum(19) => s(19), sum(18) => s(18), sum(17) => s(17)
                           , sum(16) => s(16), sum(15) => s(15), sum(14) => 
                           s(14), sum(13) => s(13), sum(12) => s(12), sum(11) 
                           => s(11), sum(10) => s(10), sum(9) => s(9), sum(8) 
                           => s(8), sum(7) => s(7), sum(6) => s(6), sum(5) => 
                           s(5), sum(4) => s(4), sum(3) => s(3), sum(2) => s(2)
                           , sum(1) => s(1), sum(0) => s(0));

end SYN_p4_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4Adder_DATA_SIZE32_SPARSITY4_6 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end P4Adder_DATA_SIZE32_SPARSITY4_6;

architecture SYN_p4_adder_arch of P4Adder_DATA_SIZE32_SPARSITY4_6 is

   component AdderSumGenerator_DATA_SIZE32_SPARSITY4_6
      port( a, b : in std_logic_vector (31 downto 0);  cin : in 
            std_logic_vector (7 downto 0);  sum : out std_logic_vector (31 
            downto 0));
   end component;
   
   component P4CarryGenerator_DATA_SIZE32_SPARSITY4_6
      port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  
            cout : out std_logic_vector (7 downto 0));
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, carry_1_port : std_logic;

begin
   
   CG0 : P4CarryGenerator_DATA_SIZE32_SPARSITY4_6 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), cin => cin, 
                           cout(7) => cout, cout(6) => carry_7_port, cout(5) =>
                           carry_6_port, cout(4) => carry_5_port, cout(3) => 
                           carry_4_port, cout(2) => carry_3_port, cout(1) => 
                           carry_2_port, cout(0) => carry_1_port);
   SG0 : AdderSumGenerator_DATA_SIZE32_SPARSITY4_6 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), cin(7) => 
                           carry_7_port, cin(6) => carry_6_port, cin(5) => 
                           carry_5_port, cin(4) => carry_4_port, cin(3) => 
                           carry_3_port, cin(2) => carry_2_port, cin(1) => 
                           carry_1_port, cin(0) => cin, sum(31) => s(31), 
                           sum(30) => s(30), sum(29) => s(29), sum(28) => s(28)
                           , sum(27) => s(27), sum(26) => s(26), sum(25) => 
                           s(25), sum(24) => s(24), sum(23) => s(23), sum(22) 
                           => s(22), sum(21) => s(21), sum(20) => s(20), 
                           sum(19) => s(19), sum(18) => s(18), sum(17) => s(17)
                           , sum(16) => s(16), sum(15) => s(15), sum(14) => 
                           s(14), sum(13) => s(13), sum(12) => s(12), sum(11) 
                           => s(11), sum(10) => s(10), sum(9) => s(9), sum(8) 
                           => s(8), sum(7) => s(7), sum(6) => s(6), sum(5) => 
                           s(5), sum(4) => s(4), sum(3) => s(3), sum(2) => s(2)
                           , sum(1) => s(1), sum(0) => s(0));

end SYN_p4_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4Adder_DATA_SIZE32_SPARSITY4_5 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end P4Adder_DATA_SIZE32_SPARSITY4_5;

architecture SYN_p4_adder_arch of P4Adder_DATA_SIZE32_SPARSITY4_5 is

   component AdderSumGenerator_DATA_SIZE32_SPARSITY4_5
      port( a, b : in std_logic_vector (31 downto 0);  cin : in 
            std_logic_vector (7 downto 0);  sum : out std_logic_vector (31 
            downto 0));
   end component;
   
   component P4CarryGenerator_DATA_SIZE32_SPARSITY4_5
      port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  
            cout : out std_logic_vector (7 downto 0));
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, carry_1_port : std_logic;

begin
   
   CG0 : P4CarryGenerator_DATA_SIZE32_SPARSITY4_5 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), cin => cin, 
                           cout(7) => cout, cout(6) => carry_7_port, cout(5) =>
                           carry_6_port, cout(4) => carry_5_port, cout(3) => 
                           carry_4_port, cout(2) => carry_3_port, cout(1) => 
                           carry_2_port, cout(0) => carry_1_port);
   SG0 : AdderSumGenerator_DATA_SIZE32_SPARSITY4_5 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), cin(7) => 
                           carry_7_port, cin(6) => carry_6_port, cin(5) => 
                           carry_5_port, cin(4) => carry_4_port, cin(3) => 
                           carry_3_port, cin(2) => carry_2_port, cin(1) => 
                           carry_1_port, cin(0) => cin, sum(31) => s(31), 
                           sum(30) => s(30), sum(29) => s(29), sum(28) => s(28)
                           , sum(27) => s(27), sum(26) => s(26), sum(25) => 
                           s(25), sum(24) => s(24), sum(23) => s(23), sum(22) 
                           => s(22), sum(21) => s(21), sum(20) => s(20), 
                           sum(19) => s(19), sum(18) => s(18), sum(17) => s(17)
                           , sum(16) => s(16), sum(15) => s(15), sum(14) => 
                           s(14), sum(13) => s(13), sum(12) => s(12), sum(11) 
                           => s(11), sum(10) => s(10), sum(9) => s(9), sum(8) 
                           => s(8), sum(7) => s(7), sum(6) => s(6), sum(5) => 
                           s(5), sum(4) => s(4), sum(3) => s(3), sum(2) => s(2)
                           , sum(1) => s(1), sum(0) => s(0));

end SYN_p4_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4Adder_DATA_SIZE32_SPARSITY4_4 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end P4Adder_DATA_SIZE32_SPARSITY4_4;

architecture SYN_p4_adder_arch of P4Adder_DATA_SIZE32_SPARSITY4_4 is

   component AdderSumGenerator_DATA_SIZE32_SPARSITY4_4
      port( a, b : in std_logic_vector (31 downto 0);  cin : in 
            std_logic_vector (7 downto 0);  sum : out std_logic_vector (31 
            downto 0));
   end component;
   
   component P4CarryGenerator_DATA_SIZE32_SPARSITY4_4
      port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  
            cout : out std_logic_vector (7 downto 0));
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, carry_1_port : std_logic;

begin
   
   CG0 : P4CarryGenerator_DATA_SIZE32_SPARSITY4_4 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), cin => cin, 
                           cout(7) => cout, cout(6) => carry_7_port, cout(5) =>
                           carry_6_port, cout(4) => carry_5_port, cout(3) => 
                           carry_4_port, cout(2) => carry_3_port, cout(1) => 
                           carry_2_port, cout(0) => carry_1_port);
   SG0 : AdderSumGenerator_DATA_SIZE32_SPARSITY4_4 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), cin(7) => 
                           carry_7_port, cin(6) => carry_6_port, cin(5) => 
                           carry_5_port, cin(4) => carry_4_port, cin(3) => 
                           carry_3_port, cin(2) => carry_2_port, cin(1) => 
                           carry_1_port, cin(0) => cin, sum(31) => s(31), 
                           sum(30) => s(30), sum(29) => s(29), sum(28) => s(28)
                           , sum(27) => s(27), sum(26) => s(26), sum(25) => 
                           s(25), sum(24) => s(24), sum(23) => s(23), sum(22) 
                           => s(22), sum(21) => s(21), sum(20) => s(20), 
                           sum(19) => s(19), sum(18) => s(18), sum(17) => s(17)
                           , sum(16) => s(16), sum(15) => s(15), sum(14) => 
                           s(14), sum(13) => s(13), sum(12) => s(12), sum(11) 
                           => s(11), sum(10) => s(10), sum(9) => s(9), sum(8) 
                           => s(8), sum(7) => s(7), sum(6) => s(6), sum(5) => 
                           s(5), sum(4) => s(4), sum(3) => s(3), sum(2) => s(2)
                           , sum(1) => s(1), sum(0) => s(0));

end SYN_p4_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4Adder_DATA_SIZE32_SPARSITY4_3 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end P4Adder_DATA_SIZE32_SPARSITY4_3;

architecture SYN_p4_adder_arch of P4Adder_DATA_SIZE32_SPARSITY4_3 is

   component AdderSumGenerator_DATA_SIZE32_SPARSITY4_3
      port( a, b : in std_logic_vector (31 downto 0);  cin : in 
            std_logic_vector (7 downto 0);  sum : out std_logic_vector (31 
            downto 0));
   end component;
   
   component P4CarryGenerator_DATA_SIZE32_SPARSITY4_3
      port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  
            cout : out std_logic_vector (7 downto 0));
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, carry_1_port : std_logic;

begin
   
   CG0 : P4CarryGenerator_DATA_SIZE32_SPARSITY4_3 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), cin => cin, 
                           cout(7) => cout, cout(6) => carry_7_port, cout(5) =>
                           carry_6_port, cout(4) => carry_5_port, cout(3) => 
                           carry_4_port, cout(2) => carry_3_port, cout(1) => 
                           carry_2_port, cout(0) => carry_1_port);
   SG0 : AdderSumGenerator_DATA_SIZE32_SPARSITY4_3 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), cin(7) => 
                           carry_7_port, cin(6) => carry_6_port, cin(5) => 
                           carry_5_port, cin(4) => carry_4_port, cin(3) => 
                           carry_3_port, cin(2) => carry_2_port, cin(1) => 
                           carry_1_port, cin(0) => cin, sum(31) => s(31), 
                           sum(30) => s(30), sum(29) => s(29), sum(28) => s(28)
                           , sum(27) => s(27), sum(26) => s(26), sum(25) => 
                           s(25), sum(24) => s(24), sum(23) => s(23), sum(22) 
                           => s(22), sum(21) => s(21), sum(20) => s(20), 
                           sum(19) => s(19), sum(18) => s(18), sum(17) => s(17)
                           , sum(16) => s(16), sum(15) => s(15), sum(14) => 
                           s(14), sum(13) => s(13), sum(12) => s(12), sum(11) 
                           => s(11), sum(10) => s(10), sum(9) => s(9), sum(8) 
                           => s(8), sum(7) => s(7), sum(6) => s(6), sum(5) => 
                           s(5), sum(4) => s(4), sum(3) => s(3), sum(2) => s(2)
                           , sum(1) => s(1), sum(0) => s(0));

end SYN_p4_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4Adder_DATA_SIZE32_SPARSITY4_2 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end P4Adder_DATA_SIZE32_SPARSITY4_2;

architecture SYN_p4_adder_arch of P4Adder_DATA_SIZE32_SPARSITY4_2 is

   component AdderSumGenerator_DATA_SIZE32_SPARSITY4_2
      port( a, b : in std_logic_vector (31 downto 0);  cin : in 
            std_logic_vector (7 downto 0);  sum : out std_logic_vector (31 
            downto 0));
   end component;
   
   component P4CarryGenerator_DATA_SIZE32_SPARSITY4_2
      port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  
            cout : out std_logic_vector (7 downto 0));
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, carry_1_port : std_logic;

begin
   
   CG0 : P4CarryGenerator_DATA_SIZE32_SPARSITY4_2 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), cin => cin, 
                           cout(7) => cout, cout(6) => carry_7_port, cout(5) =>
                           carry_6_port, cout(4) => carry_5_port, cout(3) => 
                           carry_4_port, cout(2) => carry_3_port, cout(1) => 
                           carry_2_port, cout(0) => carry_1_port);
   SG0 : AdderSumGenerator_DATA_SIZE32_SPARSITY4_2 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), cin(7) => 
                           carry_7_port, cin(6) => carry_6_port, cin(5) => 
                           carry_5_port, cin(4) => carry_4_port, cin(3) => 
                           carry_3_port, cin(2) => carry_2_port, cin(1) => 
                           carry_1_port, cin(0) => cin, sum(31) => s(31), 
                           sum(30) => s(30), sum(29) => s(29), sum(28) => s(28)
                           , sum(27) => s(27), sum(26) => s(26), sum(25) => 
                           s(25), sum(24) => s(24), sum(23) => s(23), sum(22) 
                           => s(22), sum(21) => s(21), sum(20) => s(20), 
                           sum(19) => s(19), sum(18) => s(18), sum(17) => s(17)
                           , sum(16) => s(16), sum(15) => s(15), sum(14) => 
                           s(14), sum(13) => s(13), sum(12) => s(12), sum(11) 
                           => s(11), sum(10) => s(10), sum(9) => s(9), sum(8) 
                           => s(8), sum(7) => s(7), sum(6) => s(6), sum(5) => 
                           s(5), sum(4) => s(4), sum(3) => s(3), sum(2) => s(2)
                           , sum(1) => s(1), sum(0) => s(0));

end SYN_p4_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4Adder_DATA_SIZE32_SPARSITY4_1 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end P4Adder_DATA_SIZE32_SPARSITY4_1;

architecture SYN_p4_adder_arch of P4Adder_DATA_SIZE32_SPARSITY4_1 is

   component AdderSumGenerator_DATA_SIZE32_SPARSITY4_1
      port( a, b : in std_logic_vector (31 downto 0);  cin : in 
            std_logic_vector (7 downto 0);  sum : out std_logic_vector (31 
            downto 0));
   end component;
   
   component P4CarryGenerator_DATA_SIZE32_SPARSITY4_1
      port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  
            cout : out std_logic_vector (7 downto 0));
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, carry_1_port : std_logic;

begin
   
   CG0 : P4CarryGenerator_DATA_SIZE32_SPARSITY4_1 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), cin => cin, 
                           cout(7) => cout, cout(6) => carry_7_port, cout(5) =>
                           carry_6_port, cout(4) => carry_5_port, cout(3) => 
                           carry_4_port, cout(2) => carry_3_port, cout(1) => 
                           carry_2_port, cout(0) => carry_1_port);
   SG0 : AdderSumGenerator_DATA_SIZE32_SPARSITY4_1 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), cin(7) => 
                           carry_7_port, cin(6) => carry_6_port, cin(5) => 
                           carry_5_port, cin(4) => carry_4_port, cin(3) => 
                           carry_3_port, cin(2) => carry_2_port, cin(1) => 
                           carry_1_port, cin(0) => cin, sum(31) => s(31), 
                           sum(30) => s(30), sum(29) => s(29), sum(28) => s(28)
                           , sum(27) => s(27), sum(26) => s(26), sum(25) => 
                           s(25), sum(24) => s(24), sum(23) => s(23), sum(22) 
                           => s(22), sum(21) => s(21), sum(20) => s(20), 
                           sum(19) => s(19), sum(18) => s(18), sum(17) => s(17)
                           , sum(16) => s(16), sum(15) => s(15), sum(14) => 
                           s(14), sum(13) => s(13), sum(12) => s(12), sum(11) 
                           => s(11), sum(10) => s(10), sum(9) => s(9), sum(8) 
                           => s(8), sum(7) => s(7), sum(6) => s(6), sum(5) => 
                           s(5), sum(4) => s(4), sum(3) => s(3), sum(2) => s(2)
                           , sum(1) => s(1), sum(0) => s(0));

end SYN_p4_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE5_6 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 0); 
         dout : out std_logic_vector (4 downto 0));

end Reg_DATA_SIZE5_6;

architecture SYN_reg_arch of Reg_DATA_SIZE5_6 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal dout_4_port, dout_3_port, dout_2_port, dout_1_port, dout_0_port, n1, 
      n2, n3, n4, n5, net109218, net109219, net109220, net109221, net109222 : 
      std_logic;

begin
   dout <= ( dout_4_port, dout_3_port, dout_2_port, dout_1_port, dout_0_port );
   
   dout_reg_4_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           dout_4_port, QN => net109222);
   dout_reg_3_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           dout_3_port, QN => net109221);
   dout_reg_2_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           dout_2_port, QN => net109220);
   dout_reg_1_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           dout_1_port, QN => net109219);
   dout_reg_0_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           dout_0_port, QN => net109218);
   U2 : MUX2_X1 port map( A => dout_4_port, B => din(4), S => en, Z => n1);
   U3 : MUX2_X1 port map( A => dout_3_port, B => din(3), S => en, Z => n2);
   U4 : MUX2_X1 port map( A => dout_2_port, B => din(2), S => en, Z => n3);
   U5 : MUX2_X1 port map( A => dout_1_port, B => din(1), S => en, Z => n4);
   U6 : MUX2_X1 port map( A => dout_0_port, B => din(0), S => en, Z => n5);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE5_5 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 0); 
         dout : out std_logic_vector (4 downto 0));

end Reg_DATA_SIZE5_5;

architecture SYN_reg_arch of Reg_DATA_SIZE5_5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal dout_4_port, dout_3_port, dout_2_port, dout_1_port, dout_0_port, n1, 
      n2, n3, n4, n5, net109213, net109214, net109215, net109216, net109217 : 
      std_logic;

begin
   dout <= ( dout_4_port, dout_3_port, dout_2_port, dout_1_port, dout_0_port );
   
   dout_reg_4_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           dout_4_port, QN => net109217);
   dout_reg_3_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           dout_3_port, QN => net109216);
   dout_reg_2_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           dout_2_port, QN => net109215);
   dout_reg_1_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           dout_1_port, QN => net109214);
   dout_reg_0_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           dout_0_port, QN => net109213);
   U2 : MUX2_X1 port map( A => dout_4_port, B => din(4), S => en, Z => n1);
   U3 : MUX2_X1 port map( A => dout_3_port, B => din(3), S => en, Z => n2);
   U4 : MUX2_X1 port map( A => dout_2_port, B => din(2), S => en, Z => n3);
   U5 : MUX2_X1 port map( A => dout_1_port, B => din(1), S => en, Z => n4);
   U6 : MUX2_X1 port map( A => dout_0_port, B => din(0), S => en, Z => n5);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE5_4 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 0); 
         dout : out std_logic_vector (4 downto 0));

end Reg_DATA_SIZE5_4;

architecture SYN_reg_arch of Reg_DATA_SIZE5_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal dout_4_port, dout_3_port, dout_2_port, dout_1_port, dout_0_port, n1, 
      n2, n3, n4, n5, net109208, net109209, net109210, net109211, net109212 : 
      std_logic;

begin
   dout <= ( dout_4_port, dout_3_port, dout_2_port, dout_1_port, dout_0_port );
   
   dout_reg_4_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           dout_4_port, QN => net109212);
   dout_reg_3_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           dout_3_port, QN => net109211);
   dout_reg_2_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           dout_2_port, QN => net109210);
   dout_reg_1_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           dout_1_port, QN => net109209);
   dout_reg_0_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           dout_0_port, QN => net109208);
   U2 : MUX2_X1 port map( A => dout_4_port, B => din(4), S => en, Z => n1);
   U3 : MUX2_X1 port map( A => dout_3_port, B => din(3), S => en, Z => n2);
   U4 : MUX2_X1 port map( A => dout_2_port, B => din(2), S => en, Z => n3);
   U5 : MUX2_X1 port map( A => dout_1_port, B => din(1), S => en, Z => n4);
   U6 : MUX2_X1 port map( A => dout_0_port, B => din(0), S => en, Z => n5);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE5_3 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 0); 
         dout : out std_logic_vector (4 downto 0));

end Reg_DATA_SIZE5_3;

architecture SYN_reg_arch of Reg_DATA_SIZE5_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal dout_4_port, dout_3_port, dout_2_port, dout_1_port, dout_0_port, n1, 
      n2, n3, n4, n5, net109203, net109204, net109205, net109206, net109207 : 
      std_logic;

begin
   dout <= ( dout_4_port, dout_3_port, dout_2_port, dout_1_port, dout_0_port );
   
   dout_reg_4_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           dout_4_port, QN => net109207);
   dout_reg_3_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           dout_3_port, QN => net109206);
   dout_reg_2_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           dout_2_port, QN => net109205);
   dout_reg_1_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           dout_1_port, QN => net109204);
   dout_reg_0_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           dout_0_port, QN => net109203);
   U2 : MUX2_X1 port map( A => dout_4_port, B => din(4), S => en, Z => n1);
   U3 : MUX2_X1 port map( A => dout_3_port, B => din(3), S => en, Z => n2);
   U4 : MUX2_X1 port map( A => dout_2_port, B => din(2), S => en, Z => n3);
   U5 : MUX2_X1 port map( A => dout_1_port, B => din(1), S => en, Z => n4);
   U6 : MUX2_X1 port map( A => dout_0_port, B => din(0), S => en, Z => n5);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE5_2 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 0); 
         dout : out std_logic_vector (4 downto 0));

end Reg_DATA_SIZE5_2;

architecture SYN_reg_arch of Reg_DATA_SIZE5_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal dout_4_port, dout_3_port, dout_2_port, dout_1_port, dout_0_port, n1, 
      n2, n3, n4, n5, net109198, net109199, net109200, net109201, net109202 : 
      std_logic;

begin
   dout <= ( dout_4_port, dout_3_port, dout_2_port, dout_1_port, dout_0_port );
   
   dout_reg_4_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           dout_4_port, QN => net109202);
   dout_reg_3_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           dout_3_port, QN => net109201);
   dout_reg_2_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           dout_2_port, QN => net109200);
   dout_reg_1_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           dout_1_port, QN => net109199);
   dout_reg_0_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           dout_0_port, QN => net109198);
   U2 : MUX2_X1 port map( A => dout_4_port, B => din(4), S => en, Z => n1);
   U3 : MUX2_X1 port map( A => dout_3_port, B => din(3), S => en, Z => n2);
   U4 : MUX2_X1 port map( A => dout_2_port, B => din(2), S => en, Z => n3);
   U5 : MUX2_X1 port map( A => dout_1_port, B => din(1), S => en, Z => n4);
   U6 : MUX2_X1 port map( A => dout_0_port, B => din(0), S => en, Z => n5);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE5_1 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 0); 
         dout : out std_logic_vector (4 downto 0));

end Reg_DATA_SIZE5_1;

architecture SYN_reg_arch of Reg_DATA_SIZE5_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal dout_4_port, dout_3_port, dout_2_port, dout_1_port, dout_0_port, n1, 
      n2, n3, n4, n5, net109193, net109194, net109195, net109196, net109197 : 
      std_logic;

begin
   dout <= ( dout_4_port, dout_3_port, dout_2_port, dout_1_port, dout_0_port );
   
   dout_reg_4_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           dout_4_port, QN => net109197);
   dout_reg_3_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           dout_3_port, QN => net109196);
   dout_reg_2_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           dout_2_port, QN => net109195);
   dout_reg_1_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           dout_1_port, QN => net109194);
   dout_reg_0_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           dout_0_port, QN => net109193);
   U2 : MUX2_X1 port map( A => dout_4_port, B => din(4), S => en, Z => n1);
   U3 : MUX2_X1 port map( A => dout_3_port, B => din(3), S => en, Z => n2);
   U4 : MUX2_X1 port map( A => dout_2_port, B => din(2), S => en, Z => n3);
   U5 : MUX2_X1 port map( A => dout_1_port, B => din(1), S => en, Z => n4);
   U6 : MUX2_X1 port map( A => dout_0_port, B => din(0), S => en, Z => n5);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_4 is

   port( reg_c, reg_f, reg_ff : in std_logic_vector (31 downto 0);  addr_c, 
         addr_f, addr_ff : in std_logic_vector (4 downto 0);  valid_f, valid_ff
         , dirty_f, dirty_ff, en : in std_logic;  output : out std_logic_vector
         (31 downto 0);  match_dirty_f, match_dirty_ff : out std_logic);

end FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_4;

architecture SYN_fwd_mux_2_arch of FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X4
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
      N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, 
      N106, N107, N108, N109, N110, N111, N112, n1, n2, n3, n4, n5, n6, n7, n8,
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55 : std_logic;

begin
   
   match_dirty_ff_reg : DLH_X1 port map( G => en, D => N111, Q => 
                           match_dirty_ff);
   output_reg_31_inst : DLH_X1 port map( G => en, D => N110, Q => output(31));
   output_reg_30_inst : DLH_X1 port map( G => en, D => N109, Q => output(30));
   output_reg_29_inst : DLH_X1 port map( G => en, D => N108, Q => output(29));
   output_reg_28_inst : DLH_X1 port map( G => en, D => N107, Q => output(28));
   output_reg_27_inst : DLH_X1 port map( G => en, D => N106, Q => output(27));
   output_reg_26_inst : DLH_X1 port map( G => en, D => N105, Q => output(26));
   output_reg_25_inst : DLH_X1 port map( G => en, D => N104, Q => output(25));
   output_reg_24_inst : DLH_X1 port map( G => en, D => N103, Q => output(24));
   output_reg_23_inst : DLH_X1 port map( G => en, D => N102, Q => output(23));
   output_reg_22_inst : DLH_X1 port map( G => en, D => N101, Q => output(22));
   output_reg_21_inst : DLH_X1 port map( G => en, D => N100, Q => output(21));
   output_reg_20_inst : DLH_X1 port map( G => en, D => N99, Q => output(20));
   output_reg_19_inst : DLH_X1 port map( G => en, D => N98, Q => output(19));
   output_reg_18_inst : DLH_X1 port map( G => en, D => N97, Q => output(18));
   output_reg_17_inst : DLH_X1 port map( G => en, D => N96, Q => output(17));
   output_reg_16_inst : DLH_X1 port map( G => en, D => N95, Q => output(16));
   output_reg_15_inst : DLH_X1 port map( G => en, D => N94, Q => output(15));
   output_reg_14_inst : DLH_X1 port map( G => en, D => N93, Q => output(14));
   output_reg_13_inst : DLH_X1 port map( G => en, D => N92, Q => output(13));
   output_reg_12_inst : DLH_X1 port map( G => en, D => N91, Q => output(12));
   output_reg_11_inst : DLH_X1 port map( G => en, D => N90, Q => output(11));
   output_reg_10_inst : DLH_X1 port map( G => en, D => N89, Q => output(10));
   output_reg_9_inst : DLH_X1 port map( G => en, D => N88, Q => output(9));
   output_reg_8_inst : DLH_X1 port map( G => en, D => N87, Q => output(8));
   output_reg_7_inst : DLH_X1 port map( G => en, D => N86, Q => output(7));
   output_reg_6_inst : DLH_X1 port map( G => en, D => N85, Q => output(6));
   output_reg_5_inst : DLH_X1 port map( G => en, D => N84, Q => output(5));
   output_reg_4_inst : DLH_X1 port map( G => en, D => N83, Q => output(4));
   output_reg_3_inst : DLH_X1 port map( G => en, D => N82, Q => output(3));
   output_reg_2_inst : DLH_X1 port map( G => en, D => N81, Q => output(2));
   output_reg_1_inst : DLH_X1 port map( G => en, D => N80, Q => output(1));
   output_reg_0_inst : DLH_X1 port map( G => en, D => N79, Q => output(0));
   match_dirty_f_reg : DLH_X1 port map( G => en, D => N112, Q => match_dirty_f)
                           ;
   U2 : OAI21_X4 port map( B1 => n38, B2 => n39, A => n36, ZN => n2);
   U3 : AND3_X2 port map( A1 => n36, A2 => n37, A3 => n38, ZN => n4);
   U4 : AND2_X2 port map( A1 => n39, A2 => n36, ZN => n3);
   U5 : INV_X1 port map( A => n1, ZN => N99);
   U6 : AOI222_X1 port map( A1 => reg_c(20), A2 => n2, B1 => reg_f(20), B2 => 
                           n3, C1 => reg_ff(20), C2 => n4, ZN => n1);
   U7 : INV_X1 port map( A => n5, ZN => N98);
   U8 : AOI222_X1 port map( A1 => reg_c(19), A2 => n2, B1 => reg_f(19), B2 => 
                           n3, C1 => reg_ff(19), C2 => n4, ZN => n5);
   U9 : INV_X1 port map( A => n6, ZN => N97);
   U10 : AOI222_X1 port map( A1 => reg_c(18), A2 => n2, B1 => reg_f(18), B2 => 
                           n3, C1 => reg_ff(18), C2 => n4, ZN => n6);
   U11 : INV_X1 port map( A => n7, ZN => N96);
   U12 : AOI222_X1 port map( A1 => reg_c(17), A2 => n2, B1 => reg_f(17), B2 => 
                           n3, C1 => reg_ff(17), C2 => n4, ZN => n7);
   U13 : INV_X1 port map( A => n8, ZN => N95);
   U14 : AOI222_X1 port map( A1 => reg_c(16), A2 => n2, B1 => reg_f(16), B2 => 
                           n3, C1 => reg_ff(16), C2 => n4, ZN => n8);
   U15 : INV_X1 port map( A => n9, ZN => N94);
   U16 : AOI222_X1 port map( A1 => reg_c(15), A2 => n2, B1 => reg_f(15), B2 => 
                           n3, C1 => reg_ff(15), C2 => n4, ZN => n9);
   U17 : INV_X1 port map( A => n10, ZN => N93);
   U18 : AOI222_X1 port map( A1 => reg_c(14), A2 => n2, B1 => reg_f(14), B2 => 
                           n3, C1 => reg_ff(14), C2 => n4, ZN => n10);
   U19 : INV_X1 port map( A => n11, ZN => N92);
   U20 : AOI222_X1 port map( A1 => reg_c(13), A2 => n2, B1 => reg_f(13), B2 => 
                           n3, C1 => reg_ff(13), C2 => n4, ZN => n11);
   U21 : INV_X1 port map( A => n12, ZN => N91);
   U22 : AOI222_X1 port map( A1 => reg_c(12), A2 => n2, B1 => reg_f(12), B2 => 
                           n3, C1 => reg_ff(12), C2 => n4, ZN => n12);
   U23 : INV_X1 port map( A => n13, ZN => N90);
   U24 : AOI222_X1 port map( A1 => reg_c(11), A2 => n2, B1 => reg_f(11), B2 => 
                           n3, C1 => reg_ff(11), C2 => n4, ZN => n13);
   U25 : INV_X1 port map( A => n14, ZN => N89);
   U26 : AOI222_X1 port map( A1 => reg_c(10), A2 => n2, B1 => reg_f(10), B2 => 
                           n3, C1 => reg_ff(10), C2 => n4, ZN => n14);
   U27 : INV_X1 port map( A => n15, ZN => N88);
   U28 : AOI222_X1 port map( A1 => reg_c(9), A2 => n2, B1 => reg_f(9), B2 => n3
                           , C1 => reg_ff(9), C2 => n4, ZN => n15);
   U29 : INV_X1 port map( A => n16, ZN => N87);
   U30 : AOI222_X1 port map( A1 => reg_c(8), A2 => n2, B1 => reg_f(8), B2 => n3
                           , C1 => reg_ff(8), C2 => n4, ZN => n16);
   U31 : INV_X1 port map( A => n17, ZN => N86);
   U32 : AOI222_X1 port map( A1 => reg_c(7), A2 => n2, B1 => reg_f(7), B2 => n3
                           , C1 => reg_ff(7), C2 => n4, ZN => n17);
   U33 : INV_X1 port map( A => n18, ZN => N85);
   U34 : AOI222_X1 port map( A1 => reg_c(6), A2 => n2, B1 => reg_f(6), B2 => n3
                           , C1 => reg_ff(6), C2 => n4, ZN => n18);
   U35 : INV_X1 port map( A => n19, ZN => N84);
   U36 : AOI222_X1 port map( A1 => reg_c(5), A2 => n2, B1 => reg_f(5), B2 => n3
                           , C1 => reg_ff(5), C2 => n4, ZN => n19);
   U37 : INV_X1 port map( A => n20, ZN => N83);
   U38 : AOI222_X1 port map( A1 => reg_c(4), A2 => n2, B1 => reg_f(4), B2 => n3
                           , C1 => reg_ff(4), C2 => n4, ZN => n20);
   U39 : INV_X1 port map( A => n21, ZN => N82);
   U40 : AOI222_X1 port map( A1 => reg_c(3), A2 => n2, B1 => reg_f(3), B2 => n3
                           , C1 => reg_ff(3), C2 => n4, ZN => n21);
   U41 : INV_X1 port map( A => n22, ZN => N81);
   U42 : AOI222_X1 port map( A1 => reg_c(2), A2 => n2, B1 => reg_f(2), B2 => n3
                           , C1 => reg_ff(2), C2 => n4, ZN => n22);
   U43 : INV_X1 port map( A => n23, ZN => N80);
   U44 : AOI222_X1 port map( A1 => reg_c(1), A2 => n2, B1 => reg_f(1), B2 => n3
                           , C1 => reg_ff(1), C2 => n4, ZN => n23);
   U45 : INV_X1 port map( A => n24, ZN => N79);
   U46 : AOI222_X1 port map( A1 => reg_c(0), A2 => n2, B1 => reg_f(0), B2 => n3
                           , C1 => reg_ff(0), C2 => n4, ZN => n24);
   U47 : AND2_X1 port map( A1 => dirty_f, A2 => n3, ZN => N112);
   U48 : AND2_X1 port map( A1 => dirty_ff, A2 => n4, ZN => N111);
   U49 : INV_X1 port map( A => n25, ZN => N110);
   U50 : AOI222_X1 port map( A1 => reg_c(31), A2 => n2, B1 => reg_f(31), B2 => 
                           n3, C1 => reg_ff(31), C2 => n4, ZN => n25);
   U51 : INV_X1 port map( A => n26, ZN => N109);
   U52 : AOI222_X1 port map( A1 => reg_c(30), A2 => n2, B1 => reg_f(30), B2 => 
                           n3, C1 => reg_ff(30), C2 => n4, ZN => n26);
   U53 : INV_X1 port map( A => n27, ZN => N108);
   U54 : AOI222_X1 port map( A1 => reg_c(29), A2 => n2, B1 => reg_f(29), B2 => 
                           n3, C1 => reg_ff(29), C2 => n4, ZN => n27);
   U55 : INV_X1 port map( A => n28, ZN => N107);
   U56 : AOI222_X1 port map( A1 => reg_c(28), A2 => n2, B1 => reg_f(28), B2 => 
                           n3, C1 => reg_ff(28), C2 => n4, ZN => n28);
   U57 : INV_X1 port map( A => n29, ZN => N106);
   U58 : AOI222_X1 port map( A1 => reg_c(27), A2 => n2, B1 => reg_f(27), B2 => 
                           n3, C1 => reg_ff(27), C2 => n4, ZN => n29);
   U59 : INV_X1 port map( A => n30, ZN => N105);
   U60 : AOI222_X1 port map( A1 => reg_c(26), A2 => n2, B1 => reg_f(26), B2 => 
                           n3, C1 => reg_ff(26), C2 => n4, ZN => n30);
   U61 : INV_X1 port map( A => n31, ZN => N104);
   U62 : AOI222_X1 port map( A1 => reg_c(25), A2 => n2, B1 => reg_f(25), B2 => 
                           n3, C1 => reg_ff(25), C2 => n4, ZN => n31);
   U63 : INV_X1 port map( A => n32, ZN => N103);
   U64 : AOI222_X1 port map( A1 => reg_c(24), A2 => n2, B1 => reg_f(24), B2 => 
                           n3, C1 => reg_ff(24), C2 => n4, ZN => n32);
   U65 : INV_X1 port map( A => n33, ZN => N102);
   U66 : AOI222_X1 port map( A1 => reg_c(23), A2 => n2, B1 => reg_f(23), B2 => 
                           n3, C1 => reg_ff(23), C2 => n4, ZN => n33);
   U67 : INV_X1 port map( A => n34, ZN => N101);
   U68 : AOI222_X1 port map( A1 => reg_c(22), A2 => n2, B1 => reg_f(22), B2 => 
                           n3, C1 => reg_ff(22), C2 => n4, ZN => n34);
   U69 : INV_X1 port map( A => n35, ZN => N100);
   U70 : AOI222_X1 port map( A1 => reg_c(21), A2 => n2, B1 => reg_f(21), B2 => 
                           n3, C1 => reg_ff(21), C2 => n4, ZN => n35);
   U71 : NAND4_X1 port map( A1 => n40, A2 => n41, A3 => n42, A4 => n43, ZN => 
                           n36);
   U72 : NOR2_X1 port map( A1 => addr_c(1), A2 => addr_c(0), ZN => n43);
   U73 : INV_X1 port map( A => addr_c(4), ZN => n41);
   U74 : INV_X1 port map( A => n37, ZN => n39);
   U75 : NAND4_X1 port map( A1 => n44, A2 => valid_f, A3 => n45, A4 => n46, ZN 
                           => n37);
   U76 : NOR3_X1 port map( A1 => n47, A2 => n48, A3 => n49, ZN => n46);
   U77 : XOR2_X1 port map( A => addr_f(2), B => addr_c(2), Z => n49);
   U78 : XOR2_X1 port map( A => addr_f(4), B => addr_c(4), Z => n48);
   U79 : XOR2_X1 port map( A => addr_f(3), B => addr_c(3), Z => n47);
   U80 : XNOR2_X1 port map( A => addr_c(0), B => addr_f(0), ZN => n45);
   U81 : XNOR2_X1 port map( A => addr_c(1), B => addr_f(1), ZN => n44);
   U82 : AND4_X1 port map( A1 => n50, A2 => valid_ff, A3 => n51, A4 => n52, ZN 
                           => n38);
   U83 : NOR3_X1 port map( A1 => n53, A2 => n54, A3 => n55, ZN => n52);
   U84 : XOR2_X1 port map( A => addr_ff(0), B => addr_c(0), Z => n55);
   U85 : XOR2_X1 port map( A => addr_ff(1), B => addr_c(1), Z => n54);
   U86 : XOR2_X1 port map( A => addr_ff(4), B => addr_c(4), Z => n53);
   U87 : XOR2_X1 port map( A => n40, B => addr_ff(3), Z => n51);
   U88 : INV_X1 port map( A => addr_c(3), ZN => n40);
   U89 : XOR2_X1 port map( A => n42, B => addr_ff(2), Z => n50);
   U90 : INV_X1 port map( A => addr_c(2), ZN => n42);

end SYN_fwd_mux_2_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_3 is

   port( reg_c, reg_f, reg_ff : in std_logic_vector (31 downto 0);  addr_c, 
         addr_f, addr_ff : in std_logic_vector (4 downto 0);  valid_f, valid_ff
         , dirty_f, dirty_ff, en : in std_logic;  output : out std_logic_vector
         (31 downto 0);  match_dirty_f, match_dirty_ff : out std_logic);

end FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_3;

architecture SYN_fwd_mux_2_arch of FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X4
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X2
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
      N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, 
      N106, N107, N108, N109, N110, N111, N112, n1, n2, n3, n4, n5, n6, n7, n8,
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55 : std_logic;

begin
   
   match_dirty_ff_reg : DLH_X1 port map( G => en, D => N111, Q => 
                           match_dirty_ff);
   output_reg_31_inst : DLH_X1 port map( G => en, D => N110, Q => output(31));
   output_reg_30_inst : DLH_X1 port map( G => en, D => N109, Q => output(30));
   output_reg_29_inst : DLH_X1 port map( G => en, D => N108, Q => output(29));
   output_reg_28_inst : DLH_X1 port map( G => en, D => N107, Q => output(28));
   output_reg_27_inst : DLH_X1 port map( G => en, D => N106, Q => output(27));
   output_reg_26_inst : DLH_X1 port map( G => en, D => N105, Q => output(26));
   output_reg_25_inst : DLH_X1 port map( G => en, D => N104, Q => output(25));
   output_reg_24_inst : DLH_X1 port map( G => en, D => N103, Q => output(24));
   output_reg_23_inst : DLH_X1 port map( G => en, D => N102, Q => output(23));
   output_reg_22_inst : DLH_X1 port map( G => en, D => N101, Q => output(22));
   output_reg_21_inst : DLH_X1 port map( G => en, D => N100, Q => output(21));
   output_reg_20_inst : DLH_X1 port map( G => en, D => N99, Q => output(20));
   output_reg_19_inst : DLH_X1 port map( G => en, D => N98, Q => output(19));
   output_reg_18_inst : DLH_X1 port map( G => en, D => N97, Q => output(18));
   output_reg_17_inst : DLH_X1 port map( G => en, D => N96, Q => output(17));
   output_reg_16_inst : DLH_X1 port map( G => en, D => N95, Q => output(16));
   match_dirty_f_reg : DLH_X1 port map( G => en, D => N112, Q => match_dirty_f)
                           ;
   output_reg_12_inst : DLH_X2 port map( G => en, D => N91, Q => output(12));
   output_reg_4_inst : DLH_X2 port map( G => en, D => N83, Q => output(4));
   output_reg_6_inst : DLH_X2 port map( G => en, D => N85, Q => output(6));
   output_reg_11_inst : DLH_X2 port map( G => en, D => N90, Q => output(11));
   output_reg_15_inst : DLH_X2 port map( G => en, D => N94, Q => output(15));
   output_reg_7_inst : DLH_X2 port map( G => en, D => N86, Q => output(7));
   output_reg_13_inst : DLH_X2 port map( G => en, D => N92, Q => output(13));
   output_reg_3_inst : DLH_X2 port map( G => en, D => N82, Q => output(3));
   output_reg_14_inst : DLH_X2 port map( G => en, D => N93, Q => output(14));
   output_reg_10_inst : DLH_X2 port map( G => en, D => N89, Q => output(10));
   output_reg_8_inst : DLH_X2 port map( G => en, D => N87, Q => output(8));
   output_reg_5_inst : DLH_X2 port map( G => en, D => N84, Q => output(5));
   output_reg_2_inst : DLH_X2 port map( G => en, D => N81, Q => output(2));
   output_reg_0_inst : DLH_X2 port map( G => en, D => N79, Q => output(0));
   output_reg_1_inst : DLH_X2 port map( G => en, D => N80, Q => output(1));
   output_reg_9_inst : DLH_X2 port map( G => en, D => N88, Q => output(9));
   U2 : OAI21_X4 port map( B1 => n38, B2 => n39, A => n36, ZN => n2);
   U3 : AND3_X2 port map( A1 => n36, A2 => n37, A3 => n38, ZN => n4);
   U4 : AND2_X2 port map( A1 => n39, A2 => n36, ZN => n3);
   U5 : INV_X1 port map( A => n1, ZN => N99);
   U6 : AOI222_X1 port map( A1 => reg_c(20), A2 => n2, B1 => reg_f(20), B2 => 
                           n3, C1 => reg_ff(20), C2 => n4, ZN => n1);
   U7 : INV_X1 port map( A => n5, ZN => N98);
   U8 : AOI222_X1 port map( A1 => reg_c(19), A2 => n2, B1 => reg_f(19), B2 => 
                           n3, C1 => reg_ff(19), C2 => n4, ZN => n5);
   U9 : INV_X1 port map( A => n6, ZN => N97);
   U10 : AOI222_X1 port map( A1 => reg_c(18), A2 => n2, B1 => reg_f(18), B2 => 
                           n3, C1 => reg_ff(18), C2 => n4, ZN => n6);
   U11 : INV_X1 port map( A => n7, ZN => N96);
   U12 : AOI222_X1 port map( A1 => reg_c(17), A2 => n2, B1 => reg_f(17), B2 => 
                           n3, C1 => reg_ff(17), C2 => n4, ZN => n7);
   U13 : INV_X1 port map( A => n8, ZN => N95);
   U14 : AOI222_X1 port map( A1 => reg_c(16), A2 => n2, B1 => reg_f(16), B2 => 
                           n3, C1 => reg_ff(16), C2 => n4, ZN => n8);
   U15 : INV_X1 port map( A => n9, ZN => N94);
   U16 : AOI222_X1 port map( A1 => reg_c(15), A2 => n2, B1 => reg_f(15), B2 => 
                           n3, C1 => reg_ff(15), C2 => n4, ZN => n9);
   U17 : INV_X1 port map( A => n10, ZN => N93);
   U18 : AOI222_X1 port map( A1 => reg_c(14), A2 => n2, B1 => reg_f(14), B2 => 
                           n3, C1 => reg_ff(14), C2 => n4, ZN => n10);
   U19 : INV_X1 port map( A => n11, ZN => N92);
   U20 : AOI222_X1 port map( A1 => reg_c(13), A2 => n2, B1 => reg_f(13), B2 => 
                           n3, C1 => reg_ff(13), C2 => n4, ZN => n11);
   U21 : INV_X1 port map( A => n12, ZN => N91);
   U22 : AOI222_X1 port map( A1 => reg_c(12), A2 => n2, B1 => reg_f(12), B2 => 
                           n3, C1 => reg_ff(12), C2 => n4, ZN => n12);
   U23 : INV_X1 port map( A => n13, ZN => N90);
   U24 : AOI222_X1 port map( A1 => reg_c(11), A2 => n2, B1 => reg_f(11), B2 => 
                           n3, C1 => reg_ff(11), C2 => n4, ZN => n13);
   U25 : INV_X1 port map( A => n14, ZN => N89);
   U26 : AOI222_X1 port map( A1 => reg_c(10), A2 => n2, B1 => reg_f(10), B2 => 
                           n3, C1 => reg_ff(10), C2 => n4, ZN => n14);
   U27 : INV_X1 port map( A => n15, ZN => N88);
   U28 : AOI222_X1 port map( A1 => reg_c(9), A2 => n2, B1 => reg_f(9), B2 => n3
                           , C1 => reg_ff(9), C2 => n4, ZN => n15);
   U29 : INV_X1 port map( A => n16, ZN => N87);
   U30 : AOI222_X1 port map( A1 => reg_c(8), A2 => n2, B1 => reg_f(8), B2 => n3
                           , C1 => reg_ff(8), C2 => n4, ZN => n16);
   U31 : INV_X1 port map( A => n17, ZN => N86);
   U32 : AOI222_X1 port map( A1 => reg_c(7), A2 => n2, B1 => reg_f(7), B2 => n3
                           , C1 => reg_ff(7), C2 => n4, ZN => n17);
   U33 : INV_X1 port map( A => n18, ZN => N85);
   U34 : AOI222_X1 port map( A1 => reg_c(6), A2 => n2, B1 => reg_f(6), B2 => n3
                           , C1 => reg_ff(6), C2 => n4, ZN => n18);
   U35 : INV_X1 port map( A => n19, ZN => N84);
   U36 : AOI222_X1 port map( A1 => reg_c(5), A2 => n2, B1 => reg_f(5), B2 => n3
                           , C1 => reg_ff(5), C2 => n4, ZN => n19);
   U37 : INV_X1 port map( A => n20, ZN => N83);
   U38 : AOI222_X1 port map( A1 => reg_c(4), A2 => n2, B1 => reg_f(4), B2 => n3
                           , C1 => reg_ff(4), C2 => n4, ZN => n20);
   U39 : INV_X1 port map( A => n21, ZN => N82);
   U40 : AOI222_X1 port map( A1 => reg_c(3), A2 => n2, B1 => reg_f(3), B2 => n3
                           , C1 => reg_ff(3), C2 => n4, ZN => n21);
   U41 : INV_X1 port map( A => n22, ZN => N81);
   U42 : AOI222_X1 port map( A1 => reg_c(2), A2 => n2, B1 => reg_f(2), B2 => n3
                           , C1 => reg_ff(2), C2 => n4, ZN => n22);
   U43 : INV_X1 port map( A => n23, ZN => N80);
   U44 : AOI222_X1 port map( A1 => reg_c(1), A2 => n2, B1 => reg_f(1), B2 => n3
                           , C1 => reg_ff(1), C2 => n4, ZN => n23);
   U45 : INV_X1 port map( A => n24, ZN => N79);
   U46 : AOI222_X1 port map( A1 => reg_c(0), A2 => n2, B1 => reg_f(0), B2 => n3
                           , C1 => reg_ff(0), C2 => n4, ZN => n24);
   U47 : AND2_X1 port map( A1 => dirty_f, A2 => n3, ZN => N112);
   U48 : AND2_X1 port map( A1 => dirty_ff, A2 => n4, ZN => N111);
   U49 : INV_X1 port map( A => n25, ZN => N110);
   U50 : AOI222_X1 port map( A1 => reg_c(31), A2 => n2, B1 => reg_f(31), B2 => 
                           n3, C1 => reg_ff(31), C2 => n4, ZN => n25);
   U51 : INV_X1 port map( A => n26, ZN => N109);
   U52 : AOI222_X1 port map( A1 => reg_c(30), A2 => n2, B1 => reg_f(30), B2 => 
                           n3, C1 => reg_ff(30), C2 => n4, ZN => n26);
   U53 : INV_X1 port map( A => n27, ZN => N108);
   U54 : AOI222_X1 port map( A1 => reg_c(29), A2 => n2, B1 => reg_f(29), B2 => 
                           n3, C1 => reg_ff(29), C2 => n4, ZN => n27);
   U55 : INV_X1 port map( A => n28, ZN => N107);
   U56 : AOI222_X1 port map( A1 => reg_c(28), A2 => n2, B1 => reg_f(28), B2 => 
                           n3, C1 => reg_ff(28), C2 => n4, ZN => n28);
   U57 : INV_X1 port map( A => n29, ZN => N106);
   U58 : AOI222_X1 port map( A1 => reg_c(27), A2 => n2, B1 => reg_f(27), B2 => 
                           n3, C1 => reg_ff(27), C2 => n4, ZN => n29);
   U59 : INV_X1 port map( A => n30, ZN => N105);
   U60 : AOI222_X1 port map( A1 => reg_c(26), A2 => n2, B1 => reg_f(26), B2 => 
                           n3, C1 => reg_ff(26), C2 => n4, ZN => n30);
   U61 : INV_X1 port map( A => n31, ZN => N104);
   U62 : AOI222_X1 port map( A1 => reg_c(25), A2 => n2, B1 => reg_f(25), B2 => 
                           n3, C1 => reg_ff(25), C2 => n4, ZN => n31);
   U63 : INV_X1 port map( A => n32, ZN => N103);
   U64 : AOI222_X1 port map( A1 => reg_c(24), A2 => n2, B1 => reg_f(24), B2 => 
                           n3, C1 => reg_ff(24), C2 => n4, ZN => n32);
   U65 : INV_X1 port map( A => n33, ZN => N102);
   U66 : AOI222_X1 port map( A1 => reg_c(23), A2 => n2, B1 => reg_f(23), B2 => 
                           n3, C1 => reg_ff(23), C2 => n4, ZN => n33);
   U67 : INV_X1 port map( A => n34, ZN => N101);
   U68 : AOI222_X1 port map( A1 => reg_c(22), A2 => n2, B1 => reg_f(22), B2 => 
                           n3, C1 => reg_ff(22), C2 => n4, ZN => n34);
   U69 : INV_X1 port map( A => n35, ZN => N100);
   U70 : AOI222_X1 port map( A1 => reg_c(21), A2 => n2, B1 => reg_f(21), B2 => 
                           n3, C1 => reg_ff(21), C2 => n4, ZN => n35);
   U71 : NAND4_X1 port map( A1 => n40, A2 => n41, A3 => n42, A4 => n43, ZN => 
                           n36);
   U72 : NOR2_X1 port map( A1 => addr_c(1), A2 => addr_c(0), ZN => n43);
   U73 : INV_X1 port map( A => addr_c(4), ZN => n41);
   U74 : INV_X1 port map( A => n37, ZN => n39);
   U75 : NAND4_X1 port map( A1 => n44, A2 => valid_f, A3 => n45, A4 => n46, ZN 
                           => n37);
   U76 : NOR3_X1 port map( A1 => n47, A2 => n48, A3 => n49, ZN => n46);
   U77 : XOR2_X1 port map( A => addr_f(2), B => addr_c(2), Z => n49);
   U78 : XOR2_X1 port map( A => addr_f(4), B => addr_c(4), Z => n48);
   U79 : XOR2_X1 port map( A => addr_f(3), B => addr_c(3), Z => n47);
   U80 : XNOR2_X1 port map( A => addr_c(0), B => addr_f(0), ZN => n45);
   U81 : XNOR2_X1 port map( A => addr_c(1), B => addr_f(1), ZN => n44);
   U82 : AND4_X1 port map( A1 => n50, A2 => valid_ff, A3 => n51, A4 => n52, ZN 
                           => n38);
   U83 : NOR3_X1 port map( A1 => n53, A2 => n54, A3 => n55, ZN => n52);
   U84 : XOR2_X1 port map( A => addr_ff(0), B => addr_c(0), Z => n55);
   U85 : XOR2_X1 port map( A => addr_ff(1), B => addr_c(1), Z => n54);
   U86 : XOR2_X1 port map( A => addr_ff(4), B => addr_c(4), Z => n53);
   U87 : XOR2_X1 port map( A => n40, B => addr_ff(3), Z => n51);
   U88 : INV_X1 port map( A => addr_c(3), ZN => n40);
   U89 : XOR2_X1 port map( A => n42, B => addr_ff(2), Z => n50);
   U90 : INV_X1 port map( A => addr_c(2), ZN => n42);

end SYN_fwd_mux_2_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_2 is

   port( reg_c, reg_f, reg_ff : in std_logic_vector (31 downto 0);  addr_c, 
         addr_f, addr_ff : in std_logic_vector (4 downto 0);  valid_f, valid_ff
         , dirty_f, dirty_ff, en : in std_logic;  output : out std_logic_vector
         (31 downto 0);  match_dirty_f, match_dirty_ff : out std_logic);

end FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_2;

architecture SYN_fwd_mux_2_arch of FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X4
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
      N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, 
      N106, N107, N108, N109, N110, N111, N112, n1, n2, n3, n4, n5, n6, n7, n8,
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55 : std_logic;

begin
   
   match_dirty_ff_reg : DLH_X1 port map( G => en, D => N111, Q => 
                           match_dirty_ff);
   output_reg_31_inst : DLH_X1 port map( G => en, D => N110, Q => output(31));
   output_reg_30_inst : DLH_X1 port map( G => en, D => N109, Q => output(30));
   output_reg_29_inst : DLH_X1 port map( G => en, D => N108, Q => output(29));
   output_reg_28_inst : DLH_X1 port map( G => en, D => N107, Q => output(28));
   output_reg_27_inst : DLH_X1 port map( G => en, D => N106, Q => output(27));
   output_reg_26_inst : DLH_X1 port map( G => en, D => N105, Q => output(26));
   output_reg_25_inst : DLH_X1 port map( G => en, D => N104, Q => output(25));
   output_reg_24_inst : DLH_X1 port map( G => en, D => N103, Q => output(24));
   output_reg_23_inst : DLH_X1 port map( G => en, D => N102, Q => output(23));
   output_reg_22_inst : DLH_X1 port map( G => en, D => N101, Q => output(22));
   output_reg_21_inst : DLH_X1 port map( G => en, D => N100, Q => output(21));
   output_reg_20_inst : DLH_X1 port map( G => en, D => N99, Q => output(20));
   output_reg_19_inst : DLH_X1 port map( G => en, D => N98, Q => output(19));
   output_reg_18_inst : DLH_X1 port map( G => en, D => N97, Q => output(18));
   output_reg_17_inst : DLH_X1 port map( G => en, D => N96, Q => output(17));
   output_reg_16_inst : DLH_X1 port map( G => en, D => N95, Q => output(16));
   output_reg_15_inst : DLH_X1 port map( G => en, D => N94, Q => output(15));
   output_reg_14_inst : DLH_X1 port map( G => en, D => N93, Q => output(14));
   output_reg_13_inst : DLH_X1 port map( G => en, D => N92, Q => output(13));
   output_reg_12_inst : DLH_X1 port map( G => en, D => N91, Q => output(12));
   output_reg_11_inst : DLH_X1 port map( G => en, D => N90, Q => output(11));
   output_reg_10_inst : DLH_X1 port map( G => en, D => N89, Q => output(10));
   output_reg_9_inst : DLH_X1 port map( G => en, D => N88, Q => output(9));
   output_reg_8_inst : DLH_X1 port map( G => en, D => N87, Q => output(8));
   output_reg_7_inst : DLH_X1 port map( G => en, D => N86, Q => output(7));
   output_reg_6_inst : DLH_X1 port map( G => en, D => N85, Q => output(6));
   output_reg_5_inst : DLH_X1 port map( G => en, D => N84, Q => output(5));
   output_reg_4_inst : DLH_X1 port map( G => en, D => N83, Q => output(4));
   output_reg_3_inst : DLH_X1 port map( G => en, D => N82, Q => output(3));
   output_reg_2_inst : DLH_X1 port map( G => en, D => N81, Q => output(2));
   output_reg_1_inst : DLH_X1 port map( G => en, D => N80, Q => output(1));
   output_reg_0_inst : DLH_X1 port map( G => en, D => N79, Q => output(0));
   match_dirty_f_reg : DLH_X1 port map( G => en, D => N112, Q => match_dirty_f)
                           ;
   U2 : OAI21_X4 port map( B1 => n38, B2 => n39, A => n36, ZN => n2);
   U3 : AND3_X2 port map( A1 => n36, A2 => n37, A3 => n38, ZN => n4);
   U4 : AND2_X2 port map( A1 => n39, A2 => n36, ZN => n3);
   U5 : INV_X1 port map( A => n1, ZN => N99);
   U6 : AOI222_X1 port map( A1 => reg_c(20), A2 => n2, B1 => reg_f(20), B2 => 
                           n3, C1 => reg_ff(20), C2 => n4, ZN => n1);
   U7 : INV_X1 port map( A => n5, ZN => N98);
   U8 : AOI222_X1 port map( A1 => reg_c(19), A2 => n2, B1 => reg_f(19), B2 => 
                           n3, C1 => reg_ff(19), C2 => n4, ZN => n5);
   U9 : INV_X1 port map( A => n6, ZN => N97);
   U10 : AOI222_X1 port map( A1 => reg_c(18), A2 => n2, B1 => reg_f(18), B2 => 
                           n3, C1 => reg_ff(18), C2 => n4, ZN => n6);
   U11 : INV_X1 port map( A => n7, ZN => N96);
   U12 : AOI222_X1 port map( A1 => reg_c(17), A2 => n2, B1 => reg_f(17), B2 => 
                           n3, C1 => reg_ff(17), C2 => n4, ZN => n7);
   U13 : INV_X1 port map( A => n8, ZN => N95);
   U14 : AOI222_X1 port map( A1 => reg_c(16), A2 => n2, B1 => reg_f(16), B2 => 
                           n3, C1 => reg_ff(16), C2 => n4, ZN => n8);
   U15 : INV_X1 port map( A => n9, ZN => N94);
   U16 : AOI222_X1 port map( A1 => reg_c(15), A2 => n2, B1 => reg_f(15), B2 => 
                           n3, C1 => reg_ff(15), C2 => n4, ZN => n9);
   U17 : INV_X1 port map( A => n10, ZN => N93);
   U18 : AOI222_X1 port map( A1 => reg_c(14), A2 => n2, B1 => reg_f(14), B2 => 
                           n3, C1 => reg_ff(14), C2 => n4, ZN => n10);
   U19 : INV_X1 port map( A => n11, ZN => N92);
   U20 : AOI222_X1 port map( A1 => reg_c(13), A2 => n2, B1 => reg_f(13), B2 => 
                           n3, C1 => reg_ff(13), C2 => n4, ZN => n11);
   U21 : INV_X1 port map( A => n12, ZN => N91);
   U22 : AOI222_X1 port map( A1 => reg_c(12), A2 => n2, B1 => reg_f(12), B2 => 
                           n3, C1 => reg_ff(12), C2 => n4, ZN => n12);
   U23 : INV_X1 port map( A => n13, ZN => N90);
   U24 : AOI222_X1 port map( A1 => reg_c(11), A2 => n2, B1 => reg_f(11), B2 => 
                           n3, C1 => reg_ff(11), C2 => n4, ZN => n13);
   U25 : INV_X1 port map( A => n14, ZN => N89);
   U26 : AOI222_X1 port map( A1 => reg_c(10), A2 => n2, B1 => reg_f(10), B2 => 
                           n3, C1 => reg_ff(10), C2 => n4, ZN => n14);
   U27 : INV_X1 port map( A => n15, ZN => N88);
   U28 : AOI222_X1 port map( A1 => reg_c(9), A2 => n2, B1 => reg_f(9), B2 => n3
                           , C1 => reg_ff(9), C2 => n4, ZN => n15);
   U29 : INV_X1 port map( A => n16, ZN => N87);
   U30 : AOI222_X1 port map( A1 => reg_c(8), A2 => n2, B1 => reg_f(8), B2 => n3
                           , C1 => reg_ff(8), C2 => n4, ZN => n16);
   U31 : INV_X1 port map( A => n17, ZN => N86);
   U32 : AOI222_X1 port map( A1 => reg_c(7), A2 => n2, B1 => reg_f(7), B2 => n3
                           , C1 => reg_ff(7), C2 => n4, ZN => n17);
   U33 : INV_X1 port map( A => n18, ZN => N85);
   U34 : AOI222_X1 port map( A1 => reg_c(6), A2 => n2, B1 => reg_f(6), B2 => n3
                           , C1 => reg_ff(6), C2 => n4, ZN => n18);
   U35 : INV_X1 port map( A => n19, ZN => N84);
   U36 : AOI222_X1 port map( A1 => reg_c(5), A2 => n2, B1 => reg_f(5), B2 => n3
                           , C1 => reg_ff(5), C2 => n4, ZN => n19);
   U37 : INV_X1 port map( A => n20, ZN => N83);
   U38 : AOI222_X1 port map( A1 => reg_c(4), A2 => n2, B1 => reg_f(4), B2 => n3
                           , C1 => reg_ff(4), C2 => n4, ZN => n20);
   U39 : INV_X1 port map( A => n21, ZN => N82);
   U40 : AOI222_X1 port map( A1 => reg_c(3), A2 => n2, B1 => reg_f(3), B2 => n3
                           , C1 => reg_ff(3), C2 => n4, ZN => n21);
   U41 : INV_X1 port map( A => n22, ZN => N81);
   U42 : AOI222_X1 port map( A1 => reg_c(2), A2 => n2, B1 => reg_f(2), B2 => n3
                           , C1 => reg_ff(2), C2 => n4, ZN => n22);
   U43 : INV_X1 port map( A => n23, ZN => N80);
   U44 : AOI222_X1 port map( A1 => reg_c(1), A2 => n2, B1 => reg_f(1), B2 => n3
                           , C1 => reg_ff(1), C2 => n4, ZN => n23);
   U45 : INV_X1 port map( A => n24, ZN => N79);
   U46 : AOI222_X1 port map( A1 => reg_c(0), A2 => n2, B1 => reg_f(0), B2 => n3
                           , C1 => reg_ff(0), C2 => n4, ZN => n24);
   U47 : AND2_X1 port map( A1 => dirty_f, A2 => n3, ZN => N112);
   U48 : AND2_X1 port map( A1 => dirty_ff, A2 => n4, ZN => N111);
   U49 : INV_X1 port map( A => n25, ZN => N110);
   U50 : AOI222_X1 port map( A1 => reg_c(31), A2 => n2, B1 => reg_f(31), B2 => 
                           n3, C1 => reg_ff(31), C2 => n4, ZN => n25);
   U51 : INV_X1 port map( A => n26, ZN => N109);
   U52 : AOI222_X1 port map( A1 => reg_c(30), A2 => n2, B1 => reg_f(30), B2 => 
                           n3, C1 => reg_ff(30), C2 => n4, ZN => n26);
   U53 : INV_X1 port map( A => n27, ZN => N108);
   U54 : AOI222_X1 port map( A1 => reg_c(29), A2 => n2, B1 => reg_f(29), B2 => 
                           n3, C1 => reg_ff(29), C2 => n4, ZN => n27);
   U55 : INV_X1 port map( A => n28, ZN => N107);
   U56 : AOI222_X1 port map( A1 => reg_c(28), A2 => n2, B1 => reg_f(28), B2 => 
                           n3, C1 => reg_ff(28), C2 => n4, ZN => n28);
   U57 : INV_X1 port map( A => n29, ZN => N106);
   U58 : AOI222_X1 port map( A1 => reg_c(27), A2 => n2, B1 => reg_f(27), B2 => 
                           n3, C1 => reg_ff(27), C2 => n4, ZN => n29);
   U59 : INV_X1 port map( A => n30, ZN => N105);
   U60 : AOI222_X1 port map( A1 => reg_c(26), A2 => n2, B1 => reg_f(26), B2 => 
                           n3, C1 => reg_ff(26), C2 => n4, ZN => n30);
   U61 : INV_X1 port map( A => n31, ZN => N104);
   U62 : AOI222_X1 port map( A1 => reg_c(25), A2 => n2, B1 => reg_f(25), B2 => 
                           n3, C1 => reg_ff(25), C2 => n4, ZN => n31);
   U63 : INV_X1 port map( A => n32, ZN => N103);
   U64 : AOI222_X1 port map( A1 => reg_c(24), A2 => n2, B1 => reg_f(24), B2 => 
                           n3, C1 => reg_ff(24), C2 => n4, ZN => n32);
   U65 : INV_X1 port map( A => n33, ZN => N102);
   U66 : AOI222_X1 port map( A1 => reg_c(23), A2 => n2, B1 => reg_f(23), B2 => 
                           n3, C1 => reg_ff(23), C2 => n4, ZN => n33);
   U67 : INV_X1 port map( A => n34, ZN => N101);
   U68 : AOI222_X1 port map( A1 => reg_c(22), A2 => n2, B1 => reg_f(22), B2 => 
                           n3, C1 => reg_ff(22), C2 => n4, ZN => n34);
   U69 : INV_X1 port map( A => n35, ZN => N100);
   U70 : AOI222_X1 port map( A1 => reg_c(21), A2 => n2, B1 => reg_f(21), B2 => 
                           n3, C1 => reg_ff(21), C2 => n4, ZN => n35);
   U71 : NAND4_X1 port map( A1 => n40, A2 => n41, A3 => n42, A4 => n43, ZN => 
                           n36);
   U72 : NOR2_X1 port map( A1 => addr_c(1), A2 => addr_c(0), ZN => n43);
   U73 : INV_X1 port map( A => addr_c(4), ZN => n41);
   U74 : INV_X1 port map( A => n37, ZN => n39);
   U75 : NAND4_X1 port map( A1 => n44, A2 => valid_f, A3 => n45, A4 => n46, ZN 
                           => n37);
   U76 : NOR3_X1 port map( A1 => n47, A2 => n48, A3 => n49, ZN => n46);
   U77 : XOR2_X1 port map( A => addr_f(2), B => addr_c(2), Z => n49);
   U78 : XOR2_X1 port map( A => addr_f(4), B => addr_c(4), Z => n48);
   U79 : XOR2_X1 port map( A => addr_f(3), B => addr_c(3), Z => n47);
   U80 : XNOR2_X1 port map( A => addr_c(0), B => addr_f(0), ZN => n45);
   U81 : XNOR2_X1 port map( A => addr_c(1), B => addr_f(1), ZN => n44);
   U82 : AND4_X1 port map( A1 => n50, A2 => valid_ff, A3 => n51, A4 => n52, ZN 
                           => n38);
   U83 : NOR3_X1 port map( A1 => n53, A2 => n54, A3 => n55, ZN => n52);
   U84 : XOR2_X1 port map( A => addr_ff(0), B => addr_c(0), Z => n55);
   U85 : XOR2_X1 port map( A => addr_ff(1), B => addr_c(1), Z => n54);
   U86 : XOR2_X1 port map( A => addr_ff(4), B => addr_c(4), Z => n53);
   U87 : XOR2_X1 port map( A => n40, B => addr_ff(3), Z => n51);
   U88 : INV_X1 port map( A => addr_c(3), ZN => n40);
   U89 : XOR2_X1 port map( A => n42, B => addr_ff(2), Z => n50);
   U90 : INV_X1 port map( A => addr_c(2), ZN => n42);

end SYN_fwd_mux_2_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_1 is

   port( reg_c, reg_f, reg_ff : in std_logic_vector (31 downto 0);  addr_c, 
         addr_f, addr_ff : in std_logic_vector (4 downto 0);  valid_f, valid_ff
         , dirty_f, dirty_ff, en : in std_logic;  output : out std_logic_vector
         (31 downto 0);  match_dirty_f, match_dirty_ff : out std_logic);

end FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_1;

architecture SYN_fwd_mux_2_arch of FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X4
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
      N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, 
      N106, N107, N108, N109, N110, N111, N112, n1, n2, n3, n4, n5, n6, n7, n8,
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55 : std_logic;

begin
   
   match_dirty_ff_reg : DLH_X1 port map( G => en, D => N111, Q => 
                           match_dirty_ff);
   output_reg_31_inst : DLH_X1 port map( G => en, D => N110, Q => output(31));
   output_reg_30_inst : DLH_X1 port map( G => en, D => N109, Q => output(30));
   output_reg_29_inst : DLH_X1 port map( G => en, D => N108, Q => output(29));
   output_reg_28_inst : DLH_X1 port map( G => en, D => N107, Q => output(28));
   output_reg_27_inst : DLH_X1 port map( G => en, D => N106, Q => output(27));
   output_reg_26_inst : DLH_X1 port map( G => en, D => N105, Q => output(26));
   output_reg_25_inst : DLH_X1 port map( G => en, D => N104, Q => output(25));
   output_reg_24_inst : DLH_X1 port map( G => en, D => N103, Q => output(24));
   output_reg_23_inst : DLH_X1 port map( G => en, D => N102, Q => output(23));
   output_reg_22_inst : DLH_X1 port map( G => en, D => N101, Q => output(22));
   output_reg_21_inst : DLH_X1 port map( G => en, D => N100, Q => output(21));
   output_reg_20_inst : DLH_X1 port map( G => en, D => N99, Q => output(20));
   output_reg_19_inst : DLH_X1 port map( G => en, D => N98, Q => output(19));
   output_reg_18_inst : DLH_X1 port map( G => en, D => N97, Q => output(18));
   output_reg_17_inst : DLH_X1 port map( G => en, D => N96, Q => output(17));
   output_reg_16_inst : DLH_X1 port map( G => en, D => N95, Q => output(16));
   output_reg_15_inst : DLH_X1 port map( G => en, D => N94, Q => output(15));
   output_reg_14_inst : DLH_X1 port map( G => en, D => N93, Q => output(14));
   output_reg_13_inst : DLH_X1 port map( G => en, D => N92, Q => output(13));
   output_reg_12_inst : DLH_X1 port map( G => en, D => N91, Q => output(12));
   output_reg_11_inst : DLH_X1 port map( G => en, D => N90, Q => output(11));
   output_reg_10_inst : DLH_X1 port map( G => en, D => N89, Q => output(10));
   output_reg_9_inst : DLH_X1 port map( G => en, D => N88, Q => output(9));
   output_reg_8_inst : DLH_X1 port map( G => en, D => N87, Q => output(8));
   output_reg_7_inst : DLH_X1 port map( G => en, D => N86, Q => output(7));
   output_reg_6_inst : DLH_X1 port map( G => en, D => N85, Q => output(6));
   output_reg_5_inst : DLH_X1 port map( G => en, D => N84, Q => output(5));
   output_reg_4_inst : DLH_X1 port map( G => en, D => N83, Q => output(4));
   output_reg_3_inst : DLH_X1 port map( G => en, D => N82, Q => output(3));
   output_reg_2_inst : DLH_X1 port map( G => en, D => N81, Q => output(2));
   output_reg_1_inst : DLH_X1 port map( G => en, D => N80, Q => output(1));
   output_reg_0_inst : DLH_X1 port map( G => en, D => N79, Q => output(0));
   match_dirty_f_reg : DLH_X1 port map( G => en, D => N112, Q => match_dirty_f)
                           ;
   U2 : OAI21_X4 port map( B1 => n38, B2 => n39, A => n36, ZN => n2);
   U3 : AND3_X2 port map( A1 => n36, A2 => n37, A3 => n38, ZN => n4);
   U4 : AND2_X2 port map( A1 => n39, A2 => n36, ZN => n3);
   U5 : INV_X1 port map( A => n1, ZN => N99);
   U6 : AOI222_X1 port map( A1 => reg_c(20), A2 => n2, B1 => reg_f(20), B2 => 
                           n3, C1 => reg_ff(20), C2 => n4, ZN => n1);
   U7 : INV_X1 port map( A => n5, ZN => N98);
   U8 : AOI222_X1 port map( A1 => reg_c(19), A2 => n2, B1 => reg_f(19), B2 => 
                           n3, C1 => reg_ff(19), C2 => n4, ZN => n5);
   U9 : INV_X1 port map( A => n6, ZN => N97);
   U10 : AOI222_X1 port map( A1 => reg_c(18), A2 => n2, B1 => reg_f(18), B2 => 
                           n3, C1 => reg_ff(18), C2 => n4, ZN => n6);
   U11 : INV_X1 port map( A => n7, ZN => N96);
   U12 : AOI222_X1 port map( A1 => reg_c(17), A2 => n2, B1 => reg_f(17), B2 => 
                           n3, C1 => reg_ff(17), C2 => n4, ZN => n7);
   U13 : INV_X1 port map( A => n8, ZN => N95);
   U14 : AOI222_X1 port map( A1 => reg_c(16), A2 => n2, B1 => reg_f(16), B2 => 
                           n3, C1 => reg_ff(16), C2 => n4, ZN => n8);
   U15 : INV_X1 port map( A => n9, ZN => N94);
   U16 : AOI222_X1 port map( A1 => reg_c(15), A2 => n2, B1 => reg_f(15), B2 => 
                           n3, C1 => reg_ff(15), C2 => n4, ZN => n9);
   U17 : INV_X1 port map( A => n10, ZN => N93);
   U18 : AOI222_X1 port map( A1 => reg_c(14), A2 => n2, B1 => reg_f(14), B2 => 
                           n3, C1 => reg_ff(14), C2 => n4, ZN => n10);
   U19 : INV_X1 port map( A => n11, ZN => N92);
   U20 : AOI222_X1 port map( A1 => reg_c(13), A2 => n2, B1 => reg_f(13), B2 => 
                           n3, C1 => reg_ff(13), C2 => n4, ZN => n11);
   U21 : INV_X1 port map( A => n12, ZN => N91);
   U22 : AOI222_X1 port map( A1 => reg_c(12), A2 => n2, B1 => reg_f(12), B2 => 
                           n3, C1 => reg_ff(12), C2 => n4, ZN => n12);
   U23 : INV_X1 port map( A => n13, ZN => N90);
   U24 : AOI222_X1 port map( A1 => reg_c(11), A2 => n2, B1 => reg_f(11), B2 => 
                           n3, C1 => reg_ff(11), C2 => n4, ZN => n13);
   U25 : INV_X1 port map( A => n14, ZN => N89);
   U26 : AOI222_X1 port map( A1 => reg_c(10), A2 => n2, B1 => reg_f(10), B2 => 
                           n3, C1 => reg_ff(10), C2 => n4, ZN => n14);
   U27 : INV_X1 port map( A => n15, ZN => N88);
   U28 : AOI222_X1 port map( A1 => reg_c(9), A2 => n2, B1 => reg_f(9), B2 => n3
                           , C1 => reg_ff(9), C2 => n4, ZN => n15);
   U29 : INV_X1 port map( A => n16, ZN => N87);
   U30 : AOI222_X1 port map( A1 => reg_c(8), A2 => n2, B1 => reg_f(8), B2 => n3
                           , C1 => reg_ff(8), C2 => n4, ZN => n16);
   U31 : INV_X1 port map( A => n17, ZN => N86);
   U32 : AOI222_X1 port map( A1 => reg_c(7), A2 => n2, B1 => reg_f(7), B2 => n3
                           , C1 => reg_ff(7), C2 => n4, ZN => n17);
   U33 : INV_X1 port map( A => n18, ZN => N85);
   U34 : AOI222_X1 port map( A1 => reg_c(6), A2 => n2, B1 => reg_f(6), B2 => n3
                           , C1 => reg_ff(6), C2 => n4, ZN => n18);
   U35 : INV_X1 port map( A => n19, ZN => N84);
   U36 : AOI222_X1 port map( A1 => reg_c(5), A2 => n2, B1 => reg_f(5), B2 => n3
                           , C1 => reg_ff(5), C2 => n4, ZN => n19);
   U37 : INV_X1 port map( A => n20, ZN => N83);
   U38 : AOI222_X1 port map( A1 => reg_c(4), A2 => n2, B1 => reg_f(4), B2 => n3
                           , C1 => reg_ff(4), C2 => n4, ZN => n20);
   U39 : INV_X1 port map( A => n21, ZN => N82);
   U40 : AOI222_X1 port map( A1 => reg_c(3), A2 => n2, B1 => reg_f(3), B2 => n3
                           , C1 => reg_ff(3), C2 => n4, ZN => n21);
   U41 : INV_X1 port map( A => n22, ZN => N81);
   U42 : AOI222_X1 port map( A1 => reg_c(2), A2 => n2, B1 => reg_f(2), B2 => n3
                           , C1 => reg_ff(2), C2 => n4, ZN => n22);
   U43 : INV_X1 port map( A => n23, ZN => N80);
   U44 : AOI222_X1 port map( A1 => reg_c(1), A2 => n2, B1 => reg_f(1), B2 => n3
                           , C1 => reg_ff(1), C2 => n4, ZN => n23);
   U45 : INV_X1 port map( A => n24, ZN => N79);
   U46 : AOI222_X1 port map( A1 => reg_c(0), A2 => n2, B1 => reg_f(0), B2 => n3
                           , C1 => reg_ff(0), C2 => n4, ZN => n24);
   U47 : AND2_X1 port map( A1 => dirty_f, A2 => n3, ZN => N112);
   U48 : AND2_X1 port map( A1 => dirty_ff, A2 => n4, ZN => N111);
   U49 : INV_X1 port map( A => n25, ZN => N110);
   U50 : AOI222_X1 port map( A1 => reg_c(31), A2 => n2, B1 => reg_f(31), B2 => 
                           n3, C1 => reg_ff(31), C2 => n4, ZN => n25);
   U51 : INV_X1 port map( A => n26, ZN => N109);
   U52 : AOI222_X1 port map( A1 => reg_c(30), A2 => n2, B1 => reg_f(30), B2 => 
                           n3, C1 => reg_ff(30), C2 => n4, ZN => n26);
   U53 : INV_X1 port map( A => n27, ZN => N108);
   U54 : AOI222_X1 port map( A1 => reg_c(29), A2 => n2, B1 => reg_f(29), B2 => 
                           n3, C1 => reg_ff(29), C2 => n4, ZN => n27);
   U55 : INV_X1 port map( A => n28, ZN => N107);
   U56 : AOI222_X1 port map( A1 => reg_c(28), A2 => n2, B1 => reg_f(28), B2 => 
                           n3, C1 => reg_ff(28), C2 => n4, ZN => n28);
   U57 : INV_X1 port map( A => n29, ZN => N106);
   U58 : AOI222_X1 port map( A1 => reg_c(27), A2 => n2, B1 => reg_f(27), B2 => 
                           n3, C1 => reg_ff(27), C2 => n4, ZN => n29);
   U59 : INV_X1 port map( A => n30, ZN => N105);
   U60 : AOI222_X1 port map( A1 => reg_c(26), A2 => n2, B1 => reg_f(26), B2 => 
                           n3, C1 => reg_ff(26), C2 => n4, ZN => n30);
   U61 : INV_X1 port map( A => n31, ZN => N104);
   U62 : AOI222_X1 port map( A1 => reg_c(25), A2 => n2, B1 => reg_f(25), B2 => 
                           n3, C1 => reg_ff(25), C2 => n4, ZN => n31);
   U63 : INV_X1 port map( A => n32, ZN => N103);
   U64 : AOI222_X1 port map( A1 => reg_c(24), A2 => n2, B1 => reg_f(24), B2 => 
                           n3, C1 => reg_ff(24), C2 => n4, ZN => n32);
   U65 : INV_X1 port map( A => n33, ZN => N102);
   U66 : AOI222_X1 port map( A1 => reg_c(23), A2 => n2, B1 => reg_f(23), B2 => 
                           n3, C1 => reg_ff(23), C2 => n4, ZN => n33);
   U67 : INV_X1 port map( A => n34, ZN => N101);
   U68 : AOI222_X1 port map( A1 => reg_c(22), A2 => n2, B1 => reg_f(22), B2 => 
                           n3, C1 => reg_ff(22), C2 => n4, ZN => n34);
   U69 : INV_X1 port map( A => n35, ZN => N100);
   U70 : AOI222_X1 port map( A1 => reg_c(21), A2 => n2, B1 => reg_f(21), B2 => 
                           n3, C1 => reg_ff(21), C2 => n4, ZN => n35);
   U71 : NAND4_X1 port map( A1 => n40, A2 => n41, A3 => n42, A4 => n43, ZN => 
                           n36);
   U72 : NOR2_X1 port map( A1 => addr_c(1), A2 => addr_c(0), ZN => n43);
   U73 : INV_X1 port map( A => addr_c(4), ZN => n41);
   U74 : INV_X1 port map( A => n37, ZN => n39);
   U75 : NAND4_X1 port map( A1 => n44, A2 => valid_f, A3 => n45, A4 => n46, ZN 
                           => n37);
   U76 : NOR3_X1 port map( A1 => n47, A2 => n48, A3 => n49, ZN => n46);
   U77 : XOR2_X1 port map( A => addr_f(2), B => addr_c(2), Z => n49);
   U78 : XOR2_X1 port map( A => addr_f(4), B => addr_c(4), Z => n48);
   U79 : XOR2_X1 port map( A => addr_f(3), B => addr_c(3), Z => n47);
   U80 : XNOR2_X1 port map( A => addr_c(0), B => addr_f(0), ZN => n45);
   U81 : XNOR2_X1 port map( A => addr_c(1), B => addr_f(1), ZN => n44);
   U82 : AND4_X1 port map( A1 => n50, A2 => valid_ff, A3 => n51, A4 => n52, ZN 
                           => n38);
   U83 : NOR3_X1 port map( A1 => n53, A2 => n54, A3 => n55, ZN => n52);
   U84 : XOR2_X1 port map( A => addr_ff(0), B => addr_c(0), Z => n55);
   U85 : XOR2_X1 port map( A => addr_ff(1), B => addr_c(1), Z => n54);
   U86 : XOR2_X1 port map( A => addr_ff(4), B => addr_c(4), Z => n53);
   U87 : XOR2_X1 port map( A => n40, B => addr_ff(3), Z => n51);
   U88 : INV_X1 port map( A => addr_c(3), ZN => n40);
   U89 : XOR2_X1 port map( A => n42, B => addr_ff(2), Z => n50);
   U90 : INV_X1 port map( A => addr_c(2), ZN => n42);

end SYN_fwd_mux_2_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE32_12 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 0);
         dout : out std_logic_vector (31 downto 0));

end Reg_DATA_SIZE32_12;

architecture SYN_reg_arch of Reg_DATA_SIZE32_12 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal dout_31_port, dout_30_port, dout_29_port, dout_28_port, dout_27_port,
      dout_26_port, dout_25_port, dout_24_port, dout_23_port, dout_22_port, 
      dout_21_port, dout_20_port, dout_19_port, dout_18_port, dout_17_port, 
      dout_16_port, dout_15_port, dout_14_port, dout_13_port, dout_12_port, 
      dout_11_port, dout_10_port, dout_9_port, dout_8_port, dout_7_port, 
      dout_6_port, dout_5_port, dout_4_port, dout_3_port, dout_2_port, 
      dout_1_port, dout_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, net109161, net109162, net109163, 
      net109164, net109165, net109166, net109167, net109168, net109169, 
      net109170, net109171, net109172, net109173, net109174, net109175, 
      net109176, net109177, net109178, net109179, net109180, net109181, 
      net109182, net109183, net109184, net109185, net109186, net109187, 
      net109188, net109189, net109190, net109191, net109192 : std_logic;

begin
   dout <= ( dout_31_port, dout_30_port, dout_29_port, dout_28_port, 
      dout_27_port, dout_26_port, dout_25_port, dout_24_port, dout_23_port, 
      dout_22_port, dout_21_port, dout_20_port, dout_19_port, dout_18_port, 
      dout_17_port, dout_16_port, dout_15_port, dout_14_port, dout_13_port, 
      dout_12_port, dout_11_port, dout_10_port, dout_9_port, dout_8_port, 
      dout_7_port, dout_6_port, dout_5_port, dout_4_port, dout_3_port, 
      dout_2_port, dout_1_port, dout_0_port );
   
   dout_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           dout_31_port, QN => net109192);
   dout_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           dout_30_port, QN => net109191);
   dout_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           dout_29_port, QN => net109190);
   dout_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           dout_28_port, QN => net109189);
   dout_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           dout_27_port, QN => net109188);
   dout_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => rst, Q => 
                           dout_26_port, QN => net109187);
   dout_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => rst, Q => 
                           dout_25_port, QN => net109186);
   dout_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => rst, Q => 
                           dout_24_port, QN => net109185);
   dout_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => rst, Q => 
                           dout_23_port, QN => net109184);
   dout_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => rst, Q => 
                           dout_22_port, QN => net109183);
   dout_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => rst, Q => 
                           dout_21_port, QN => net109182);
   dout_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => rst, Q => 
                           dout_20_port, QN => net109181);
   dout_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => rst, Q => 
                           dout_19_port, QN => net109180);
   dout_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => rst, Q => 
                           dout_18_port, QN => net109179);
   dout_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => rst, Q => 
                           dout_17_port, QN => net109178);
   dout_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => rst, Q => 
                           dout_16_port, QN => net109177);
   dout_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => rst, Q => 
                           dout_15_port, QN => net109176);
   dout_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => rst, Q => 
                           dout_14_port, QN => net109175);
   dout_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => rst, Q => 
                           dout_13_port, QN => net109174);
   dout_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => rst, Q => 
                           dout_12_port, QN => net109173);
   dout_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => rst, Q => 
                           dout_11_port, QN => net109172);
   dout_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => rst, Q => 
                           dout_10_port, QN => net109171);
   dout_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => rst, Q => 
                           dout_9_port, QN => net109170);
   dout_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => rst, Q => 
                           dout_8_port, QN => net109169);
   dout_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => rst, Q => 
                           dout_7_port, QN => net109168);
   dout_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => rst, Q => 
                           dout_6_port, QN => net109167);
   dout_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => rst, Q => 
                           dout_5_port, QN => net109166);
   dout_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => rst, Q => 
                           dout_4_port, QN => net109165);
   dout_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => rst, Q => 
                           dout_3_port, QN => net109164);
   dout_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => rst, Q => 
                           dout_2_port, QN => net109163);
   dout_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => rst, Q => 
                           dout_1_port, QN => net109162);
   dout_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => rst, Q => 
                           dout_0_port, QN => net109161);
   U2 : MUX2_X1 port map( A => dout_31_port, B => din(31), S => en, Z => n1);
   U3 : MUX2_X1 port map( A => dout_30_port, B => din(30), S => en, Z => n2);
   U4 : MUX2_X1 port map( A => dout_29_port, B => din(29), S => en, Z => n3);
   U5 : MUX2_X1 port map( A => dout_28_port, B => din(28), S => en, Z => n4);
   U6 : MUX2_X1 port map( A => dout_27_port, B => din(27), S => en, Z => n5);
   U7 : MUX2_X1 port map( A => dout_26_port, B => din(26), S => en, Z => n6);
   U8 : MUX2_X1 port map( A => dout_25_port, B => din(25), S => en, Z => n7);
   U9 : MUX2_X1 port map( A => dout_24_port, B => din(24), S => en, Z => n8);
   U10 : MUX2_X1 port map( A => dout_23_port, B => din(23), S => en, Z => n9);
   U11 : MUX2_X1 port map( A => dout_22_port, B => din(22), S => en, Z => n10);
   U12 : MUX2_X1 port map( A => dout_21_port, B => din(21), S => en, Z => n11);
   U13 : MUX2_X1 port map( A => dout_20_port, B => din(20), S => en, Z => n12);
   U14 : MUX2_X1 port map( A => dout_19_port, B => din(19), S => en, Z => n13);
   U15 : MUX2_X1 port map( A => dout_18_port, B => din(18), S => en, Z => n14);
   U16 : MUX2_X1 port map( A => dout_17_port, B => din(17), S => en, Z => n15);
   U17 : MUX2_X1 port map( A => dout_16_port, B => din(16), S => en, Z => n16);
   U18 : MUX2_X1 port map( A => dout_15_port, B => din(15), S => en, Z => n17);
   U19 : MUX2_X1 port map( A => dout_14_port, B => din(14), S => en, Z => n18);
   U20 : MUX2_X1 port map( A => dout_13_port, B => din(13), S => en, Z => n19);
   U21 : MUX2_X1 port map( A => dout_12_port, B => din(12), S => en, Z => n20);
   U22 : MUX2_X1 port map( A => dout_11_port, B => din(11), S => en, Z => n21);
   U23 : MUX2_X1 port map( A => dout_10_port, B => din(10), S => en, Z => n22);
   U24 : MUX2_X1 port map( A => dout_9_port, B => din(9), S => en, Z => n23);
   U25 : MUX2_X1 port map( A => dout_8_port, B => din(8), S => en, Z => n24);
   U26 : MUX2_X1 port map( A => dout_7_port, B => din(7), S => en, Z => n25);
   U27 : MUX2_X1 port map( A => dout_6_port, B => din(6), S => en, Z => n26);
   U28 : MUX2_X1 port map( A => dout_5_port, B => din(5), S => en, Z => n27);
   U29 : MUX2_X1 port map( A => dout_4_port, B => din(4), S => en, Z => n28);
   U30 : MUX2_X1 port map( A => dout_3_port, B => din(3), S => en, Z => n29);
   U31 : MUX2_X1 port map( A => dout_2_port, B => din(2), S => en, Z => n30);
   U32 : MUX2_X1 port map( A => dout_1_port, B => din(1), S => en, Z => n31);
   U33 : MUX2_X1 port map( A => dout_0_port, B => din(0), S => en, Z => n32);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE32_11 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 0);
         dout : out std_logic_vector (31 downto 0));

end Reg_DATA_SIZE32_11;

architecture SYN_reg_arch of Reg_DATA_SIZE32_11 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal dout_31_port, dout_30_port, dout_29_port, dout_28_port, dout_27_port,
      dout_26_port, dout_25_port, dout_24_port, dout_23_port, dout_22_port, 
      dout_21_port, dout_20_port, dout_19_port, dout_18_port, dout_17_port, 
      dout_16_port, dout_15_port, dout_14_port, dout_13_port, dout_12_port, 
      dout_11_port, dout_10_port, dout_9_port, dout_8_port, dout_7_port, 
      dout_6_port, dout_5_port, dout_4_port, dout_3_port, dout_2_port, 
      dout_1_port, dout_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, net109129, net109130, net109131, 
      net109132, net109133, net109134, net109135, net109136, net109137, 
      net109138, net109139, net109140, net109141, net109142, net109143, 
      net109144, net109145, net109146, net109147, net109148, net109149, 
      net109150, net109151, net109152, net109153, net109154, net109155, 
      net109156, net109157, net109158, net109159, net109160 : std_logic;

begin
   dout <= ( dout_31_port, dout_30_port, dout_29_port, dout_28_port, 
      dout_27_port, dout_26_port, dout_25_port, dout_24_port, dout_23_port, 
      dout_22_port, dout_21_port, dout_20_port, dout_19_port, dout_18_port, 
      dout_17_port, dout_16_port, dout_15_port, dout_14_port, dout_13_port, 
      dout_12_port, dout_11_port, dout_10_port, dout_9_port, dout_8_port, 
      dout_7_port, dout_6_port, dout_5_port, dout_4_port, dout_3_port, 
      dout_2_port, dout_1_port, dout_0_port );
   
   dout_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           dout_31_port, QN => net109160);
   dout_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           dout_30_port, QN => net109159);
   dout_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           dout_29_port, QN => net109158);
   dout_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           dout_28_port, QN => net109157);
   dout_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           dout_27_port, QN => net109156);
   dout_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => rst, Q => 
                           dout_26_port, QN => net109155);
   dout_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => rst, Q => 
                           dout_25_port, QN => net109154);
   dout_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => rst, Q => 
                           dout_24_port, QN => net109153);
   dout_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => rst, Q => 
                           dout_23_port, QN => net109152);
   dout_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => rst, Q => 
                           dout_22_port, QN => net109151);
   dout_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => rst, Q => 
                           dout_21_port, QN => net109150);
   dout_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => rst, Q => 
                           dout_20_port, QN => net109149);
   dout_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => rst, Q => 
                           dout_19_port, QN => net109148);
   dout_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => rst, Q => 
                           dout_18_port, QN => net109147);
   dout_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => rst, Q => 
                           dout_17_port, QN => net109146);
   dout_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => rst, Q => 
                           dout_16_port, QN => net109145);
   dout_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => rst, Q => 
                           dout_15_port, QN => net109144);
   dout_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => rst, Q => 
                           dout_14_port, QN => net109143);
   dout_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => rst, Q => 
                           dout_13_port, QN => net109142);
   dout_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => rst, Q => 
                           dout_12_port, QN => net109141);
   dout_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => rst, Q => 
                           dout_11_port, QN => net109140);
   dout_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => rst, Q => 
                           dout_10_port, QN => net109139);
   dout_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => rst, Q => 
                           dout_9_port, QN => net109138);
   dout_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => rst, Q => 
                           dout_8_port, QN => net109137);
   dout_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => rst, Q => 
                           dout_7_port, QN => net109136);
   dout_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => rst, Q => 
                           dout_6_port, QN => net109135);
   dout_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => rst, Q => 
                           dout_5_port, QN => net109134);
   dout_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => rst, Q => 
                           dout_4_port, QN => net109133);
   dout_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => rst, Q => 
                           dout_3_port, QN => net109132);
   dout_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => rst, Q => 
                           dout_2_port, QN => net109131);
   dout_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => rst, Q => 
                           dout_1_port, QN => net109130);
   dout_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => rst, Q => 
                           dout_0_port, QN => net109129);
   U2 : MUX2_X1 port map( A => dout_31_port, B => din(31), S => en, Z => n1);
   U3 : MUX2_X1 port map( A => dout_30_port, B => din(30), S => en, Z => n2);
   U4 : MUX2_X1 port map( A => dout_29_port, B => din(29), S => en, Z => n3);
   U5 : MUX2_X1 port map( A => dout_28_port, B => din(28), S => en, Z => n4);
   U6 : MUX2_X1 port map( A => dout_27_port, B => din(27), S => en, Z => n5);
   U7 : MUX2_X1 port map( A => dout_26_port, B => din(26), S => en, Z => n6);
   U8 : MUX2_X1 port map( A => dout_25_port, B => din(25), S => en, Z => n7);
   U9 : MUX2_X1 port map( A => dout_24_port, B => din(24), S => en, Z => n8);
   U10 : MUX2_X1 port map( A => dout_23_port, B => din(23), S => en, Z => n9);
   U11 : MUX2_X1 port map( A => dout_22_port, B => din(22), S => en, Z => n10);
   U12 : MUX2_X1 port map( A => dout_21_port, B => din(21), S => en, Z => n11);
   U13 : MUX2_X1 port map( A => dout_20_port, B => din(20), S => en, Z => n12);
   U14 : MUX2_X1 port map( A => dout_19_port, B => din(19), S => en, Z => n13);
   U15 : MUX2_X1 port map( A => dout_18_port, B => din(18), S => en, Z => n14);
   U16 : MUX2_X1 port map( A => dout_17_port, B => din(17), S => en, Z => n15);
   U17 : MUX2_X1 port map( A => dout_16_port, B => din(16), S => en, Z => n16);
   U18 : MUX2_X1 port map( A => dout_15_port, B => din(15), S => en, Z => n17);
   U19 : MUX2_X1 port map( A => dout_14_port, B => din(14), S => en, Z => n18);
   U20 : MUX2_X1 port map( A => dout_13_port, B => din(13), S => en, Z => n19);
   U21 : MUX2_X1 port map( A => dout_12_port, B => din(12), S => en, Z => n20);
   U22 : MUX2_X1 port map( A => dout_11_port, B => din(11), S => en, Z => n21);
   U23 : MUX2_X1 port map( A => dout_10_port, B => din(10), S => en, Z => n22);
   U24 : MUX2_X1 port map( A => dout_9_port, B => din(9), S => en, Z => n23);
   U25 : MUX2_X1 port map( A => dout_8_port, B => din(8), S => en, Z => n24);
   U26 : MUX2_X1 port map( A => dout_7_port, B => din(7), S => en, Z => n25);
   U27 : MUX2_X1 port map( A => dout_6_port, B => din(6), S => en, Z => n26);
   U28 : MUX2_X1 port map( A => dout_5_port, B => din(5), S => en, Z => n27);
   U29 : MUX2_X1 port map( A => dout_4_port, B => din(4), S => en, Z => n28);
   U30 : MUX2_X1 port map( A => dout_3_port, B => din(3), S => en, Z => n29);
   U31 : MUX2_X1 port map( A => dout_2_port, B => din(2), S => en, Z => n30);
   U32 : MUX2_X1 port map( A => dout_1_port, B => din(1), S => en, Z => n31);
   U33 : MUX2_X1 port map( A => dout_0_port, B => din(0), S => en, Z => n32);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE32_10 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 0);
         dout : out std_logic_vector (31 downto 0));

end Reg_DATA_SIZE32_10;

architecture SYN_reg_arch of Reg_DATA_SIZE32_10 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal dout_31_port, dout_30_port, dout_29_port, dout_28_port, dout_27_port,
      dout_26_port, dout_25_port, dout_24_port, dout_23_port, dout_22_port, 
      dout_21_port, dout_20_port, dout_19_port, dout_18_port, dout_17_port, 
      dout_16_port, dout_15_port, dout_14_port, dout_13_port, dout_12_port, 
      dout_11_port, dout_10_port, dout_9_port, dout_8_port, dout_7_port, 
      dout_6_port, dout_5_port, dout_4_port, dout_3_port, dout_2_port, 
      dout_1_port, dout_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, net109097, net109098, net109099, 
      net109100, net109101, net109102, net109103, net109104, net109105, 
      net109106, net109107, net109108, net109109, net109110, net109111, 
      net109112, net109113, net109114, net109115, net109116, net109117, 
      net109118, net109119, net109120, net109121, net109122, net109123, 
      net109124, net109125, net109126, net109127, net109128 : std_logic;

begin
   dout <= ( dout_31_port, dout_30_port, dout_29_port, dout_28_port, 
      dout_27_port, dout_26_port, dout_25_port, dout_24_port, dout_23_port, 
      dout_22_port, dout_21_port, dout_20_port, dout_19_port, dout_18_port, 
      dout_17_port, dout_16_port, dout_15_port, dout_14_port, dout_13_port, 
      dout_12_port, dout_11_port, dout_10_port, dout_9_port, dout_8_port, 
      dout_7_port, dout_6_port, dout_5_port, dout_4_port, dout_3_port, 
      dout_2_port, dout_1_port, dout_0_port );
   
   dout_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           dout_31_port, QN => net109128);
   dout_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           dout_30_port, QN => net109127);
   dout_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           dout_29_port, QN => net109126);
   dout_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           dout_28_port, QN => net109125);
   dout_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           dout_27_port, QN => net109124);
   dout_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => rst, Q => 
                           dout_26_port, QN => net109123);
   dout_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => rst, Q => 
                           dout_25_port, QN => net109122);
   dout_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => rst, Q => 
                           dout_24_port, QN => net109121);
   dout_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => rst, Q => 
                           dout_23_port, QN => net109120);
   dout_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => rst, Q => 
                           dout_22_port, QN => net109119);
   dout_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => rst, Q => 
                           dout_21_port, QN => net109118);
   dout_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => rst, Q => 
                           dout_20_port, QN => net109117);
   dout_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => rst, Q => 
                           dout_19_port, QN => net109116);
   dout_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => rst, Q => 
                           dout_18_port, QN => net109115);
   dout_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => rst, Q => 
                           dout_17_port, QN => net109114);
   dout_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => rst, Q => 
                           dout_16_port, QN => net109113);
   dout_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => rst, Q => 
                           dout_15_port, QN => net109112);
   dout_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => rst, Q => 
                           dout_14_port, QN => net109111);
   dout_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => rst, Q => 
                           dout_13_port, QN => net109110);
   dout_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => rst, Q => 
                           dout_12_port, QN => net109109);
   dout_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => rst, Q => 
                           dout_11_port, QN => net109108);
   dout_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => rst, Q => 
                           dout_10_port, QN => net109107);
   dout_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => rst, Q => 
                           dout_9_port, QN => net109106);
   dout_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => rst, Q => 
                           dout_8_port, QN => net109105);
   dout_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => rst, Q => 
                           dout_7_port, QN => net109104);
   dout_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => rst, Q => 
                           dout_6_port, QN => net109103);
   dout_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => rst, Q => 
                           dout_5_port, QN => net109102);
   dout_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => rst, Q => 
                           dout_4_port, QN => net109101);
   dout_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => rst, Q => 
                           dout_3_port, QN => net109100);
   dout_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => rst, Q => 
                           dout_2_port, QN => net109099);
   dout_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => rst, Q => 
                           dout_1_port, QN => net109098);
   dout_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => rst, Q => 
                           dout_0_port, QN => net109097);
   U2 : MUX2_X1 port map( A => dout_31_port, B => din(31), S => en, Z => n1);
   U3 : MUX2_X1 port map( A => dout_30_port, B => din(30), S => en, Z => n2);
   U4 : MUX2_X1 port map( A => dout_29_port, B => din(29), S => en, Z => n3);
   U5 : MUX2_X1 port map( A => dout_28_port, B => din(28), S => en, Z => n4);
   U6 : MUX2_X1 port map( A => dout_27_port, B => din(27), S => en, Z => n5);
   U7 : MUX2_X1 port map( A => dout_26_port, B => din(26), S => en, Z => n6);
   U8 : MUX2_X1 port map( A => dout_25_port, B => din(25), S => en, Z => n7);
   U9 : MUX2_X1 port map( A => dout_24_port, B => din(24), S => en, Z => n8);
   U10 : MUX2_X1 port map( A => dout_23_port, B => din(23), S => en, Z => n9);
   U11 : MUX2_X1 port map( A => dout_22_port, B => din(22), S => en, Z => n10);
   U12 : MUX2_X1 port map( A => dout_21_port, B => din(21), S => en, Z => n11);
   U13 : MUX2_X1 port map( A => dout_20_port, B => din(20), S => en, Z => n12);
   U14 : MUX2_X1 port map( A => dout_19_port, B => din(19), S => en, Z => n13);
   U15 : MUX2_X1 port map( A => dout_18_port, B => din(18), S => en, Z => n14);
   U16 : MUX2_X1 port map( A => dout_17_port, B => din(17), S => en, Z => n15);
   U17 : MUX2_X1 port map( A => dout_16_port, B => din(16), S => en, Z => n16);
   U18 : MUX2_X1 port map( A => dout_15_port, B => din(15), S => en, Z => n17);
   U19 : MUX2_X1 port map( A => dout_14_port, B => din(14), S => en, Z => n18);
   U20 : MUX2_X1 port map( A => dout_13_port, B => din(13), S => en, Z => n19);
   U21 : MUX2_X1 port map( A => dout_12_port, B => din(12), S => en, Z => n20);
   U22 : MUX2_X1 port map( A => dout_11_port, B => din(11), S => en, Z => n21);
   U23 : MUX2_X1 port map( A => dout_10_port, B => din(10), S => en, Z => n22);
   U24 : MUX2_X1 port map( A => dout_9_port, B => din(9), S => en, Z => n23);
   U25 : MUX2_X1 port map( A => dout_8_port, B => din(8), S => en, Z => n24);
   U26 : MUX2_X1 port map( A => dout_7_port, B => din(7), S => en, Z => n25);
   U27 : MUX2_X1 port map( A => dout_6_port, B => din(6), S => en, Z => n26);
   U28 : MUX2_X1 port map( A => dout_5_port, B => din(5), S => en, Z => n27);
   U29 : MUX2_X1 port map( A => dout_4_port, B => din(4), S => en, Z => n28);
   U30 : MUX2_X1 port map( A => dout_3_port, B => din(3), S => en, Z => n29);
   U31 : MUX2_X1 port map( A => dout_2_port, B => din(2), S => en, Z => n30);
   U32 : MUX2_X1 port map( A => dout_1_port, B => din(1), S => en, Z => n31);
   U33 : MUX2_X1 port map( A => dout_0_port, B => din(0), S => en, Z => n32);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE32_9 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 0);
         dout : out std_logic_vector (31 downto 0));

end Reg_DATA_SIZE32_9;

architecture SYN_reg_arch of Reg_DATA_SIZE32_9 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal dout_31_port, dout_30_port, dout_29_port, dout_28_port, dout_27_port,
      dout_26_port, dout_25_port, dout_24_port, dout_23_port, dout_22_port, 
      dout_21_port, dout_20_port, dout_19_port, dout_18_port, dout_17_port, 
      dout_16_port, dout_15_port, dout_14_port, dout_13_port, dout_12_port, 
      dout_11_port, dout_10_port, dout_9_port, dout_8_port, dout_7_port, 
      dout_6_port, dout_5_port, dout_4_port, dout_3_port, dout_2_port, 
      dout_1_port, dout_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, net109065, net109066, net109067, 
      net109068, net109069, net109070, net109071, net109072, net109073, 
      net109074, net109075, net109076, net109077, net109078, net109079, 
      net109080, net109081, net109082, net109083, net109084, net109085, 
      net109086, net109087, net109088, net109089, net109090, net109091, 
      net109092, net109093, net109094, net109095, net109096 : std_logic;

begin
   dout <= ( dout_31_port, dout_30_port, dout_29_port, dout_28_port, 
      dout_27_port, dout_26_port, dout_25_port, dout_24_port, dout_23_port, 
      dout_22_port, dout_21_port, dout_20_port, dout_19_port, dout_18_port, 
      dout_17_port, dout_16_port, dout_15_port, dout_14_port, dout_13_port, 
      dout_12_port, dout_11_port, dout_10_port, dout_9_port, dout_8_port, 
      dout_7_port, dout_6_port, dout_5_port, dout_4_port, dout_3_port, 
      dout_2_port, dout_1_port, dout_0_port );
   
   dout_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           dout_31_port, QN => net109096);
   dout_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           dout_30_port, QN => net109095);
   dout_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           dout_29_port, QN => net109094);
   dout_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           dout_28_port, QN => net109093);
   dout_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           dout_27_port, QN => net109092);
   dout_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => rst, Q => 
                           dout_26_port, QN => net109091);
   dout_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => rst, Q => 
                           dout_25_port, QN => net109090);
   dout_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => rst, Q => 
                           dout_24_port, QN => net109089);
   dout_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => rst, Q => 
                           dout_23_port, QN => net109088);
   dout_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => rst, Q => 
                           dout_22_port, QN => net109087);
   dout_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => rst, Q => 
                           dout_21_port, QN => net109086);
   dout_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => rst, Q => 
                           dout_20_port, QN => net109085);
   dout_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => rst, Q => 
                           dout_19_port, QN => net109084);
   dout_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => rst, Q => 
                           dout_18_port, QN => net109083);
   dout_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => rst, Q => 
                           dout_17_port, QN => net109082);
   dout_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => rst, Q => 
                           dout_16_port, QN => net109081);
   dout_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => rst, Q => 
                           dout_15_port, QN => net109080);
   dout_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => rst, Q => 
                           dout_14_port, QN => net109079);
   dout_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => rst, Q => 
                           dout_13_port, QN => net109078);
   dout_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => rst, Q => 
                           dout_12_port, QN => net109077);
   dout_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => rst, Q => 
                           dout_11_port, QN => net109076);
   dout_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => rst, Q => 
                           dout_10_port, QN => net109075);
   dout_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => rst, Q => 
                           dout_9_port, QN => net109074);
   dout_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => rst, Q => 
                           dout_8_port, QN => net109073);
   dout_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => rst, Q => 
                           dout_7_port, QN => net109072);
   dout_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => rst, Q => 
                           dout_6_port, QN => net109071);
   dout_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => rst, Q => 
                           dout_5_port, QN => net109070);
   dout_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => rst, Q => 
                           dout_4_port, QN => net109069);
   dout_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => rst, Q => 
                           dout_3_port, QN => net109068);
   dout_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => rst, Q => 
                           dout_2_port, QN => net109067);
   dout_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => rst, Q => 
                           dout_1_port, QN => net109066);
   dout_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => rst, Q => 
                           dout_0_port, QN => net109065);
   U2 : MUX2_X1 port map( A => dout_31_port, B => din(31), S => en, Z => n1);
   U3 : MUX2_X1 port map( A => dout_30_port, B => din(30), S => en, Z => n2);
   U4 : MUX2_X1 port map( A => dout_29_port, B => din(29), S => en, Z => n3);
   U5 : MUX2_X1 port map( A => dout_28_port, B => din(28), S => en, Z => n4);
   U6 : MUX2_X1 port map( A => dout_27_port, B => din(27), S => en, Z => n5);
   U7 : MUX2_X1 port map( A => dout_26_port, B => din(26), S => en, Z => n6);
   U8 : MUX2_X1 port map( A => dout_25_port, B => din(25), S => en, Z => n7);
   U9 : MUX2_X1 port map( A => dout_24_port, B => din(24), S => en, Z => n8);
   U10 : MUX2_X1 port map( A => dout_23_port, B => din(23), S => en, Z => n9);
   U11 : MUX2_X1 port map( A => dout_22_port, B => din(22), S => en, Z => n10);
   U12 : MUX2_X1 port map( A => dout_21_port, B => din(21), S => en, Z => n11);
   U13 : MUX2_X1 port map( A => dout_20_port, B => din(20), S => en, Z => n12);
   U14 : MUX2_X1 port map( A => dout_19_port, B => din(19), S => en, Z => n13);
   U15 : MUX2_X1 port map( A => dout_18_port, B => din(18), S => en, Z => n14);
   U16 : MUX2_X1 port map( A => dout_17_port, B => din(17), S => en, Z => n15);
   U17 : MUX2_X1 port map( A => dout_16_port, B => din(16), S => en, Z => n16);
   U18 : MUX2_X1 port map( A => dout_15_port, B => din(15), S => en, Z => n17);
   U19 : MUX2_X1 port map( A => dout_14_port, B => din(14), S => en, Z => n18);
   U20 : MUX2_X1 port map( A => dout_13_port, B => din(13), S => en, Z => n19);
   U21 : MUX2_X1 port map( A => dout_12_port, B => din(12), S => en, Z => n20);
   U22 : MUX2_X1 port map( A => dout_11_port, B => din(11), S => en, Z => n21);
   U23 : MUX2_X1 port map( A => dout_10_port, B => din(10), S => en, Z => n22);
   U24 : MUX2_X1 port map( A => dout_9_port, B => din(9), S => en, Z => n23);
   U25 : MUX2_X1 port map( A => dout_8_port, B => din(8), S => en, Z => n24);
   U26 : MUX2_X1 port map( A => dout_7_port, B => din(7), S => en, Z => n25);
   U27 : MUX2_X1 port map( A => dout_6_port, B => din(6), S => en, Z => n26);
   U28 : MUX2_X1 port map( A => dout_5_port, B => din(5), S => en, Z => n27);
   U29 : MUX2_X1 port map( A => dout_4_port, B => din(4), S => en, Z => n28);
   U30 : MUX2_X1 port map( A => dout_3_port, B => din(3), S => en, Z => n29);
   U31 : MUX2_X1 port map( A => dout_2_port, B => din(2), S => en, Z => n30);
   U32 : MUX2_X1 port map( A => dout_1_port, B => din(1), S => en, Z => n31);
   U33 : MUX2_X1 port map( A => dout_0_port, B => din(0), S => en, Z => n32);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE32_8 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 0);
         dout : out std_logic_vector (31 downto 0));

end Reg_DATA_SIZE32_8;

architecture SYN_reg_arch of Reg_DATA_SIZE32_8 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal dout_31_port, dout_30_port, dout_29_port, dout_28_port, dout_27_port,
      dout_26_port, dout_25_port, dout_24_port, dout_23_port, dout_22_port, 
      dout_21_port, dout_20_port, dout_19_port, dout_18_port, dout_17_port, 
      dout_16_port, dout_15_port, dout_14_port, dout_13_port, dout_12_port, 
      dout_11_port, dout_10_port, dout_9_port, dout_8_port, dout_7_port, 
      dout_6_port, dout_5_port, dout_4_port, dout_3_port, dout_2_port, 
      dout_1_port, dout_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, net109033, net109034, net109035, 
      net109036, net109037, net109038, net109039, net109040, net109041, 
      net109042, net109043, net109044, net109045, net109046, net109047, 
      net109048, net109049, net109050, net109051, net109052, net109053, 
      net109054, net109055, net109056, net109057, net109058, net109059, 
      net109060, net109061, net109062, net109063, net109064 : std_logic;

begin
   dout <= ( dout_31_port, dout_30_port, dout_29_port, dout_28_port, 
      dout_27_port, dout_26_port, dout_25_port, dout_24_port, dout_23_port, 
      dout_22_port, dout_21_port, dout_20_port, dout_19_port, dout_18_port, 
      dout_17_port, dout_16_port, dout_15_port, dout_14_port, dout_13_port, 
      dout_12_port, dout_11_port, dout_10_port, dout_9_port, dout_8_port, 
      dout_7_port, dout_6_port, dout_5_port, dout_4_port, dout_3_port, 
      dout_2_port, dout_1_port, dout_0_port );
   
   dout_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           dout_31_port, QN => net109064);
   dout_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           dout_30_port, QN => net109063);
   dout_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           dout_29_port, QN => net109062);
   dout_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           dout_28_port, QN => net109061);
   dout_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           dout_27_port, QN => net109060);
   dout_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => rst, Q => 
                           dout_26_port, QN => net109059);
   dout_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => rst, Q => 
                           dout_25_port, QN => net109058);
   dout_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => rst, Q => 
                           dout_24_port, QN => net109057);
   dout_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => rst, Q => 
                           dout_23_port, QN => net109056);
   dout_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => rst, Q => 
                           dout_22_port, QN => net109055);
   dout_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => rst, Q => 
                           dout_21_port, QN => net109054);
   dout_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => rst, Q => 
                           dout_20_port, QN => net109053);
   dout_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => rst, Q => 
                           dout_19_port, QN => net109052);
   dout_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => rst, Q => 
                           dout_18_port, QN => net109051);
   dout_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => rst, Q => 
                           dout_17_port, QN => net109050);
   dout_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => rst, Q => 
                           dout_16_port, QN => net109049);
   dout_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => rst, Q => 
                           dout_15_port, QN => net109048);
   dout_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => rst, Q => 
                           dout_14_port, QN => net109047);
   dout_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => rst, Q => 
                           dout_13_port, QN => net109046);
   dout_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => rst, Q => 
                           dout_12_port, QN => net109045);
   dout_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => rst, Q => 
                           dout_11_port, QN => net109044);
   dout_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => rst, Q => 
                           dout_10_port, QN => net109043);
   dout_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => rst, Q => 
                           dout_9_port, QN => net109042);
   dout_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => rst, Q => 
                           dout_8_port, QN => net109041);
   dout_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => rst, Q => 
                           dout_7_port, QN => net109040);
   dout_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => rst, Q => 
                           dout_6_port, QN => net109039);
   dout_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => rst, Q => 
                           dout_5_port, QN => net109038);
   dout_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => rst, Q => 
                           dout_4_port, QN => net109037);
   dout_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => rst, Q => 
                           dout_3_port, QN => net109036);
   dout_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => rst, Q => 
                           dout_2_port, QN => net109035);
   dout_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => rst, Q => 
                           dout_1_port, QN => net109034);
   dout_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => rst, Q => 
                           dout_0_port, QN => net109033);
   U2 : MUX2_X1 port map( A => dout_31_port, B => din(31), S => en, Z => n1);
   U3 : MUX2_X1 port map( A => dout_30_port, B => din(30), S => en, Z => n2);
   U4 : MUX2_X1 port map( A => dout_29_port, B => din(29), S => en, Z => n3);
   U5 : MUX2_X1 port map( A => dout_28_port, B => din(28), S => en, Z => n4);
   U6 : MUX2_X1 port map( A => dout_27_port, B => din(27), S => en, Z => n5);
   U7 : MUX2_X1 port map( A => dout_26_port, B => din(26), S => en, Z => n6);
   U8 : MUX2_X1 port map( A => dout_25_port, B => din(25), S => en, Z => n7);
   U9 : MUX2_X1 port map( A => dout_24_port, B => din(24), S => en, Z => n8);
   U10 : MUX2_X1 port map( A => dout_23_port, B => din(23), S => en, Z => n9);
   U11 : MUX2_X1 port map( A => dout_22_port, B => din(22), S => en, Z => n10);
   U12 : MUX2_X1 port map( A => dout_21_port, B => din(21), S => en, Z => n11);
   U13 : MUX2_X1 port map( A => dout_20_port, B => din(20), S => en, Z => n12);
   U14 : MUX2_X1 port map( A => dout_19_port, B => din(19), S => en, Z => n13);
   U15 : MUX2_X1 port map( A => dout_18_port, B => din(18), S => en, Z => n14);
   U16 : MUX2_X1 port map( A => dout_17_port, B => din(17), S => en, Z => n15);
   U17 : MUX2_X1 port map( A => dout_16_port, B => din(16), S => en, Z => n16);
   U18 : MUX2_X1 port map( A => dout_15_port, B => din(15), S => en, Z => n17);
   U19 : MUX2_X1 port map( A => dout_14_port, B => din(14), S => en, Z => n18);
   U20 : MUX2_X1 port map( A => dout_13_port, B => din(13), S => en, Z => n19);
   U21 : MUX2_X1 port map( A => dout_12_port, B => din(12), S => en, Z => n20);
   U22 : MUX2_X1 port map( A => dout_11_port, B => din(11), S => en, Z => n21);
   U23 : MUX2_X1 port map( A => dout_10_port, B => din(10), S => en, Z => n22);
   U24 : MUX2_X1 port map( A => dout_9_port, B => din(9), S => en, Z => n23);
   U25 : MUX2_X1 port map( A => dout_8_port, B => din(8), S => en, Z => n24);
   U26 : MUX2_X1 port map( A => dout_7_port, B => din(7), S => en, Z => n25);
   U27 : MUX2_X1 port map( A => dout_6_port, B => din(6), S => en, Z => n26);
   U28 : MUX2_X1 port map( A => dout_5_port, B => din(5), S => en, Z => n27);
   U29 : MUX2_X1 port map( A => dout_4_port, B => din(4), S => en, Z => n28);
   U30 : MUX2_X1 port map( A => dout_3_port, B => din(3), S => en, Z => n29);
   U31 : MUX2_X1 port map( A => dout_2_port, B => din(2), S => en, Z => n30);
   U32 : MUX2_X1 port map( A => dout_1_port, B => din(1), S => en, Z => n31);
   U33 : MUX2_X1 port map( A => dout_0_port, B => din(0), S => en, Z => n32);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE32_7 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 0);
         dout : out std_logic_vector (31 downto 0));

end Reg_DATA_SIZE32_7;

architecture SYN_reg_arch of Reg_DATA_SIZE32_7 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal dout_31_port, dout_30_port, dout_29_port, dout_28_port, dout_27_port,
      dout_26_port, dout_25_port, dout_24_port, dout_23_port, dout_22_port, 
      dout_21_port, dout_20_port, dout_19_port, dout_18_port, dout_17_port, 
      dout_16_port, dout_15_port, dout_14_port, dout_13_port, dout_12_port, 
      dout_11_port, dout_10_port, dout_9_port, dout_8_port, dout_7_port, 
      dout_6_port, dout_5_port, dout_4_port, dout_3_port, dout_2_port, 
      dout_1_port, dout_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, net109001, net109002, net109003, 
      net109004, net109005, net109006, net109007, net109008, net109009, 
      net109010, net109011, net109012, net109013, net109014, net109015, 
      net109016, net109017, net109018, net109019, net109020, net109021, 
      net109022, net109023, net109024, net109025, net109026, net109027, 
      net109028, net109029, net109030, net109031, net109032 : std_logic;

begin
   dout <= ( dout_31_port, dout_30_port, dout_29_port, dout_28_port, 
      dout_27_port, dout_26_port, dout_25_port, dout_24_port, dout_23_port, 
      dout_22_port, dout_21_port, dout_20_port, dout_19_port, dout_18_port, 
      dout_17_port, dout_16_port, dout_15_port, dout_14_port, dout_13_port, 
      dout_12_port, dout_11_port, dout_10_port, dout_9_port, dout_8_port, 
      dout_7_port, dout_6_port, dout_5_port, dout_4_port, dout_3_port, 
      dout_2_port, dout_1_port, dout_0_port );
   
   dout_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           dout_31_port, QN => net109032);
   dout_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           dout_30_port, QN => net109031);
   dout_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           dout_29_port, QN => net109030);
   dout_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           dout_28_port, QN => net109029);
   dout_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           dout_27_port, QN => net109028);
   dout_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => rst, Q => 
                           dout_26_port, QN => net109027);
   dout_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => rst, Q => 
                           dout_25_port, QN => net109026);
   dout_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => rst, Q => 
                           dout_24_port, QN => net109025);
   dout_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => rst, Q => 
                           dout_23_port, QN => net109024);
   dout_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => rst, Q => 
                           dout_22_port, QN => net109023);
   dout_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => rst, Q => 
                           dout_21_port, QN => net109022);
   dout_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => rst, Q => 
                           dout_20_port, QN => net109021);
   dout_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => rst, Q => 
                           dout_19_port, QN => net109020);
   dout_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => rst, Q => 
                           dout_18_port, QN => net109019);
   dout_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => rst, Q => 
                           dout_17_port, QN => net109018);
   dout_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => rst, Q => 
                           dout_16_port, QN => net109017);
   dout_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => rst, Q => 
                           dout_15_port, QN => net109016);
   dout_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => rst, Q => 
                           dout_14_port, QN => net109015);
   dout_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => rst, Q => 
                           dout_13_port, QN => net109014);
   dout_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => rst, Q => 
                           dout_12_port, QN => net109013);
   dout_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => rst, Q => 
                           dout_11_port, QN => net109012);
   dout_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => rst, Q => 
                           dout_10_port, QN => net109011);
   dout_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => rst, Q => 
                           dout_9_port, QN => net109010);
   dout_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => rst, Q => 
                           dout_8_port, QN => net109009);
   dout_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => rst, Q => 
                           dout_7_port, QN => net109008);
   dout_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => rst, Q => 
                           dout_6_port, QN => net109007);
   dout_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => rst, Q => 
                           dout_5_port, QN => net109006);
   dout_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => rst, Q => 
                           dout_4_port, QN => net109005);
   dout_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => rst, Q => 
                           dout_3_port, QN => net109004);
   dout_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => rst, Q => 
                           dout_2_port, QN => net109003);
   dout_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => rst, Q => 
                           dout_1_port, QN => net109002);
   dout_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => rst, Q => 
                           dout_0_port, QN => net109001);
   U2 : MUX2_X1 port map( A => dout_31_port, B => din(31), S => en, Z => n1);
   U3 : MUX2_X1 port map( A => dout_30_port, B => din(30), S => en, Z => n2);
   U4 : MUX2_X1 port map( A => dout_29_port, B => din(29), S => en, Z => n3);
   U5 : MUX2_X1 port map( A => dout_28_port, B => din(28), S => en, Z => n4);
   U6 : MUX2_X1 port map( A => dout_27_port, B => din(27), S => en, Z => n5);
   U7 : MUX2_X1 port map( A => dout_26_port, B => din(26), S => en, Z => n6);
   U8 : MUX2_X1 port map( A => dout_25_port, B => din(25), S => en, Z => n7);
   U9 : MUX2_X1 port map( A => dout_24_port, B => din(24), S => en, Z => n8);
   U10 : MUX2_X1 port map( A => dout_23_port, B => din(23), S => en, Z => n9);
   U11 : MUX2_X1 port map( A => dout_22_port, B => din(22), S => en, Z => n10);
   U12 : MUX2_X1 port map( A => dout_21_port, B => din(21), S => en, Z => n11);
   U13 : MUX2_X1 port map( A => dout_20_port, B => din(20), S => en, Z => n12);
   U14 : MUX2_X1 port map( A => dout_19_port, B => din(19), S => en, Z => n13);
   U15 : MUX2_X1 port map( A => dout_18_port, B => din(18), S => en, Z => n14);
   U16 : MUX2_X1 port map( A => dout_17_port, B => din(17), S => en, Z => n15);
   U17 : MUX2_X1 port map( A => dout_16_port, B => din(16), S => en, Z => n16);
   U18 : MUX2_X1 port map( A => dout_15_port, B => din(15), S => en, Z => n17);
   U19 : MUX2_X1 port map( A => dout_14_port, B => din(14), S => en, Z => n18);
   U20 : MUX2_X1 port map( A => dout_13_port, B => din(13), S => en, Z => n19);
   U21 : MUX2_X1 port map( A => dout_12_port, B => din(12), S => en, Z => n20);
   U22 : MUX2_X1 port map( A => dout_11_port, B => din(11), S => en, Z => n21);
   U23 : MUX2_X1 port map( A => dout_10_port, B => din(10), S => en, Z => n22);
   U24 : MUX2_X1 port map( A => dout_9_port, B => din(9), S => en, Z => n23);
   U25 : MUX2_X1 port map( A => dout_8_port, B => din(8), S => en, Z => n24);
   U26 : MUX2_X1 port map( A => dout_7_port, B => din(7), S => en, Z => n25);
   U27 : MUX2_X1 port map( A => dout_6_port, B => din(6), S => en, Z => n26);
   U28 : MUX2_X1 port map( A => dout_5_port, B => din(5), S => en, Z => n27);
   U29 : MUX2_X1 port map( A => dout_4_port, B => din(4), S => en, Z => n28);
   U30 : MUX2_X1 port map( A => dout_3_port, B => din(3), S => en, Z => n29);
   U31 : MUX2_X1 port map( A => dout_2_port, B => din(2), S => en, Z => n30);
   U32 : MUX2_X1 port map( A => dout_1_port, B => din(1), S => en, Z => n31);
   U33 : MUX2_X1 port map( A => dout_0_port, B => din(0), S => en, Z => n32);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE32_6 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 0);
         dout : out std_logic_vector (31 downto 0));

end Reg_DATA_SIZE32_6;

architecture SYN_reg_arch of Reg_DATA_SIZE32_6 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal dout_31_port, dout_30_port, dout_29_port, dout_28_port, dout_27_port,
      dout_26_port, dout_25_port, dout_24_port, dout_23_port, dout_22_port, 
      dout_21_port, dout_20_port, dout_19_port, dout_18_port, dout_17_port, 
      dout_16_port, dout_15_port, dout_14_port, dout_13_port, dout_12_port, 
      dout_11_port, dout_10_port, dout_9_port, dout_8_port, dout_7_port, 
      dout_6_port, dout_5_port, dout_4_port, dout_3_port, dout_2_port, 
      dout_1_port, dout_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, net108969, net108970, net108971, 
      net108972, net108973, net108974, net108975, net108976, net108977, 
      net108978, net108979, net108980, net108981, net108982, net108983, 
      net108984, net108985, net108986, net108987, net108988, net108989, 
      net108990, net108991, net108992, net108993, net108994, net108995, 
      net108996, net108997, net108998, net108999, net109000 : std_logic;

begin
   dout <= ( dout_31_port, dout_30_port, dout_29_port, dout_28_port, 
      dout_27_port, dout_26_port, dout_25_port, dout_24_port, dout_23_port, 
      dout_22_port, dout_21_port, dout_20_port, dout_19_port, dout_18_port, 
      dout_17_port, dout_16_port, dout_15_port, dout_14_port, dout_13_port, 
      dout_12_port, dout_11_port, dout_10_port, dout_9_port, dout_8_port, 
      dout_7_port, dout_6_port, dout_5_port, dout_4_port, dout_3_port, 
      dout_2_port, dout_1_port, dout_0_port );
   
   dout_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           dout_31_port, QN => net109000);
   dout_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           dout_30_port, QN => net108999);
   dout_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           dout_29_port, QN => net108998);
   dout_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           dout_28_port, QN => net108997);
   dout_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           dout_27_port, QN => net108996);
   dout_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => rst, Q => 
                           dout_26_port, QN => net108995);
   dout_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => rst, Q => 
                           dout_25_port, QN => net108994);
   dout_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => rst, Q => 
                           dout_24_port, QN => net108993);
   dout_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => rst, Q => 
                           dout_23_port, QN => net108992);
   dout_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => rst, Q => 
                           dout_22_port, QN => net108991);
   dout_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => rst, Q => 
                           dout_21_port, QN => net108990);
   dout_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => rst, Q => 
                           dout_20_port, QN => net108989);
   dout_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => rst, Q => 
                           dout_19_port, QN => net108988);
   dout_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => rst, Q => 
                           dout_18_port, QN => net108987);
   dout_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => rst, Q => 
                           dout_17_port, QN => net108986);
   dout_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => rst, Q => 
                           dout_16_port, QN => net108985);
   dout_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => rst, Q => 
                           dout_15_port, QN => net108984);
   dout_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => rst, Q => 
                           dout_14_port, QN => net108983);
   dout_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => rst, Q => 
                           dout_13_port, QN => net108982);
   dout_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => rst, Q => 
                           dout_12_port, QN => net108981);
   dout_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => rst, Q => 
                           dout_11_port, QN => net108980);
   dout_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => rst, Q => 
                           dout_10_port, QN => net108979);
   dout_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => rst, Q => 
                           dout_9_port, QN => net108978);
   dout_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => rst, Q => 
                           dout_8_port, QN => net108977);
   dout_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => rst, Q => 
                           dout_7_port, QN => net108976);
   dout_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => rst, Q => 
                           dout_6_port, QN => net108975);
   dout_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => rst, Q => 
                           dout_5_port, QN => net108974);
   dout_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => rst, Q => 
                           dout_4_port, QN => net108973);
   dout_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => rst, Q => 
                           dout_3_port, QN => net108972);
   dout_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => rst, Q => 
                           dout_2_port, QN => net108971);
   dout_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => rst, Q => 
                           dout_1_port, QN => net108970);
   dout_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => rst, Q => 
                           dout_0_port, QN => net108969);
   U2 : MUX2_X1 port map( A => dout_31_port, B => din(31), S => en, Z => n1);
   U3 : MUX2_X1 port map( A => dout_30_port, B => din(30), S => en, Z => n2);
   U4 : MUX2_X1 port map( A => dout_29_port, B => din(29), S => en, Z => n3);
   U5 : MUX2_X1 port map( A => dout_28_port, B => din(28), S => en, Z => n4);
   U6 : MUX2_X1 port map( A => dout_27_port, B => din(27), S => en, Z => n5);
   U7 : MUX2_X1 port map( A => dout_26_port, B => din(26), S => en, Z => n6);
   U8 : MUX2_X1 port map( A => dout_25_port, B => din(25), S => en, Z => n7);
   U9 : MUX2_X1 port map( A => dout_24_port, B => din(24), S => en, Z => n8);
   U10 : MUX2_X1 port map( A => dout_23_port, B => din(23), S => en, Z => n9);
   U11 : MUX2_X1 port map( A => dout_22_port, B => din(22), S => en, Z => n10);
   U12 : MUX2_X1 port map( A => dout_21_port, B => din(21), S => en, Z => n11);
   U13 : MUX2_X1 port map( A => dout_20_port, B => din(20), S => en, Z => n12);
   U14 : MUX2_X1 port map( A => dout_19_port, B => din(19), S => en, Z => n13);
   U15 : MUX2_X1 port map( A => dout_18_port, B => din(18), S => en, Z => n14);
   U16 : MUX2_X1 port map( A => dout_17_port, B => din(17), S => en, Z => n15);
   U17 : MUX2_X1 port map( A => dout_16_port, B => din(16), S => en, Z => n16);
   U18 : MUX2_X1 port map( A => dout_15_port, B => din(15), S => en, Z => n17);
   U19 : MUX2_X1 port map( A => dout_14_port, B => din(14), S => en, Z => n18);
   U20 : MUX2_X1 port map( A => dout_13_port, B => din(13), S => en, Z => n19);
   U21 : MUX2_X1 port map( A => dout_12_port, B => din(12), S => en, Z => n20);
   U22 : MUX2_X1 port map( A => dout_11_port, B => din(11), S => en, Z => n21);
   U23 : MUX2_X1 port map( A => dout_10_port, B => din(10), S => en, Z => n22);
   U24 : MUX2_X1 port map( A => dout_9_port, B => din(9), S => en, Z => n23);
   U25 : MUX2_X1 port map( A => dout_8_port, B => din(8), S => en, Z => n24);
   U26 : MUX2_X1 port map( A => dout_7_port, B => din(7), S => en, Z => n25);
   U27 : MUX2_X1 port map( A => dout_6_port, B => din(6), S => en, Z => n26);
   U28 : MUX2_X1 port map( A => dout_5_port, B => din(5), S => en, Z => n27);
   U29 : MUX2_X1 port map( A => dout_4_port, B => din(4), S => en, Z => n28);
   U30 : MUX2_X1 port map( A => dout_3_port, B => din(3), S => en, Z => n29);
   U31 : MUX2_X1 port map( A => dout_2_port, B => din(2), S => en, Z => n30);
   U32 : MUX2_X1 port map( A => dout_1_port, B => din(1), S => en, Z => n31);
   U33 : MUX2_X1 port map( A => dout_0_port, B => din(0), S => en, Z => n32);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE32_5 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 0);
         dout : out std_logic_vector (31 downto 0));

end Reg_DATA_SIZE32_5;

architecture SYN_reg_arch of Reg_DATA_SIZE32_5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal dout_31_port, dout_30_port, dout_29_port, dout_28_port, dout_27_port,
      dout_26_port, dout_25_port, dout_24_port, dout_23_port, dout_22_port, 
      dout_21_port, dout_20_port, dout_19_port, dout_18_port, dout_17_port, 
      dout_16_port, dout_15_port, dout_14_port, dout_13_port, dout_12_port, 
      dout_11_port, dout_10_port, dout_9_port, dout_8_port, dout_7_port, 
      dout_6_port, dout_5_port, dout_4_port, dout_3_port, dout_2_port, 
      dout_1_port, dout_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, net108937, net108938, net108939, 
      net108940, net108941, net108942, net108943, net108944, net108945, 
      net108946, net108947, net108948, net108949, net108950, net108951, 
      net108952, net108953, net108954, net108955, net108956, net108957, 
      net108958, net108959, net108960, net108961, net108962, net108963, 
      net108964, net108965, net108966, net108967, net108968 : std_logic;

begin
   dout <= ( dout_31_port, dout_30_port, dout_29_port, dout_28_port, 
      dout_27_port, dout_26_port, dout_25_port, dout_24_port, dout_23_port, 
      dout_22_port, dout_21_port, dout_20_port, dout_19_port, dout_18_port, 
      dout_17_port, dout_16_port, dout_15_port, dout_14_port, dout_13_port, 
      dout_12_port, dout_11_port, dout_10_port, dout_9_port, dout_8_port, 
      dout_7_port, dout_6_port, dout_5_port, dout_4_port, dout_3_port, 
      dout_2_port, dout_1_port, dout_0_port );
   
   dout_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           dout_31_port, QN => net108968);
   dout_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           dout_30_port, QN => net108967);
   dout_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           dout_29_port, QN => net108966);
   dout_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           dout_28_port, QN => net108965);
   dout_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           dout_27_port, QN => net108964);
   dout_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => rst, Q => 
                           dout_26_port, QN => net108963);
   dout_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => rst, Q => 
                           dout_25_port, QN => net108962);
   dout_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => rst, Q => 
                           dout_24_port, QN => net108961);
   dout_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => rst, Q => 
                           dout_23_port, QN => net108960);
   dout_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => rst, Q => 
                           dout_22_port, QN => net108959);
   dout_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => rst, Q => 
                           dout_21_port, QN => net108958);
   dout_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => rst, Q => 
                           dout_20_port, QN => net108957);
   dout_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => rst, Q => 
                           dout_19_port, QN => net108956);
   dout_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => rst, Q => 
                           dout_18_port, QN => net108955);
   dout_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => rst, Q => 
                           dout_17_port, QN => net108954);
   dout_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => rst, Q => 
                           dout_16_port, QN => net108953);
   dout_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => rst, Q => 
                           dout_15_port, QN => net108952);
   dout_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => rst, Q => 
                           dout_14_port, QN => net108951);
   dout_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => rst, Q => 
                           dout_13_port, QN => net108950);
   dout_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => rst, Q => 
                           dout_12_port, QN => net108949);
   dout_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => rst, Q => 
                           dout_11_port, QN => net108948);
   dout_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => rst, Q => 
                           dout_10_port, QN => net108947);
   dout_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => rst, Q => 
                           dout_9_port, QN => net108946);
   dout_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => rst, Q => 
                           dout_8_port, QN => net108945);
   dout_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => rst, Q => 
                           dout_7_port, QN => net108944);
   dout_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => rst, Q => 
                           dout_6_port, QN => net108943);
   dout_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => rst, Q => 
                           dout_5_port, QN => net108942);
   dout_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => rst, Q => 
                           dout_4_port, QN => net108941);
   dout_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => rst, Q => 
                           dout_3_port, QN => net108940);
   dout_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => rst, Q => 
                           dout_2_port, QN => net108939);
   dout_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => rst, Q => 
                           dout_1_port, QN => net108938);
   dout_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => rst, Q => 
                           dout_0_port, QN => net108937);
   U2 : MUX2_X1 port map( A => dout_31_port, B => din(31), S => en, Z => n1);
   U3 : MUX2_X1 port map( A => dout_30_port, B => din(30), S => en, Z => n2);
   U4 : MUX2_X1 port map( A => dout_29_port, B => din(29), S => en, Z => n3);
   U5 : MUX2_X1 port map( A => dout_28_port, B => din(28), S => en, Z => n4);
   U6 : MUX2_X1 port map( A => dout_27_port, B => din(27), S => en, Z => n5);
   U7 : MUX2_X1 port map( A => dout_26_port, B => din(26), S => en, Z => n6);
   U8 : MUX2_X1 port map( A => dout_25_port, B => din(25), S => en, Z => n7);
   U9 : MUX2_X1 port map( A => dout_24_port, B => din(24), S => en, Z => n8);
   U10 : MUX2_X1 port map( A => dout_23_port, B => din(23), S => en, Z => n9);
   U11 : MUX2_X1 port map( A => dout_22_port, B => din(22), S => en, Z => n10);
   U12 : MUX2_X1 port map( A => dout_21_port, B => din(21), S => en, Z => n11);
   U13 : MUX2_X1 port map( A => dout_20_port, B => din(20), S => en, Z => n12);
   U14 : MUX2_X1 port map( A => dout_19_port, B => din(19), S => en, Z => n13);
   U15 : MUX2_X1 port map( A => dout_18_port, B => din(18), S => en, Z => n14);
   U16 : MUX2_X1 port map( A => dout_17_port, B => din(17), S => en, Z => n15);
   U17 : MUX2_X1 port map( A => dout_16_port, B => din(16), S => en, Z => n16);
   U18 : MUX2_X1 port map( A => dout_15_port, B => din(15), S => en, Z => n17);
   U19 : MUX2_X1 port map( A => dout_14_port, B => din(14), S => en, Z => n18);
   U20 : MUX2_X1 port map( A => dout_13_port, B => din(13), S => en, Z => n19);
   U21 : MUX2_X1 port map( A => dout_12_port, B => din(12), S => en, Z => n20);
   U22 : MUX2_X1 port map( A => dout_11_port, B => din(11), S => en, Z => n21);
   U23 : MUX2_X1 port map( A => dout_10_port, B => din(10), S => en, Z => n22);
   U24 : MUX2_X1 port map( A => dout_9_port, B => din(9), S => en, Z => n23);
   U25 : MUX2_X1 port map( A => dout_8_port, B => din(8), S => en, Z => n24);
   U26 : MUX2_X1 port map( A => dout_7_port, B => din(7), S => en, Z => n25);
   U27 : MUX2_X1 port map( A => dout_6_port, B => din(6), S => en, Z => n26);
   U28 : MUX2_X1 port map( A => dout_5_port, B => din(5), S => en, Z => n27);
   U29 : MUX2_X1 port map( A => dout_4_port, B => din(4), S => en, Z => n28);
   U30 : MUX2_X1 port map( A => dout_3_port, B => din(3), S => en, Z => n29);
   U31 : MUX2_X1 port map( A => dout_2_port, B => din(2), S => en, Z => n30);
   U32 : MUX2_X1 port map( A => dout_1_port, B => din(1), S => en, Z => n31);
   U33 : MUX2_X1 port map( A => dout_0_port, B => din(0), S => en, Z => n32);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE32_4 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 0);
         dout : out std_logic_vector (31 downto 0));

end Reg_DATA_SIZE32_4;

architecture SYN_reg_arch of Reg_DATA_SIZE32_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal dout_31_port, dout_30_port, dout_29_port, dout_28_port, dout_27_port,
      dout_26_port, dout_25_port, dout_24_port, dout_23_port, dout_22_port, 
      dout_21_port, dout_20_port, dout_19_port, dout_18_port, dout_17_port, 
      dout_16_port, dout_15_port, dout_14_port, dout_13_port, dout_12_port, 
      dout_11_port, dout_10_port, dout_9_port, dout_8_port, dout_7_port, 
      dout_6_port, dout_5_port, dout_4_port, dout_3_port, dout_2_port, 
      dout_1_port, dout_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, net108905, net108906, net108907, 
      net108908, net108909, net108910, net108911, net108912, net108913, 
      net108914, net108915, net108916, net108917, net108918, net108919, 
      net108920, net108921, net108922, net108923, net108924, net108925, 
      net108926, net108927, net108928, net108929, net108930, net108931, 
      net108932, net108933, net108934, net108935, net108936 : std_logic;

begin
   dout <= ( dout_31_port, dout_30_port, dout_29_port, dout_28_port, 
      dout_27_port, dout_26_port, dout_25_port, dout_24_port, dout_23_port, 
      dout_22_port, dout_21_port, dout_20_port, dout_19_port, dout_18_port, 
      dout_17_port, dout_16_port, dout_15_port, dout_14_port, dout_13_port, 
      dout_12_port, dout_11_port, dout_10_port, dout_9_port, dout_8_port, 
      dout_7_port, dout_6_port, dout_5_port, dout_4_port, dout_3_port, 
      dout_2_port, dout_1_port, dout_0_port );
   
   dout_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           dout_31_port, QN => net108936);
   dout_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           dout_30_port, QN => net108935);
   dout_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           dout_29_port, QN => net108934);
   dout_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           dout_28_port, QN => net108933);
   dout_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           dout_27_port, QN => net108932);
   dout_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => rst, Q => 
                           dout_26_port, QN => net108931);
   dout_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => rst, Q => 
                           dout_25_port, QN => net108930);
   dout_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => rst, Q => 
                           dout_24_port, QN => net108929);
   dout_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => rst, Q => 
                           dout_23_port, QN => net108928);
   dout_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => rst, Q => 
                           dout_22_port, QN => net108927);
   dout_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => rst, Q => 
                           dout_21_port, QN => net108926);
   dout_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => rst, Q => 
                           dout_20_port, QN => net108925);
   dout_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => rst, Q => 
                           dout_19_port, QN => net108924);
   dout_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => rst, Q => 
                           dout_18_port, QN => net108923);
   dout_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => rst, Q => 
                           dout_17_port, QN => net108922);
   dout_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => rst, Q => 
                           dout_16_port, QN => net108921);
   dout_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => rst, Q => 
                           dout_15_port, QN => net108920);
   dout_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => rst, Q => 
                           dout_14_port, QN => net108919);
   dout_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => rst, Q => 
                           dout_13_port, QN => net108918);
   dout_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => rst, Q => 
                           dout_12_port, QN => net108917);
   dout_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => rst, Q => 
                           dout_11_port, QN => net108916);
   dout_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => rst, Q => 
                           dout_10_port, QN => net108915);
   dout_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => rst, Q => 
                           dout_9_port, QN => net108914);
   dout_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => rst, Q => 
                           dout_8_port, QN => net108913);
   dout_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => rst, Q => 
                           dout_7_port, QN => net108912);
   dout_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => rst, Q => 
                           dout_6_port, QN => net108911);
   dout_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => rst, Q => 
                           dout_5_port, QN => net108910);
   dout_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => rst, Q => 
                           dout_4_port, QN => net108909);
   dout_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => rst, Q => 
                           dout_3_port, QN => net108908);
   dout_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => rst, Q => 
                           dout_2_port, QN => net108907);
   dout_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => rst, Q => 
                           dout_1_port, QN => net108906);
   dout_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => rst, Q => 
                           dout_0_port, QN => net108905);
   U2 : MUX2_X1 port map( A => dout_31_port, B => din(31), S => en, Z => n1);
   U3 : MUX2_X1 port map( A => dout_30_port, B => din(30), S => en, Z => n2);
   U4 : MUX2_X1 port map( A => dout_29_port, B => din(29), S => en, Z => n3);
   U5 : MUX2_X1 port map( A => dout_28_port, B => din(28), S => en, Z => n4);
   U6 : MUX2_X1 port map( A => dout_27_port, B => din(27), S => en, Z => n5);
   U7 : MUX2_X1 port map( A => dout_26_port, B => din(26), S => en, Z => n6);
   U8 : MUX2_X1 port map( A => dout_25_port, B => din(25), S => en, Z => n7);
   U9 : MUX2_X1 port map( A => dout_24_port, B => din(24), S => en, Z => n8);
   U10 : MUX2_X1 port map( A => dout_23_port, B => din(23), S => en, Z => n9);
   U11 : MUX2_X1 port map( A => dout_22_port, B => din(22), S => en, Z => n10);
   U12 : MUX2_X1 port map( A => dout_21_port, B => din(21), S => en, Z => n11);
   U13 : MUX2_X1 port map( A => dout_20_port, B => din(20), S => en, Z => n12);
   U14 : MUX2_X1 port map( A => dout_19_port, B => din(19), S => en, Z => n13);
   U15 : MUX2_X1 port map( A => dout_18_port, B => din(18), S => en, Z => n14);
   U16 : MUX2_X1 port map( A => dout_17_port, B => din(17), S => en, Z => n15);
   U17 : MUX2_X1 port map( A => dout_16_port, B => din(16), S => en, Z => n16);
   U18 : MUX2_X1 port map( A => dout_15_port, B => din(15), S => en, Z => n17);
   U19 : MUX2_X1 port map( A => dout_14_port, B => din(14), S => en, Z => n18);
   U20 : MUX2_X1 port map( A => dout_13_port, B => din(13), S => en, Z => n19);
   U21 : MUX2_X1 port map( A => dout_12_port, B => din(12), S => en, Z => n20);
   U22 : MUX2_X1 port map( A => dout_11_port, B => din(11), S => en, Z => n21);
   U23 : MUX2_X1 port map( A => dout_10_port, B => din(10), S => en, Z => n22);
   U24 : MUX2_X1 port map( A => dout_9_port, B => din(9), S => en, Z => n23);
   U25 : MUX2_X1 port map( A => dout_8_port, B => din(8), S => en, Z => n24);
   U26 : MUX2_X1 port map( A => dout_7_port, B => din(7), S => en, Z => n25);
   U27 : MUX2_X1 port map( A => dout_6_port, B => din(6), S => en, Z => n26);
   U28 : MUX2_X1 port map( A => dout_5_port, B => din(5), S => en, Z => n27);
   U29 : MUX2_X1 port map( A => dout_4_port, B => din(4), S => en, Z => n28);
   U30 : MUX2_X1 port map( A => dout_3_port, B => din(3), S => en, Z => n29);
   U31 : MUX2_X1 port map( A => dout_2_port, B => din(2), S => en, Z => n30);
   U32 : MUX2_X1 port map( A => dout_1_port, B => din(1), S => en, Z => n31);
   U33 : MUX2_X1 port map( A => dout_0_port, B => din(0), S => en, Z => n32);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE32_3 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 0);
         dout : out std_logic_vector (31 downto 0));

end Reg_DATA_SIZE32_3;

architecture SYN_reg_arch of Reg_DATA_SIZE32_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal dout_31_port, dout_30_port, dout_29_port, dout_28_port, dout_27_port,
      dout_26_port, dout_25_port, dout_24_port, dout_23_port, dout_22_port, 
      dout_21_port, dout_20_port, dout_19_port, dout_18_port, dout_17_port, 
      dout_16_port, dout_15_port, dout_14_port, dout_13_port, dout_12_port, 
      dout_11_port, dout_10_port, dout_9_port, dout_8_port, dout_7_port, 
      dout_6_port, dout_5_port, dout_4_port, dout_3_port, dout_2_port, 
      dout_1_port, dout_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, 
      n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55
      , n56, n57, n58, n59, n60, n61, n62, n63, n64 : std_logic;

begin
   dout <= ( dout_31_port, dout_30_port, dout_29_port, dout_28_port, 
      dout_27_port, dout_26_port, dout_25_port, dout_24_port, dout_23_port, 
      dout_22_port, dout_21_port, dout_20_port, dout_19_port, dout_18_port, 
      dout_17_port, dout_16_port, dout_15_port, dout_14_port, dout_13_port, 
      dout_12_port, dout_11_port, dout_10_port, dout_9_port, dout_8_port, 
      dout_7_port, dout_6_port, dout_5_port, dout_4_port, dout_3_port, 
      dout_2_port, dout_1_port, dout_0_port );
   
   dout_reg_0_inst : DFFR_X2 port map( D => n64, CK => clk, RN => rst, Q => 
                           dout_0_port, QN => n32);
   dout_reg_1_inst : DFFR_X2 port map( D => n63, CK => clk, RN => rst, Q => 
                           dout_1_port, QN => n31);
   dout_reg_2_inst : DFFR_X2 port map( D => n62, CK => clk, RN => rst, Q => 
                           dout_2_port, QN => n30);
   dout_reg_3_inst : DFFR_X2 port map( D => n61, CK => clk, RN => rst, Q => 
                           dout_3_port, QN => n29);
   dout_reg_4_inst : DFFR_X2 port map( D => n60, CK => clk, RN => rst, Q => 
                           dout_4_port, QN => n28);
   dout_reg_5_inst : DFFR_X2 port map( D => n59, CK => clk, RN => rst, Q => 
                           dout_5_port, QN => n27);
   dout_reg_6_inst : DFFR_X2 port map( D => n58, CK => clk, RN => rst, Q => 
                           dout_6_port, QN => n26);
   dout_reg_7_inst : DFFR_X2 port map( D => n57, CK => clk, RN => rst, Q => 
                           dout_7_port, QN => n25);
   dout_reg_8_inst : DFFR_X2 port map( D => n56, CK => clk, RN => rst, Q => 
                           dout_8_port, QN => n24);
   dout_reg_9_inst : DFFR_X2 port map( D => n55, CK => clk, RN => rst, Q => 
                           dout_9_port, QN => n23);
   dout_reg_10_inst : DFFR_X2 port map( D => n54, CK => clk, RN => rst, Q => 
                           dout_10_port, QN => n22);
   dout_reg_11_inst : DFFR_X2 port map( D => n53, CK => clk, RN => rst, Q => 
                           dout_11_port, QN => n21);
   dout_reg_12_inst : DFFR_X2 port map( D => n52, CK => clk, RN => rst, Q => 
                           dout_12_port, QN => n20);
   dout_reg_13_inst : DFFR_X2 port map( D => n51, CK => clk, RN => rst, Q => 
                           dout_13_port, QN => n19);
   dout_reg_14_inst : DFFR_X2 port map( D => n50, CK => clk, RN => rst, Q => 
                           dout_14_port, QN => n18);
   dout_reg_15_inst : DFFR_X2 port map( D => n49, CK => clk, RN => rst, Q => 
                           dout_15_port, QN => n17);
   dout_reg_16_inst : DFFR_X2 port map( D => n48, CK => clk, RN => rst, Q => 
                           dout_16_port, QN => n16);
   dout_reg_17_inst : DFFR_X2 port map( D => n47, CK => clk, RN => rst, Q => 
                           dout_17_port, QN => n15);
   dout_reg_18_inst : DFFR_X2 port map( D => n46, CK => clk, RN => rst, Q => 
                           dout_18_port, QN => n14);
   dout_reg_19_inst : DFFR_X2 port map( D => n45, CK => clk, RN => rst, Q => 
                           dout_19_port, QN => n13);
   dout_reg_20_inst : DFFR_X2 port map( D => n44, CK => clk, RN => rst, Q => 
                           dout_20_port, QN => n12);
   dout_reg_21_inst : DFFR_X2 port map( D => n43, CK => clk, RN => rst, Q => 
                           dout_21_port, QN => n11);
   dout_reg_22_inst : DFFR_X2 port map( D => n42, CK => clk, RN => rst, Q => 
                           dout_22_port, QN => n10);
   dout_reg_23_inst : DFFR_X2 port map( D => n41, CK => clk, RN => rst, Q => 
                           dout_23_port, QN => n9);
   dout_reg_24_inst : DFFR_X2 port map( D => n40, CK => clk, RN => rst, Q => 
                           dout_24_port, QN => n8);
   dout_reg_25_inst : DFFR_X2 port map( D => n39, CK => clk, RN => rst, Q => 
                           dout_25_port, QN => n7);
   dout_reg_26_inst : DFFR_X2 port map( D => n38, CK => clk, RN => rst, Q => 
                           dout_26_port, QN => n6);
   dout_reg_27_inst : DFFR_X2 port map( D => n37, CK => clk, RN => rst, Q => 
                           dout_27_port, QN => n5);
   dout_reg_28_inst : DFFR_X2 port map( D => n36, CK => clk, RN => rst, Q => 
                           dout_28_port, QN => n4);
   dout_reg_29_inst : DFFR_X2 port map( D => n35, CK => clk, RN => rst, Q => 
                           dout_29_port, QN => n3);
   dout_reg_30_inst : DFFR_X2 port map( D => n34, CK => clk, RN => rst, Q => 
                           dout_30_port, QN => n2);
   dout_reg_31_inst : DFFR_X2 port map( D => n33, CK => clk, RN => rst, Q => 
                           dout_31_port, QN => n1);
   U2 : MUX2_X1 port map( A => dout_31_port, B => din(31), S => en, Z => n33);
   U3 : MUX2_X1 port map( A => dout_30_port, B => din(30), S => en, Z => n34);
   U4 : MUX2_X1 port map( A => dout_29_port, B => din(29), S => en, Z => n35);
   U5 : MUX2_X1 port map( A => dout_28_port, B => din(28), S => en, Z => n36);
   U6 : MUX2_X1 port map( A => dout_27_port, B => din(27), S => en, Z => n37);
   U7 : MUX2_X1 port map( A => dout_26_port, B => din(26), S => en, Z => n38);
   U8 : MUX2_X1 port map( A => dout_25_port, B => din(25), S => en, Z => n39);
   U9 : MUX2_X1 port map( A => dout_24_port, B => din(24), S => en, Z => n40);
   U10 : MUX2_X1 port map( A => dout_23_port, B => din(23), S => en, Z => n41);
   U11 : MUX2_X1 port map( A => dout_22_port, B => din(22), S => en, Z => n42);
   U12 : MUX2_X1 port map( A => dout_21_port, B => din(21), S => en, Z => n43);
   U13 : MUX2_X1 port map( A => dout_20_port, B => din(20), S => en, Z => n44);
   U14 : MUX2_X1 port map( A => dout_19_port, B => din(19), S => en, Z => n45);
   U15 : MUX2_X1 port map( A => dout_18_port, B => din(18), S => en, Z => n46);
   U16 : MUX2_X1 port map( A => dout_17_port, B => din(17), S => en, Z => n47);
   U17 : MUX2_X1 port map( A => dout_16_port, B => din(16), S => en, Z => n48);
   U18 : MUX2_X1 port map( A => dout_15_port, B => din(15), S => en, Z => n49);
   U19 : MUX2_X1 port map( A => dout_14_port, B => din(14), S => en, Z => n50);
   U20 : MUX2_X1 port map( A => dout_13_port, B => din(13), S => en, Z => n51);
   U21 : MUX2_X1 port map( A => dout_12_port, B => din(12), S => en, Z => n52);
   U22 : MUX2_X1 port map( A => dout_11_port, B => din(11), S => en, Z => n53);
   U23 : MUX2_X1 port map( A => dout_10_port, B => din(10), S => en, Z => n54);
   U24 : MUX2_X1 port map( A => dout_9_port, B => din(9), S => en, Z => n55);
   U25 : MUX2_X1 port map( A => dout_8_port, B => din(8), S => en, Z => n56);
   U26 : MUX2_X1 port map( A => dout_7_port, B => din(7), S => en, Z => n57);
   U27 : MUX2_X1 port map( A => dout_6_port, B => din(6), S => en, Z => n58);
   U28 : MUX2_X1 port map( A => dout_5_port, B => din(5), S => en, Z => n59);
   U29 : MUX2_X1 port map( A => dout_4_port, B => din(4), S => en, Z => n60);
   U30 : MUX2_X1 port map( A => dout_3_port, B => din(3), S => en, Z => n61);
   U31 : MUX2_X1 port map( A => dout_2_port, B => din(2), S => en, Z => n62);
   U32 : MUX2_X1 port map( A => dout_1_port, B => din(1), S => en, Z => n63);
   U33 : MUX2_X1 port map( A => dout_0_port, B => din(0), S => en, Z => n64);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE32_2 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 0);
         dout : out std_logic_vector (31 downto 0));

end Reg_DATA_SIZE32_2;

architecture SYN_reg_arch of Reg_DATA_SIZE32_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal dout_31_port, dout_30_port, dout_29_port, dout_28_port, dout_27_port,
      dout_26_port, dout_25_port, dout_24_port, dout_23_port, dout_22_port, 
      dout_21_port, dout_20_port, dout_19_port, dout_18_port, dout_17_port, 
      dout_16_port, dout_15_port, dout_14_port, dout_13_port, dout_12_port, 
      dout_11_port, dout_10_port, dout_9_port, dout_8_port, dout_7_port, 
      dout_6_port, dout_5_port, dout_4_port, dout_3_port, dout_2_port, 
      dout_1_port, dout_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, net108873, net108874, net108875, 
      net108876, net108877, net108878, net108879, net108880, net108881, 
      net108882, net108883, net108884, net108885, net108886, net108887, 
      net108888, net108889, net108890, net108891, net108892, net108893, 
      net108894, net108895, net108896, net108897, net108898, net108899, 
      net108900, net108901, net108902, net108903, net108904 : std_logic;

begin
   dout <= ( dout_31_port, dout_30_port, dout_29_port, dout_28_port, 
      dout_27_port, dout_26_port, dout_25_port, dout_24_port, dout_23_port, 
      dout_22_port, dout_21_port, dout_20_port, dout_19_port, dout_18_port, 
      dout_17_port, dout_16_port, dout_15_port, dout_14_port, dout_13_port, 
      dout_12_port, dout_11_port, dout_10_port, dout_9_port, dout_8_port, 
      dout_7_port, dout_6_port, dout_5_port, dout_4_port, dout_3_port, 
      dout_2_port, dout_1_port, dout_0_port );
   
   dout_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           dout_31_port, QN => net108904);
   dout_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           dout_30_port, QN => net108903);
   dout_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           dout_29_port, QN => net108902);
   dout_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           dout_28_port, QN => net108901);
   dout_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           dout_27_port, QN => net108900);
   dout_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => rst, Q => 
                           dout_26_port, QN => net108899);
   dout_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => rst, Q => 
                           dout_25_port, QN => net108898);
   dout_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => rst, Q => 
                           dout_24_port, QN => net108897);
   dout_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => rst, Q => 
                           dout_23_port, QN => net108896);
   dout_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => rst, Q => 
                           dout_22_port, QN => net108895);
   dout_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => rst, Q => 
                           dout_21_port, QN => net108894);
   dout_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => rst, Q => 
                           dout_20_port, QN => net108893);
   dout_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => rst, Q => 
                           dout_19_port, QN => net108892);
   dout_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => rst, Q => 
                           dout_18_port, QN => net108891);
   dout_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => rst, Q => 
                           dout_17_port, QN => net108890);
   dout_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => rst, Q => 
                           dout_16_port, QN => net108889);
   dout_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => rst, Q => 
                           dout_15_port, QN => net108888);
   dout_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => rst, Q => 
                           dout_14_port, QN => net108887);
   dout_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => rst, Q => 
                           dout_13_port, QN => net108886);
   dout_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => rst, Q => 
                           dout_12_port, QN => net108885);
   dout_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => rst, Q => 
                           dout_11_port, QN => net108884);
   dout_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => rst, Q => 
                           dout_10_port, QN => net108883);
   dout_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => rst, Q => 
                           dout_9_port, QN => net108882);
   dout_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => rst, Q => 
                           dout_8_port, QN => net108881);
   dout_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => rst, Q => 
                           dout_7_port, QN => net108880);
   dout_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => rst, Q => 
                           dout_6_port, QN => net108879);
   dout_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => rst, Q => 
                           dout_5_port, QN => net108878);
   dout_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => rst, Q => 
                           dout_4_port, QN => net108877);
   dout_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => rst, Q => 
                           dout_3_port, QN => net108876);
   dout_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => rst, Q => 
                           dout_2_port, QN => net108875);
   dout_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => rst, Q => 
                           dout_1_port, QN => net108874);
   dout_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => rst, Q => 
                           dout_0_port, QN => net108873);
   U2 : MUX2_X1 port map( A => dout_31_port, B => din(31), S => en, Z => n1);
   U3 : MUX2_X1 port map( A => dout_30_port, B => din(30), S => en, Z => n2);
   U4 : MUX2_X1 port map( A => dout_29_port, B => din(29), S => en, Z => n3);
   U5 : MUX2_X1 port map( A => dout_28_port, B => din(28), S => en, Z => n4);
   U6 : MUX2_X1 port map( A => dout_27_port, B => din(27), S => en, Z => n5);
   U7 : MUX2_X1 port map( A => dout_26_port, B => din(26), S => en, Z => n6);
   U8 : MUX2_X1 port map( A => dout_25_port, B => din(25), S => en, Z => n7);
   U9 : MUX2_X1 port map( A => dout_24_port, B => din(24), S => en, Z => n8);
   U10 : MUX2_X1 port map( A => dout_23_port, B => din(23), S => en, Z => n9);
   U11 : MUX2_X1 port map( A => dout_22_port, B => din(22), S => en, Z => n10);
   U12 : MUX2_X1 port map( A => dout_21_port, B => din(21), S => en, Z => n11);
   U13 : MUX2_X1 port map( A => dout_20_port, B => din(20), S => en, Z => n12);
   U14 : MUX2_X1 port map( A => dout_19_port, B => din(19), S => en, Z => n13);
   U15 : MUX2_X1 port map( A => dout_18_port, B => din(18), S => en, Z => n14);
   U16 : MUX2_X1 port map( A => dout_17_port, B => din(17), S => en, Z => n15);
   U17 : MUX2_X1 port map( A => dout_16_port, B => din(16), S => en, Z => n16);
   U18 : MUX2_X1 port map( A => dout_15_port, B => din(15), S => en, Z => n17);
   U19 : MUX2_X1 port map( A => dout_14_port, B => din(14), S => en, Z => n18);
   U20 : MUX2_X1 port map( A => dout_13_port, B => din(13), S => en, Z => n19);
   U21 : MUX2_X1 port map( A => dout_12_port, B => din(12), S => en, Z => n20);
   U22 : MUX2_X1 port map( A => dout_11_port, B => din(11), S => en, Z => n21);
   U23 : MUX2_X1 port map( A => dout_10_port, B => din(10), S => en, Z => n22);
   U24 : MUX2_X1 port map( A => dout_9_port, B => din(9), S => en, Z => n23);
   U25 : MUX2_X1 port map( A => dout_8_port, B => din(8), S => en, Z => n24);
   U26 : MUX2_X1 port map( A => dout_7_port, B => din(7), S => en, Z => n25);
   U27 : MUX2_X1 port map( A => dout_6_port, B => din(6), S => en, Z => n26);
   U28 : MUX2_X1 port map( A => dout_5_port, B => din(5), S => en, Z => n27);
   U29 : MUX2_X1 port map( A => dout_4_port, B => din(4), S => en, Z => n28);
   U30 : MUX2_X1 port map( A => dout_3_port, B => din(3), S => en, Z => n29);
   U31 : MUX2_X1 port map( A => dout_2_port, B => din(2), S => en, Z => n30);
   U32 : MUX2_X1 port map( A => dout_1_port, B => din(1), S => en, Z => n31);
   U33 : MUX2_X1 port map( A => dout_0_port, B => din(0), S => en, Z => n32);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE32_1 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 0);
         dout : out std_logic_vector (31 downto 0));

end Reg_DATA_SIZE32_1;

architecture SYN_reg_arch of Reg_DATA_SIZE32_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal dout_31_port, dout_30_port, dout_29_port, dout_28_port, dout_27_port,
      dout_26_port, dout_25_port, dout_24_port, dout_23_port, dout_22_port, 
      dout_21_port, dout_20_port, dout_19_port, dout_18_port, dout_17_port, 
      dout_16_port, dout_15_port, dout_14_port, dout_13_port, dout_12_port, 
      dout_11_port, dout_10_port, dout_9_port, dout_8_port, dout_7_port, 
      dout_6_port, dout_5_port, dout_4_port, dout_3_port, dout_2_port, 
      dout_1_port, dout_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, 
      n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, net108841, net108842, net108843, 
      net108844, net108845, net108846, net108847, net108848, net108849, 
      net108850, net108851, net108852, net108853, net108854, net108855, 
      net108856, net108857, net108858, net108859, net108860, net108861, 
      net108862, net108863, net108864, net108865, net108866, net108867, 
      net108868, net108869, net108870, net108871, net108872 : std_logic;

begin
   dout <= ( dout_31_port, dout_30_port, dout_29_port, dout_28_port, 
      dout_27_port, dout_26_port, dout_25_port, dout_24_port, dout_23_port, 
      dout_22_port, dout_21_port, dout_20_port, dout_19_port, dout_18_port, 
      dout_17_port, dout_16_port, dout_15_port, dout_14_port, dout_13_port, 
      dout_12_port, dout_11_port, dout_10_port, dout_9_port, dout_8_port, 
      dout_7_port, dout_6_port, dout_5_port, dout_4_port, dout_3_port, 
      dout_2_port, dout_1_port, dout_0_port );
   
   dout_reg_31_inst : DFFR_X1 port map( D => n1, CK => clk, RN => rst, Q => 
                           dout_31_port, QN => net108872);
   dout_reg_30_inst : DFFR_X1 port map( D => n2, CK => clk, RN => rst, Q => 
                           dout_30_port, QN => net108871);
   dout_reg_29_inst : DFFR_X1 port map( D => n3, CK => clk, RN => rst, Q => 
                           dout_29_port, QN => net108870);
   dout_reg_28_inst : DFFR_X1 port map( D => n4, CK => clk, RN => rst, Q => 
                           dout_28_port, QN => net108869);
   dout_reg_27_inst : DFFR_X1 port map( D => n5, CK => clk, RN => rst, Q => 
                           dout_27_port, QN => net108868);
   dout_reg_26_inst : DFFR_X1 port map( D => n6, CK => clk, RN => rst, Q => 
                           dout_26_port, QN => net108867);
   dout_reg_25_inst : DFFR_X1 port map( D => n7, CK => clk, RN => rst, Q => 
                           dout_25_port, QN => net108866);
   dout_reg_24_inst : DFFR_X1 port map( D => n8, CK => clk, RN => rst, Q => 
                           dout_24_port, QN => net108865);
   dout_reg_23_inst : DFFR_X1 port map( D => n9, CK => clk, RN => rst, Q => 
                           dout_23_port, QN => net108864);
   dout_reg_22_inst : DFFR_X1 port map( D => n10, CK => clk, RN => rst, Q => 
                           dout_22_port, QN => net108863);
   dout_reg_21_inst : DFFR_X1 port map( D => n11, CK => clk, RN => rst, Q => 
                           dout_21_port, QN => net108862);
   dout_reg_20_inst : DFFR_X1 port map( D => n12, CK => clk, RN => rst, Q => 
                           dout_20_port, QN => net108861);
   dout_reg_19_inst : DFFR_X1 port map( D => n13, CK => clk, RN => rst, Q => 
                           dout_19_port, QN => net108860);
   dout_reg_18_inst : DFFR_X1 port map( D => n14, CK => clk, RN => rst, Q => 
                           dout_18_port, QN => net108859);
   dout_reg_17_inst : DFFR_X1 port map( D => n15, CK => clk, RN => rst, Q => 
                           dout_17_port, QN => net108858);
   dout_reg_16_inst : DFFR_X1 port map( D => n16, CK => clk, RN => rst, Q => 
                           dout_16_port, QN => net108857);
   dout_reg_15_inst : DFFR_X1 port map( D => n17, CK => clk, RN => rst, Q => 
                           dout_15_port, QN => net108856);
   dout_reg_14_inst : DFFR_X1 port map( D => n18, CK => clk, RN => rst, Q => 
                           dout_14_port, QN => net108855);
   dout_reg_13_inst : DFFR_X1 port map( D => n19, CK => clk, RN => rst, Q => 
                           dout_13_port, QN => net108854);
   dout_reg_12_inst : DFFR_X1 port map( D => n20, CK => clk, RN => rst, Q => 
                           dout_12_port, QN => net108853);
   dout_reg_11_inst : DFFR_X1 port map( D => n21, CK => clk, RN => rst, Q => 
                           dout_11_port, QN => net108852);
   dout_reg_10_inst : DFFR_X1 port map( D => n22, CK => clk, RN => rst, Q => 
                           dout_10_port, QN => net108851);
   dout_reg_9_inst : DFFR_X1 port map( D => n23, CK => clk, RN => rst, Q => 
                           dout_9_port, QN => net108850);
   dout_reg_8_inst : DFFR_X1 port map( D => n24, CK => clk, RN => rst, Q => 
                           dout_8_port, QN => net108849);
   dout_reg_7_inst : DFFR_X1 port map( D => n25, CK => clk, RN => rst, Q => 
                           dout_7_port, QN => net108848);
   dout_reg_6_inst : DFFR_X1 port map( D => n26, CK => clk, RN => rst, Q => 
                           dout_6_port, QN => net108847);
   dout_reg_5_inst : DFFR_X1 port map( D => n27, CK => clk, RN => rst, Q => 
                           dout_5_port, QN => net108846);
   dout_reg_4_inst : DFFR_X1 port map( D => n28, CK => clk, RN => rst, Q => 
                           dout_4_port, QN => net108845);
   dout_reg_3_inst : DFFR_X1 port map( D => n29, CK => clk, RN => rst, Q => 
                           dout_3_port, QN => net108844);
   dout_reg_2_inst : DFFR_X1 port map( D => n30, CK => clk, RN => rst, Q => 
                           dout_2_port, QN => net108843);
   dout_reg_1_inst : DFFR_X1 port map( D => n31, CK => clk, RN => rst, Q => 
                           dout_1_port, QN => net108842);
   dout_reg_0_inst : DFFR_X1 port map( D => n32, CK => clk, RN => rst, Q => 
                           dout_0_port, QN => net108841);
   U2 : MUX2_X1 port map( A => dout_31_port, B => din(31), S => en, Z => n1);
   U3 : MUX2_X1 port map( A => dout_30_port, B => din(30), S => en, Z => n2);
   U4 : MUX2_X1 port map( A => dout_29_port, B => din(29), S => en, Z => n3);
   U5 : MUX2_X1 port map( A => dout_28_port, B => din(28), S => en, Z => n4);
   U6 : MUX2_X1 port map( A => dout_27_port, B => din(27), S => en, Z => n5);
   U7 : MUX2_X1 port map( A => dout_26_port, B => din(26), S => en, Z => n6);
   U8 : MUX2_X1 port map( A => dout_25_port, B => din(25), S => en, Z => n7);
   U9 : MUX2_X1 port map( A => dout_24_port, B => din(24), S => en, Z => n8);
   U10 : MUX2_X1 port map( A => dout_23_port, B => din(23), S => en, Z => n9);
   U11 : MUX2_X1 port map( A => dout_22_port, B => din(22), S => en, Z => n10);
   U12 : MUX2_X1 port map( A => dout_21_port, B => din(21), S => en, Z => n11);
   U13 : MUX2_X1 port map( A => dout_20_port, B => din(20), S => en, Z => n12);
   U14 : MUX2_X1 port map( A => dout_19_port, B => din(19), S => en, Z => n13);
   U15 : MUX2_X1 port map( A => dout_18_port, B => din(18), S => en, Z => n14);
   U16 : MUX2_X1 port map( A => dout_17_port, B => din(17), S => en, Z => n15);
   U17 : MUX2_X1 port map( A => dout_16_port, B => din(16), S => en, Z => n16);
   U18 : MUX2_X1 port map( A => dout_15_port, B => din(15), S => en, Z => n17);
   U19 : MUX2_X1 port map( A => dout_14_port, B => din(14), S => en, Z => n18);
   U20 : MUX2_X1 port map( A => dout_13_port, B => din(13), S => en, Z => n19);
   U21 : MUX2_X1 port map( A => dout_12_port, B => din(12), S => en, Z => n20);
   U22 : MUX2_X1 port map( A => dout_11_port, B => din(11), S => en, Z => n21);
   U23 : MUX2_X1 port map( A => dout_10_port, B => din(10), S => en, Z => n22);
   U24 : MUX2_X1 port map( A => dout_9_port, B => din(9), S => en, Z => n23);
   U25 : MUX2_X1 port map( A => dout_8_port, B => din(8), S => en, Z => n24);
   U26 : MUX2_X1 port map( A => dout_7_port, B => din(7), S => en, Z => n25);
   U27 : MUX2_X1 port map( A => dout_6_port, B => din(6), S => en, Z => n26);
   U28 : MUX2_X1 port map( A => dout_5_port, B => din(5), S => en, Z => n27);
   U29 : MUX2_X1 port map( A => dout_4_port, B => din(4), S => en, Z => n28);
   U30 : MUX2_X1 port map( A => dout_3_port, B => din(3), S => en, Z => n29);
   U31 : MUX2_X1 port map( A => dout_2_port, B => din(2), S => en, Z => n30);
   U32 : MUX2_X1 port map( A => dout_1_port, B => din(1), S => en, Z => n31);
   U33 : MUX2_X1 port map( A => dout_0_port, B => din(0), S => en, Z => n32);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE32_9 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0);  
         dout : out std_logic_vector (31 downto 0));

end Mux_DATA_SIZE32_9;

architecture SYN_mux_arch of Mux_DATA_SIZE32_9 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(9), B => din1(9), S => sel, Z => dout(9));
   U2 : MUX2_X1 port map( A => din0(8), B => din1(8), S => sel, Z => dout(8));
   U3 : MUX2_X1 port map( A => din0(7), B => din1(7), S => sel, Z => dout(7));
   U4 : MUX2_X1 port map( A => din0(6), B => din1(6), S => sel, Z => dout(6));
   U5 : MUX2_X1 port map( A => din0(5), B => din1(5), S => sel, Z => dout(5));
   U6 : MUX2_X1 port map( A => din0(4), B => din1(4), S => sel, Z => dout(4));
   U7 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U8 : MUX2_X1 port map( A => din0(31), B => din1(31), S => sel, Z => dout(31)
                           );
   U9 : MUX2_X1 port map( A => din0(30), B => din1(30), S => sel, Z => dout(30)
                           );
   U10 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U11 : MUX2_X1 port map( A => din0(29), B => din1(29), S => sel, Z => 
                           dout(29));
   U12 : MUX2_X1 port map( A => din0(28), B => din1(28), S => sel, Z => 
                           dout(28));
   U13 : MUX2_X1 port map( A => din0(27), B => din1(27), S => sel, Z => 
                           dout(27));
   U14 : MUX2_X1 port map( A => din0(26), B => din1(26), S => sel, Z => 
                           dout(26));
   U15 : MUX2_X1 port map( A => din0(25), B => din1(25), S => sel, Z => 
                           dout(25));
   U16 : MUX2_X1 port map( A => din0(24), B => din1(24), S => sel, Z => 
                           dout(24));
   U17 : MUX2_X1 port map( A => din0(23), B => din1(23), S => sel, Z => 
                           dout(23));
   U18 : MUX2_X1 port map( A => din0(22), B => din1(22), S => sel, Z => 
                           dout(22));
   U19 : MUX2_X1 port map( A => din0(21), B => din1(21), S => sel, Z => 
                           dout(21));
   U20 : MUX2_X1 port map( A => din0(20), B => din1(20), S => sel, Z => 
                           dout(20));
   U21 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U22 : MUX2_X1 port map( A => din0(19), B => din1(19), S => sel, Z => 
                           dout(19));
   U23 : MUX2_X1 port map( A => din0(18), B => din1(18), S => sel, Z => 
                           dout(18));
   U24 : MUX2_X1 port map( A => din0(17), B => din1(17), S => sel, Z => 
                           dout(17));
   U25 : MUX2_X1 port map( A => din0(16), B => din1(16), S => sel, Z => 
                           dout(16));
   U26 : MUX2_X1 port map( A => din0(15), B => din1(15), S => sel, Z => 
                           dout(15));
   U27 : MUX2_X1 port map( A => din0(14), B => din1(14), S => sel, Z => 
                           dout(14));
   U28 : MUX2_X1 port map( A => din0(13), B => din1(13), S => sel, Z => 
                           dout(13));
   U29 : MUX2_X1 port map( A => din0(12), B => din1(12), S => sel, Z => 
                           dout(12));
   U30 : MUX2_X1 port map( A => din0(11), B => din1(11), S => sel, Z => 
                           dout(11));
   U31 : MUX2_X1 port map( A => din0(10), B => din1(10), S => sel, Z => 
                           dout(10));
   U32 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE32_8 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0);  
         dout : out std_logic_vector (31 downto 0));

end Mux_DATA_SIZE32_8;

architecture SYN_mux_arch of Mux_DATA_SIZE32_8 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(9), B => din1(9), S => sel, Z => dout(9));
   U2 : MUX2_X1 port map( A => din0(8), B => din1(8), S => sel, Z => dout(8));
   U3 : MUX2_X1 port map( A => din0(7), B => din1(7), S => sel, Z => dout(7));
   U4 : MUX2_X1 port map( A => din0(6), B => din1(6), S => sel, Z => dout(6));
   U5 : MUX2_X1 port map( A => din0(5), B => din1(5), S => sel, Z => dout(5));
   U6 : MUX2_X1 port map( A => din0(4), B => din1(4), S => sel, Z => dout(4));
   U7 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U8 : MUX2_X1 port map( A => din0(31), B => din1(31), S => sel, Z => dout(31)
                           );
   U9 : MUX2_X1 port map( A => din0(30), B => din1(30), S => sel, Z => dout(30)
                           );
   U10 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U11 : MUX2_X1 port map( A => din0(29), B => din1(29), S => sel, Z => 
                           dout(29));
   U12 : MUX2_X1 port map( A => din0(28), B => din1(28), S => sel, Z => 
                           dout(28));
   U13 : MUX2_X1 port map( A => din0(27), B => din1(27), S => sel, Z => 
                           dout(27));
   U14 : MUX2_X1 port map( A => din0(26), B => din1(26), S => sel, Z => 
                           dout(26));
   U15 : MUX2_X1 port map( A => din0(25), B => din1(25), S => sel, Z => 
                           dout(25));
   U16 : MUX2_X1 port map( A => din0(24), B => din1(24), S => sel, Z => 
                           dout(24));
   U17 : MUX2_X1 port map( A => din0(23), B => din1(23), S => sel, Z => 
                           dout(23));
   U18 : MUX2_X1 port map( A => din0(22), B => din1(22), S => sel, Z => 
                           dout(22));
   U19 : MUX2_X1 port map( A => din0(21), B => din1(21), S => sel, Z => 
                           dout(21));
   U20 : MUX2_X1 port map( A => din0(20), B => din1(20), S => sel, Z => 
                           dout(20));
   U21 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U22 : MUX2_X1 port map( A => din0(19), B => din1(19), S => sel, Z => 
                           dout(19));
   U23 : MUX2_X1 port map( A => din0(18), B => din1(18), S => sel, Z => 
                           dout(18));
   U24 : MUX2_X1 port map( A => din0(17), B => din1(17), S => sel, Z => 
                           dout(17));
   U25 : MUX2_X1 port map( A => din0(16), B => din1(16), S => sel, Z => 
                           dout(16));
   U26 : MUX2_X1 port map( A => din0(15), B => din1(15), S => sel, Z => 
                           dout(15));
   U27 : MUX2_X1 port map( A => din0(14), B => din1(14), S => sel, Z => 
                           dout(14));
   U28 : MUX2_X1 port map( A => din0(13), B => din1(13), S => sel, Z => 
                           dout(13));
   U29 : MUX2_X1 port map( A => din0(12), B => din1(12), S => sel, Z => 
                           dout(12));
   U30 : MUX2_X1 port map( A => din0(11), B => din1(11), S => sel, Z => 
                           dout(11));
   U31 : MUX2_X1 port map( A => din0(10), B => din1(10), S => sel, Z => 
                           dout(10));
   U32 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE32_7 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0);  
         dout : out std_logic_vector (31 downto 0));

end Mux_DATA_SIZE32_7;

architecture SYN_mux_arch of Mux_DATA_SIZE32_7 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(9), B => din1(9), S => sel, Z => dout(9));
   U2 : MUX2_X1 port map( A => din0(8), B => din1(8), S => sel, Z => dout(8));
   U3 : MUX2_X1 port map( A => din0(7), B => din1(7), S => sel, Z => dout(7));
   U4 : MUX2_X1 port map( A => din0(6), B => din1(6), S => sel, Z => dout(6));
   U5 : MUX2_X1 port map( A => din0(5), B => din1(5), S => sel, Z => dout(5));
   U6 : MUX2_X1 port map( A => din0(4), B => din1(4), S => sel, Z => dout(4));
   U7 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U8 : MUX2_X1 port map( A => din0(31), B => din1(31), S => sel, Z => dout(31)
                           );
   U9 : MUX2_X1 port map( A => din0(30), B => din1(30), S => sel, Z => dout(30)
                           );
   U10 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U11 : MUX2_X1 port map( A => din0(29), B => din1(29), S => sel, Z => 
                           dout(29));
   U12 : MUX2_X1 port map( A => din0(28), B => din1(28), S => sel, Z => 
                           dout(28));
   U13 : MUX2_X1 port map( A => din0(27), B => din1(27), S => sel, Z => 
                           dout(27));
   U14 : MUX2_X1 port map( A => din0(26), B => din1(26), S => sel, Z => 
                           dout(26));
   U15 : MUX2_X1 port map( A => din0(25), B => din1(25), S => sel, Z => 
                           dout(25));
   U16 : MUX2_X1 port map( A => din0(24), B => din1(24), S => sel, Z => 
                           dout(24));
   U17 : MUX2_X1 port map( A => din0(23), B => din1(23), S => sel, Z => 
                           dout(23));
   U18 : MUX2_X1 port map( A => din0(22), B => din1(22), S => sel, Z => 
                           dout(22));
   U19 : MUX2_X1 port map( A => din0(21), B => din1(21), S => sel, Z => 
                           dout(21));
   U20 : MUX2_X1 port map( A => din0(20), B => din1(20), S => sel, Z => 
                           dout(20));
   U21 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U22 : MUX2_X1 port map( A => din0(19), B => din1(19), S => sel, Z => 
                           dout(19));
   U23 : MUX2_X1 port map( A => din0(18), B => din1(18), S => sel, Z => 
                           dout(18));
   U24 : MUX2_X1 port map( A => din0(17), B => din1(17), S => sel, Z => 
                           dout(17));
   U25 : MUX2_X1 port map( A => din0(16), B => din1(16), S => sel, Z => 
                           dout(16));
   U26 : MUX2_X1 port map( A => din0(15), B => din1(15), S => sel, Z => 
                           dout(15));
   U27 : MUX2_X1 port map( A => din0(14), B => din1(14), S => sel, Z => 
                           dout(14));
   U28 : MUX2_X1 port map( A => din0(13), B => din1(13), S => sel, Z => 
                           dout(13));
   U29 : MUX2_X1 port map( A => din0(12), B => din1(12), S => sel, Z => 
                           dout(12));
   U30 : MUX2_X1 port map( A => din0(11), B => din1(11), S => sel, Z => 
                           dout(11));
   U31 : MUX2_X1 port map( A => din0(10), B => din1(10), S => sel, Z => 
                           dout(10));
   U32 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE32_6 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0);  
         dout : out std_logic_vector (31 downto 0));

end Mux_DATA_SIZE32_6;

architecture SYN_mux_arch of Mux_DATA_SIZE32_6 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(9), B => din1(9), S => sel, Z => dout(9));
   U2 : MUX2_X1 port map( A => din0(8), B => din1(8), S => sel, Z => dout(8));
   U3 : MUX2_X1 port map( A => din0(7), B => din1(7), S => sel, Z => dout(7));
   U4 : MUX2_X1 port map( A => din0(6), B => din1(6), S => sel, Z => dout(6));
   U5 : MUX2_X1 port map( A => din0(5), B => din1(5), S => sel, Z => dout(5));
   U6 : MUX2_X1 port map( A => din0(4), B => din1(4), S => sel, Z => dout(4));
   U7 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U8 : MUX2_X1 port map( A => din0(31), B => din1(31), S => sel, Z => dout(31)
                           );
   U9 : MUX2_X1 port map( A => din0(30), B => din1(30), S => sel, Z => dout(30)
                           );
   U10 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U11 : MUX2_X1 port map( A => din0(29), B => din1(29), S => sel, Z => 
                           dout(29));
   U12 : MUX2_X1 port map( A => din0(28), B => din1(28), S => sel, Z => 
                           dout(28));
   U13 : MUX2_X1 port map( A => din0(27), B => din1(27), S => sel, Z => 
                           dout(27));
   U14 : MUX2_X1 port map( A => din0(26), B => din1(26), S => sel, Z => 
                           dout(26));
   U15 : MUX2_X1 port map( A => din0(25), B => din1(25), S => sel, Z => 
                           dout(25));
   U16 : MUX2_X1 port map( A => din0(24), B => din1(24), S => sel, Z => 
                           dout(24));
   U17 : MUX2_X1 port map( A => din0(23), B => din1(23), S => sel, Z => 
                           dout(23));
   U18 : MUX2_X1 port map( A => din0(22), B => din1(22), S => sel, Z => 
                           dout(22));
   U19 : MUX2_X1 port map( A => din0(21), B => din1(21), S => sel, Z => 
                           dout(21));
   U20 : MUX2_X1 port map( A => din0(20), B => din1(20), S => sel, Z => 
                           dout(20));
   U21 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U22 : MUX2_X1 port map( A => din0(19), B => din1(19), S => sel, Z => 
                           dout(19));
   U23 : MUX2_X1 port map( A => din0(18), B => din1(18), S => sel, Z => 
                           dout(18));
   U24 : MUX2_X1 port map( A => din0(17), B => din1(17), S => sel, Z => 
                           dout(17));
   U25 : MUX2_X1 port map( A => din0(16), B => din1(16), S => sel, Z => 
                           dout(16));
   U26 : MUX2_X1 port map( A => din0(15), B => din1(15), S => sel, Z => 
                           dout(15));
   U27 : MUX2_X1 port map( A => din0(14), B => din1(14), S => sel, Z => 
                           dout(14));
   U28 : MUX2_X1 port map( A => din0(13), B => din1(13), S => sel, Z => 
                           dout(13));
   U29 : MUX2_X1 port map( A => din0(12), B => din1(12), S => sel, Z => 
                           dout(12));
   U30 : MUX2_X1 port map( A => din0(11), B => din1(11), S => sel, Z => 
                           dout(11));
   U31 : MUX2_X1 port map( A => din0(10), B => din1(10), S => sel, Z => 
                           dout(10));
   U32 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE32_5 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0);  
         dout : out std_logic_vector (31 downto 0));

end Mux_DATA_SIZE32_5;

architecture SYN_mux_arch of Mux_DATA_SIZE32_5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(9), B => din1(9), S => sel, Z => dout(9));
   U2 : MUX2_X1 port map( A => din0(8), B => din1(8), S => sel, Z => dout(8));
   U3 : MUX2_X1 port map( A => din0(7), B => din1(7), S => sel, Z => dout(7));
   U4 : MUX2_X1 port map( A => din0(6), B => din1(6), S => sel, Z => dout(6));
   U5 : MUX2_X1 port map( A => din0(5), B => din1(5), S => sel, Z => dout(5));
   U6 : MUX2_X1 port map( A => din0(4), B => din1(4), S => sel, Z => dout(4));
   U7 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U8 : MUX2_X1 port map( A => din0(31), B => din1(31), S => sel, Z => dout(31)
                           );
   U9 : MUX2_X1 port map( A => din0(30), B => din1(30), S => sel, Z => dout(30)
                           );
   U10 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U11 : MUX2_X1 port map( A => din0(29), B => din1(29), S => sel, Z => 
                           dout(29));
   U12 : MUX2_X1 port map( A => din0(28), B => din1(28), S => sel, Z => 
                           dout(28));
   U13 : MUX2_X1 port map( A => din0(27), B => din1(27), S => sel, Z => 
                           dout(27));
   U14 : MUX2_X1 port map( A => din0(26), B => din1(26), S => sel, Z => 
                           dout(26));
   U15 : MUX2_X1 port map( A => din0(25), B => din1(25), S => sel, Z => 
                           dout(25));
   U16 : MUX2_X1 port map( A => din0(24), B => din1(24), S => sel, Z => 
                           dout(24));
   U17 : MUX2_X1 port map( A => din0(23), B => din1(23), S => sel, Z => 
                           dout(23));
   U18 : MUX2_X1 port map( A => din0(22), B => din1(22), S => sel, Z => 
                           dout(22));
   U19 : MUX2_X1 port map( A => din0(21), B => din1(21), S => sel, Z => 
                           dout(21));
   U20 : MUX2_X1 port map( A => din0(20), B => din1(20), S => sel, Z => 
                           dout(20));
   U21 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U22 : MUX2_X1 port map( A => din0(19), B => din1(19), S => sel, Z => 
                           dout(19));
   U23 : MUX2_X1 port map( A => din0(18), B => din1(18), S => sel, Z => 
                           dout(18));
   U24 : MUX2_X1 port map( A => din0(17), B => din1(17), S => sel, Z => 
                           dout(17));
   U25 : MUX2_X1 port map( A => din0(16), B => din1(16), S => sel, Z => 
                           dout(16));
   U26 : MUX2_X1 port map( A => din0(15), B => din1(15), S => sel, Z => 
                           dout(15));
   U27 : MUX2_X1 port map( A => din0(14), B => din1(14), S => sel, Z => 
                           dout(14));
   U28 : MUX2_X1 port map( A => din0(13), B => din1(13), S => sel, Z => 
                           dout(13));
   U29 : MUX2_X1 port map( A => din0(12), B => din1(12), S => sel, Z => 
                           dout(12));
   U30 : MUX2_X1 port map( A => din0(11), B => din1(11), S => sel, Z => 
                           dout(11));
   U31 : MUX2_X1 port map( A => din0(10), B => din1(10), S => sel, Z => 
                           dout(10));
   U32 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE32_4 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0);  
         dout : out std_logic_vector (31 downto 0));

end Mux_DATA_SIZE32_4;

architecture SYN_mux_arch of Mux_DATA_SIZE32_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(9), B => din1(9), S => sel, Z => dout(9));
   U2 : MUX2_X1 port map( A => din0(8), B => din1(8), S => sel, Z => dout(8));
   U3 : MUX2_X1 port map( A => din0(7), B => din1(7), S => sel, Z => dout(7));
   U4 : MUX2_X1 port map( A => din0(6), B => din1(6), S => sel, Z => dout(6));
   U5 : MUX2_X1 port map( A => din0(5), B => din1(5), S => sel, Z => dout(5));
   U6 : MUX2_X1 port map( A => din0(4), B => din1(4), S => sel, Z => dout(4));
   U7 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U8 : MUX2_X1 port map( A => din0(31), B => din1(31), S => sel, Z => dout(31)
                           );
   U9 : MUX2_X1 port map( A => din0(30), B => din1(30), S => sel, Z => dout(30)
                           );
   U10 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U11 : MUX2_X1 port map( A => din0(29), B => din1(29), S => sel, Z => 
                           dout(29));
   U12 : MUX2_X1 port map( A => din0(28), B => din1(28), S => sel, Z => 
                           dout(28));
   U13 : MUX2_X1 port map( A => din0(27), B => din1(27), S => sel, Z => 
                           dout(27));
   U14 : MUX2_X1 port map( A => din0(26), B => din1(26), S => sel, Z => 
                           dout(26));
   U15 : MUX2_X1 port map( A => din0(25), B => din1(25), S => sel, Z => 
                           dout(25));
   U16 : MUX2_X1 port map( A => din0(24), B => din1(24), S => sel, Z => 
                           dout(24));
   U17 : MUX2_X1 port map( A => din0(23), B => din1(23), S => sel, Z => 
                           dout(23));
   U18 : MUX2_X1 port map( A => din0(22), B => din1(22), S => sel, Z => 
                           dout(22));
   U19 : MUX2_X1 port map( A => din0(21), B => din1(21), S => sel, Z => 
                           dout(21));
   U20 : MUX2_X1 port map( A => din0(20), B => din1(20), S => sel, Z => 
                           dout(20));
   U21 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U22 : MUX2_X1 port map( A => din0(19), B => din1(19), S => sel, Z => 
                           dout(19));
   U23 : MUX2_X1 port map( A => din0(18), B => din1(18), S => sel, Z => 
                           dout(18));
   U24 : MUX2_X1 port map( A => din0(17), B => din1(17), S => sel, Z => 
                           dout(17));
   U25 : MUX2_X1 port map( A => din0(16), B => din1(16), S => sel, Z => 
                           dout(16));
   U26 : MUX2_X1 port map( A => din0(15), B => din1(15), S => sel, Z => 
                           dout(15));
   U27 : MUX2_X1 port map( A => din0(14), B => din1(14), S => sel, Z => 
                           dout(14));
   U28 : MUX2_X1 port map( A => din0(13), B => din1(13), S => sel, Z => 
                           dout(13));
   U29 : MUX2_X1 port map( A => din0(12), B => din1(12), S => sel, Z => 
                           dout(12));
   U30 : MUX2_X1 port map( A => din0(11), B => din1(11), S => sel, Z => 
                           dout(11));
   U31 : MUX2_X1 port map( A => din0(10), B => din1(10), S => sel, Z => 
                           dout(10));
   U32 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE32_3 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0);  
         dout : out std_logic_vector (31 downto 0));

end Mux_DATA_SIZE32_3;

architecture SYN_mux_arch of Mux_DATA_SIZE32_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X8
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11, n12, n1, n3, n5, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n10, ZN => n1);
   U2 : INV_X8 port map( A => n1, ZN => dout(2));
   U3 : INV_X1 port map( A => n9, ZN => n3);
   U4 : INV_X8 port map( A => n3, ZN => dout(3));
   U5 : INV_X1 port map( A => n12, ZN => n5);
   U6 : INV_X8 port map( A => n5, ZN => dout(0));
   U7 : INV_X1 port map( A => n11, ZN => n7);
   U8 : INV_X8 port map( A => n7, ZN => dout(1));
   U9 : MUX2_X1 port map( A => din0(9), B => din1(9), S => sel, Z => dout(9));
   U10 : MUX2_X1 port map( A => din0(8), B => din1(8), S => sel, Z => dout(8));
   U11 : MUX2_X1 port map( A => din0(7), B => din1(7), S => sel, Z => dout(7));
   U12 : MUX2_X1 port map( A => din0(6), B => din1(6), S => sel, Z => dout(6));
   U13 : MUX2_X1 port map( A => din0(5), B => din1(5), S => sel, Z => dout(5));
   U14 : MUX2_X1 port map( A => din0(4), B => din1(4), S => sel, Z => dout(4));
   U15 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => n9);
   U16 : MUX2_X1 port map( A => din0(31), B => din1(31), S => sel, Z => 
                           dout(31));
   U17 : MUX2_X1 port map( A => din0(30), B => din1(30), S => sel, Z => 
                           dout(30));
   U18 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => n10);
   U19 : MUX2_X1 port map( A => din0(29), B => din1(29), S => sel, Z => 
                           dout(29));
   U20 : MUX2_X1 port map( A => din0(28), B => din1(28), S => sel, Z => 
                           dout(28));
   U21 : MUX2_X1 port map( A => din0(27), B => din1(27), S => sel, Z => 
                           dout(27));
   U22 : MUX2_X1 port map( A => din0(26), B => din1(26), S => sel, Z => 
                           dout(26));
   U23 : MUX2_X1 port map( A => din0(25), B => din1(25), S => sel, Z => 
                           dout(25));
   U24 : MUX2_X1 port map( A => din0(24), B => din1(24), S => sel, Z => 
                           dout(24));
   U25 : MUX2_X1 port map( A => din0(23), B => din1(23), S => sel, Z => 
                           dout(23));
   U26 : MUX2_X1 port map( A => din0(22), B => din1(22), S => sel, Z => 
                           dout(22));
   U27 : MUX2_X1 port map( A => din0(21), B => din1(21), S => sel, Z => 
                           dout(21));
   U28 : MUX2_X1 port map( A => din0(20), B => din1(20), S => sel, Z => 
                           dout(20));
   U29 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => n11);
   U30 : MUX2_X1 port map( A => din0(19), B => din1(19), S => sel, Z => 
                           dout(19));
   U31 : MUX2_X1 port map( A => din0(18), B => din1(18), S => sel, Z => 
                           dout(18));
   U32 : MUX2_X1 port map( A => din0(17), B => din1(17), S => sel, Z => 
                           dout(17));
   U33 : MUX2_X1 port map( A => din0(16), B => din1(16), S => sel, Z => 
                           dout(16));
   U34 : MUX2_X1 port map( A => din0(15), B => din1(15), S => sel, Z => 
                           dout(15));
   U35 : MUX2_X1 port map( A => din0(14), B => din1(14), S => sel, Z => 
                           dout(14));
   U36 : MUX2_X1 port map( A => din0(13), B => din1(13), S => sel, Z => 
                           dout(13));
   U37 : MUX2_X1 port map( A => din0(12), B => din1(12), S => sel, Z => 
                           dout(12));
   U38 : MUX2_X1 port map( A => din0(11), B => din1(11), S => sel, Z => 
                           dout(11));
   U39 : MUX2_X1 port map( A => din0(10), B => din1(10), S => sel, Z => 
                           dout(10));
   U40 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => n12);

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE32_2 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0);  
         dout : out std_logic_vector (31 downto 0));

end Mux_DATA_SIZE32_2;

architecture SYN_mux_arch of Mux_DATA_SIZE32_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(9), B => din1(9), S => sel, Z => dout(9));
   U2 : MUX2_X1 port map( A => din0(8), B => din1(8), S => sel, Z => dout(8));
   U3 : MUX2_X1 port map( A => din0(7), B => din1(7), S => sel, Z => dout(7));
   U4 : MUX2_X1 port map( A => din0(6), B => din1(6), S => sel, Z => dout(6));
   U5 : MUX2_X1 port map( A => din0(5), B => din1(5), S => sel, Z => dout(5));
   U6 : MUX2_X1 port map( A => din0(4), B => din1(4), S => sel, Z => dout(4));
   U7 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U8 : MUX2_X1 port map( A => din0(31), B => din1(31), S => sel, Z => dout(31)
                           );
   U9 : MUX2_X1 port map( A => din0(30), B => din1(30), S => sel, Z => dout(30)
                           );
   U10 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U11 : MUX2_X1 port map( A => din0(29), B => din1(29), S => sel, Z => 
                           dout(29));
   U12 : MUX2_X1 port map( A => din0(28), B => din1(28), S => sel, Z => 
                           dout(28));
   U13 : MUX2_X1 port map( A => din0(27), B => din1(27), S => sel, Z => 
                           dout(27));
   U14 : MUX2_X1 port map( A => din0(26), B => din1(26), S => sel, Z => 
                           dout(26));
   U15 : MUX2_X1 port map( A => din0(25), B => din1(25), S => sel, Z => 
                           dout(25));
   U16 : MUX2_X1 port map( A => din0(24), B => din1(24), S => sel, Z => 
                           dout(24));
   U17 : MUX2_X1 port map( A => din0(23), B => din1(23), S => sel, Z => 
                           dout(23));
   U18 : MUX2_X1 port map( A => din0(22), B => din1(22), S => sel, Z => 
                           dout(22));
   U19 : MUX2_X1 port map( A => din0(21), B => din1(21), S => sel, Z => 
                           dout(21));
   U20 : MUX2_X1 port map( A => din0(20), B => din1(20), S => sel, Z => 
                           dout(20));
   U21 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U22 : MUX2_X1 port map( A => din0(19), B => din1(19), S => sel, Z => 
                           dout(19));
   U23 : MUX2_X1 port map( A => din0(18), B => din1(18), S => sel, Z => 
                           dout(18));
   U24 : MUX2_X1 port map( A => din0(17), B => din1(17), S => sel, Z => 
                           dout(17));
   U25 : MUX2_X1 port map( A => din0(16), B => din1(16), S => sel, Z => 
                           dout(16));
   U26 : MUX2_X1 port map( A => din0(15), B => din1(15), S => sel, Z => 
                           dout(15));
   U27 : MUX2_X1 port map( A => din0(14), B => din1(14), S => sel, Z => 
                           dout(14));
   U28 : MUX2_X1 port map( A => din0(13), B => din1(13), S => sel, Z => 
                           dout(13));
   U29 : MUX2_X1 port map( A => din0(12), B => din1(12), S => sel, Z => 
                           dout(12));
   U30 : MUX2_X1 port map( A => din0(11), B => din1(11), S => sel, Z => 
                           dout(11));
   U31 : MUX2_X1 port map( A => din0(10), B => din1(10), S => sel, Z => 
                           dout(10));
   U32 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE32_1 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0);  
         dout : out std_logic_vector (31 downto 0));

end Mux_DATA_SIZE32_1;

architecture SYN_mux_arch of Mux_DATA_SIZE32_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(9), B => din1(9), S => sel, Z => dout(9));
   U2 : MUX2_X1 port map( A => din0(8), B => din1(8), S => sel, Z => dout(8));
   U3 : MUX2_X1 port map( A => din0(7), B => din1(7), S => sel, Z => dout(7));
   U4 : MUX2_X1 port map( A => din0(6), B => din1(6), S => sel, Z => dout(6));
   U5 : MUX2_X1 port map( A => din0(5), B => din1(5), S => sel, Z => dout(5));
   U6 : MUX2_X1 port map( A => din0(4), B => din1(4), S => sel, Z => dout(4));
   U7 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U8 : MUX2_X1 port map( A => din0(31), B => din1(31), S => sel, Z => dout(31)
                           );
   U9 : MUX2_X1 port map( A => din0(30), B => din1(30), S => sel, Z => dout(30)
                           );
   U10 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U11 : MUX2_X1 port map( A => din0(29), B => din1(29), S => sel, Z => 
                           dout(29));
   U12 : MUX2_X1 port map( A => din0(28), B => din1(28), S => sel, Z => 
                           dout(28));
   U13 : MUX2_X1 port map( A => din0(27), B => din1(27), S => sel, Z => 
                           dout(27));
   U14 : MUX2_X1 port map( A => din0(26), B => din1(26), S => sel, Z => 
                           dout(26));
   U15 : MUX2_X1 port map( A => din0(25), B => din1(25), S => sel, Z => 
                           dout(25));
   U16 : MUX2_X1 port map( A => din0(24), B => din1(24), S => sel, Z => 
                           dout(24));
   U17 : MUX2_X1 port map( A => din0(23), B => din1(23), S => sel, Z => 
                           dout(23));
   U18 : MUX2_X1 port map( A => din0(22), B => din1(22), S => sel, Z => 
                           dout(22));
   U19 : MUX2_X1 port map( A => din0(21), B => din1(21), S => sel, Z => 
                           dout(21));
   U20 : MUX2_X1 port map( A => din0(20), B => din1(20), S => sel, Z => 
                           dout(20));
   U21 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U22 : MUX2_X1 port map( A => din0(19), B => din1(19), S => sel, Z => 
                           dout(19));
   U23 : MUX2_X1 port map( A => din0(18), B => din1(18), S => sel, Z => 
                           dout(18));
   U24 : MUX2_X1 port map( A => din0(17), B => din1(17), S => sel, Z => 
                           dout(17));
   U25 : MUX2_X1 port map( A => din0(16), B => din1(16), S => sel, Z => 
                           dout(16));
   U26 : MUX2_X1 port map( A => din0(15), B => din1(15), S => sel, Z => 
                           dout(15));
   U27 : MUX2_X1 port map( A => din0(14), B => din1(14), S => sel, Z => 
                           dout(14));
   U28 : MUX2_X1 port map( A => din0(13), B => din1(13), S => sel, Z => 
                           dout(13));
   U29 : MUX2_X1 port map( A => din0(12), B => din1(12), S => sel, Z => 
                           dout(12));
   U30 : MUX2_X1 port map( A => din0(11), B => din1(11), S => sel, Z => 
                           dout(11));
   U31 : MUX2_X1 port map( A => din0(10), B => din1(10), S => sel, Z => 
                           dout(10));
   U32 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Adder_DATA_SIZE32_7 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end Adder_DATA_SIZE32_7;

architecture SYN_adder_arch of Adder_DATA_SIZE32_7 is

   component P4Adder_DATA_SIZE32_SPARSITY4_7
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;

begin
   
   ADDER0 : P4Adder_DATA_SIZE32_SPARSITY4_7 port map( cin => cin, a(31) => 
                           a(31), a(30) => a(30), a(29) => a(29), a(28) => 
                           a(28), a(27) => a(27), a(26) => a(26), a(25) => 
                           a(25), a(24) => a(24), a(23) => a(23), a(22) => 
                           a(22), a(21) => a(21), a(20) => a(20), a(19) => 
                           a(19), a(18) => a(18), a(17) => a(17), a(16) => 
                           a(16), a(15) => a(15), a(14) => a(14), a(13) => 
                           a(13), a(12) => a(12), a(11) => a(11), a(10) => 
                           a(10), a(9) => a(9), a(8) => a(8), a(7) => a(7), 
                           a(6) => a(6), a(5) => a(5), a(4) => a(4), a(3) => 
                           a(3), a(2) => a(2), a(1) => a(1), a(0) => a(0), 
                           b(31) => b(31), b(30) => b(30), b(29) => b(29), 
                           b(28) => b(28), b(27) => b(27), b(26) => b(26), 
                           b(25) => b(25), b(24) => b(24), b(23) => b(23), 
                           b(22) => b(22), b(21) => b(21), b(20) => b(20), 
                           b(19) => b(19), b(18) => b(18), b(17) => b(17), 
                           b(16) => b(16), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           s(31) => s(31), s(30) => s(30), s(29) => s(29), 
                           s(28) => s(28), s(27) => s(27), s(26) => s(26), 
                           s(25) => s(25), s(24) => s(24), s(23) => s(23), 
                           s(22) => s(22), s(21) => s(21), s(20) => s(20), 
                           s(19) => s(19), s(18) => s(18), s(17) => s(17), 
                           s(16) => s(16), s(15) => s(15), s(14) => s(14), 
                           s(13) => s(13), s(12) => s(12), s(11) => s(11), 
                           s(10) => s(10), s(9) => s(9), s(8) => s(8), s(7) => 
                           s(7), s(6) => s(6), s(5) => s(5), s(4) => s(4), s(3)
                           => s(3), s(2) => s(2), s(1) => s(1), s(0) => s(0), 
                           cout => cout);

end SYN_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Adder_DATA_SIZE32_6 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end Adder_DATA_SIZE32_6;

architecture SYN_adder_arch of Adder_DATA_SIZE32_6 is

   component P4Adder_DATA_SIZE32_SPARSITY4_6
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;

begin
   
   ADDER0 : P4Adder_DATA_SIZE32_SPARSITY4_6 port map( cin => cin, a(31) => 
                           a(31), a(30) => a(30), a(29) => a(29), a(28) => 
                           a(28), a(27) => a(27), a(26) => a(26), a(25) => 
                           a(25), a(24) => a(24), a(23) => a(23), a(22) => 
                           a(22), a(21) => a(21), a(20) => a(20), a(19) => 
                           a(19), a(18) => a(18), a(17) => a(17), a(16) => 
                           a(16), a(15) => a(15), a(14) => a(14), a(13) => 
                           a(13), a(12) => a(12), a(11) => a(11), a(10) => 
                           a(10), a(9) => a(9), a(8) => a(8), a(7) => a(7), 
                           a(6) => a(6), a(5) => a(5), a(4) => a(4), a(3) => 
                           a(3), a(2) => a(2), a(1) => a(1), a(0) => a(0), 
                           b(31) => b(31), b(30) => b(30), b(29) => b(29), 
                           b(28) => b(28), b(27) => b(27), b(26) => b(26), 
                           b(25) => b(25), b(24) => b(24), b(23) => b(23), 
                           b(22) => b(22), b(21) => b(21), b(20) => b(20), 
                           b(19) => b(19), b(18) => b(18), b(17) => b(17), 
                           b(16) => b(16), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           s(31) => s(31), s(30) => s(30), s(29) => s(29), 
                           s(28) => s(28), s(27) => s(27), s(26) => s(26), 
                           s(25) => s(25), s(24) => s(24), s(23) => s(23), 
                           s(22) => s(22), s(21) => s(21), s(20) => s(20), 
                           s(19) => s(19), s(18) => s(18), s(17) => s(17), 
                           s(16) => s(16), s(15) => s(15), s(14) => s(14), 
                           s(13) => s(13), s(12) => s(12), s(11) => s(11), 
                           s(10) => s(10), s(9) => s(9), s(8) => s(8), s(7) => 
                           s(7), s(6) => s(6), s(5) => s(5), s(4) => s(4), s(3)
                           => s(3), s(2) => s(2), s(1) => s(1), s(0) => s(0), 
                           cout => cout);

end SYN_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Adder_DATA_SIZE32_5 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end Adder_DATA_SIZE32_5;

architecture SYN_adder_arch of Adder_DATA_SIZE32_5 is

   component P4Adder_DATA_SIZE32_SPARSITY4_5
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;

begin
   
   ADDER0 : P4Adder_DATA_SIZE32_SPARSITY4_5 port map( cin => cin, a(31) => 
                           a(31), a(30) => a(30), a(29) => a(29), a(28) => 
                           a(28), a(27) => a(27), a(26) => a(26), a(25) => 
                           a(25), a(24) => a(24), a(23) => a(23), a(22) => 
                           a(22), a(21) => a(21), a(20) => a(20), a(19) => 
                           a(19), a(18) => a(18), a(17) => a(17), a(16) => 
                           a(16), a(15) => a(15), a(14) => a(14), a(13) => 
                           a(13), a(12) => a(12), a(11) => a(11), a(10) => 
                           a(10), a(9) => a(9), a(8) => a(8), a(7) => a(7), 
                           a(6) => a(6), a(5) => a(5), a(4) => a(4), a(3) => 
                           a(3), a(2) => a(2), a(1) => a(1), a(0) => a(0), 
                           b(31) => b(31), b(30) => b(30), b(29) => b(29), 
                           b(28) => b(28), b(27) => b(27), b(26) => b(26), 
                           b(25) => b(25), b(24) => b(24), b(23) => b(23), 
                           b(22) => b(22), b(21) => b(21), b(20) => b(20), 
                           b(19) => b(19), b(18) => b(18), b(17) => b(17), 
                           b(16) => b(16), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           s(31) => s(31), s(30) => s(30), s(29) => s(29), 
                           s(28) => s(28), s(27) => s(27), s(26) => s(26), 
                           s(25) => s(25), s(24) => s(24), s(23) => s(23), 
                           s(22) => s(22), s(21) => s(21), s(20) => s(20), 
                           s(19) => s(19), s(18) => s(18), s(17) => s(17), 
                           s(16) => s(16), s(15) => s(15), s(14) => s(14), 
                           s(13) => s(13), s(12) => s(12), s(11) => s(11), 
                           s(10) => s(10), s(9) => s(9), s(8) => s(8), s(7) => 
                           s(7), s(6) => s(6), s(5) => s(5), s(4) => s(4), s(3)
                           => s(3), s(2) => s(2), s(1) => s(1), s(0) => s(0), 
                           cout => cout);

end SYN_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Adder_DATA_SIZE32_4 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end Adder_DATA_SIZE32_4;

architecture SYN_adder_arch of Adder_DATA_SIZE32_4 is

   component P4Adder_DATA_SIZE32_SPARSITY4_4
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;

begin
   
   ADDER0 : P4Adder_DATA_SIZE32_SPARSITY4_4 port map( cin => cin, a(31) => 
                           a(31), a(30) => a(30), a(29) => a(29), a(28) => 
                           a(28), a(27) => a(27), a(26) => a(26), a(25) => 
                           a(25), a(24) => a(24), a(23) => a(23), a(22) => 
                           a(22), a(21) => a(21), a(20) => a(20), a(19) => 
                           a(19), a(18) => a(18), a(17) => a(17), a(16) => 
                           a(16), a(15) => a(15), a(14) => a(14), a(13) => 
                           a(13), a(12) => a(12), a(11) => a(11), a(10) => 
                           a(10), a(9) => a(9), a(8) => a(8), a(7) => a(7), 
                           a(6) => a(6), a(5) => a(5), a(4) => a(4), a(3) => 
                           a(3), a(2) => a(2), a(1) => a(1), a(0) => a(0), 
                           b(31) => b(31), b(30) => b(30), b(29) => b(29), 
                           b(28) => b(28), b(27) => b(27), b(26) => b(26), 
                           b(25) => b(25), b(24) => b(24), b(23) => b(23), 
                           b(22) => b(22), b(21) => b(21), b(20) => b(20), 
                           b(19) => b(19), b(18) => b(18), b(17) => b(17), 
                           b(16) => b(16), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           s(31) => s(31), s(30) => s(30), s(29) => s(29), 
                           s(28) => s(28), s(27) => s(27), s(26) => s(26), 
                           s(25) => s(25), s(24) => s(24), s(23) => s(23), 
                           s(22) => s(22), s(21) => s(21), s(20) => s(20), 
                           s(19) => s(19), s(18) => s(18), s(17) => s(17), 
                           s(16) => s(16), s(15) => s(15), s(14) => s(14), 
                           s(13) => s(13), s(12) => s(12), s(11) => s(11), 
                           s(10) => s(10), s(9) => s(9), s(8) => s(8), s(7) => 
                           s(7), s(6) => s(6), s(5) => s(5), s(4) => s(4), s(3)
                           => s(3), s(2) => s(2), s(1) => s(1), s(0) => s(0), 
                           cout => cout);

end SYN_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Adder_DATA_SIZE32_3 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end Adder_DATA_SIZE32_3;

architecture SYN_adder_arch of Adder_DATA_SIZE32_3 is

   component P4Adder_DATA_SIZE32_SPARSITY4_3
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;

begin
   
   ADDER0 : P4Adder_DATA_SIZE32_SPARSITY4_3 port map( cin => cin, a(31) => 
                           a(31), a(30) => a(30), a(29) => a(29), a(28) => 
                           a(28), a(27) => a(27), a(26) => a(26), a(25) => 
                           a(25), a(24) => a(24), a(23) => a(23), a(22) => 
                           a(22), a(21) => a(21), a(20) => a(20), a(19) => 
                           a(19), a(18) => a(18), a(17) => a(17), a(16) => 
                           a(16), a(15) => a(15), a(14) => a(14), a(13) => 
                           a(13), a(12) => a(12), a(11) => a(11), a(10) => 
                           a(10), a(9) => a(9), a(8) => a(8), a(7) => a(7), 
                           a(6) => a(6), a(5) => a(5), a(4) => a(4), a(3) => 
                           a(3), a(2) => a(2), a(1) => a(1), a(0) => a(0), 
                           b(31) => b(31), b(30) => b(30), b(29) => b(29), 
                           b(28) => b(28), b(27) => b(27), b(26) => b(26), 
                           b(25) => b(25), b(24) => b(24), b(23) => b(23), 
                           b(22) => b(22), b(21) => b(21), b(20) => b(20), 
                           b(19) => b(19), b(18) => b(18), b(17) => b(17), 
                           b(16) => b(16), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           s(31) => s(31), s(30) => s(30), s(29) => s(29), 
                           s(28) => s(28), s(27) => s(27), s(26) => s(26), 
                           s(25) => s(25), s(24) => s(24), s(23) => s(23), 
                           s(22) => s(22), s(21) => s(21), s(20) => s(20), 
                           s(19) => s(19), s(18) => s(18), s(17) => s(17), 
                           s(16) => s(16), s(15) => s(15), s(14) => s(14), 
                           s(13) => s(13), s(12) => s(12), s(11) => s(11), 
                           s(10) => s(10), s(9) => s(9), s(8) => s(8), s(7) => 
                           s(7), s(6) => s(6), s(5) => s(5), s(4) => s(4), s(3)
                           => s(3), s(2) => s(2), s(1) => s(1), s(0) => s(0), 
                           cout => cout);

end SYN_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Adder_DATA_SIZE32_2 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end Adder_DATA_SIZE32_2;

architecture SYN_adder_arch of Adder_DATA_SIZE32_2 is

   component P4Adder_DATA_SIZE32_SPARSITY4_2
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;

begin
   
   ADDER0 : P4Adder_DATA_SIZE32_SPARSITY4_2 port map( cin => cin, a(31) => 
                           a(31), a(30) => a(30), a(29) => a(29), a(28) => 
                           a(28), a(27) => a(27), a(26) => a(26), a(25) => 
                           a(25), a(24) => a(24), a(23) => a(23), a(22) => 
                           a(22), a(21) => a(21), a(20) => a(20), a(19) => 
                           a(19), a(18) => a(18), a(17) => a(17), a(16) => 
                           a(16), a(15) => a(15), a(14) => a(14), a(13) => 
                           a(13), a(12) => a(12), a(11) => a(11), a(10) => 
                           a(10), a(9) => a(9), a(8) => a(8), a(7) => a(7), 
                           a(6) => a(6), a(5) => a(5), a(4) => a(4), a(3) => 
                           a(3), a(2) => a(2), a(1) => a(1), a(0) => a(0), 
                           b(31) => b(31), b(30) => b(30), b(29) => b(29), 
                           b(28) => b(28), b(27) => b(27), b(26) => b(26), 
                           b(25) => b(25), b(24) => b(24), b(23) => b(23), 
                           b(22) => b(22), b(21) => b(21), b(20) => b(20), 
                           b(19) => b(19), b(18) => b(18), b(17) => b(17), 
                           b(16) => b(16), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           s(31) => s(31), s(30) => s(30), s(29) => s(29), 
                           s(28) => s(28), s(27) => s(27), s(26) => s(26), 
                           s(25) => s(25), s(24) => s(24), s(23) => s(23), 
                           s(22) => s(22), s(21) => s(21), s(20) => s(20), 
                           s(19) => s(19), s(18) => s(18), s(17) => s(17), 
                           s(16) => s(16), s(15) => s(15), s(14) => s(14), 
                           s(13) => s(13), s(12) => s(12), s(11) => s(11), 
                           s(10) => s(10), s(9) => s(9), s(8) => s(8), s(7) => 
                           s(7), s(6) => s(6), s(5) => s(5), s(4) => s(4), s(3)
                           => s(3), s(2) => s(2), s(1) => s(1), s(0) => s(0), 
                           cout => cout);

end SYN_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Adder_DATA_SIZE32_1 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end Adder_DATA_SIZE32_1;

architecture SYN_adder_arch of Adder_DATA_SIZE32_1 is

   component P4Adder_DATA_SIZE32_SPARSITY4_1
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;

begin
   
   ADDER0 : P4Adder_DATA_SIZE32_SPARSITY4_1 port map( cin => cin, a(31) => 
                           a(31), a(30) => a(30), a(29) => a(29), a(28) => 
                           a(28), a(27) => a(27), a(26) => a(26), a(25) => 
                           a(25), a(24) => a(24), a(23) => a(23), a(22) => 
                           a(22), a(21) => a(21), a(20) => a(20), a(19) => 
                           a(19), a(18) => a(18), a(17) => a(17), a(16) => 
                           a(16), a(15) => a(15), a(14) => a(14), a(13) => 
                           a(13), a(12) => a(12), a(11) => a(11), a(10) => 
                           a(10), a(9) => a(9), a(8) => a(8), a(7) => a(7), 
                           a(6) => a(6), a(5) => a(5), a(4) => a(4), a(3) => 
                           a(3), a(2) => a(2), a(1) => a(1), a(0) => a(0), 
                           b(31) => b(31), b(30) => b(30), b(29) => b(29), 
                           b(28) => b(28), b(27) => b(27), b(26) => b(26), 
                           b(25) => b(25), b(24) => b(24), b(23) => b(23), 
                           b(22) => b(22), b(21) => b(21), b(20) => b(20), 
                           b(19) => b(19), b(18) => b(18), b(17) => b(17), 
                           b(16) => b(16), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           s(31) => s(31), s(30) => s(30), s(29) => s(29), 
                           s(28) => s(28), s(27) => s(27), s(26) => s(26), 
                           s(25) => s(25), s(24) => s(24), s(23) => s(23), 
                           s(22) => s(22), s(21) => s(21), s(20) => s(20), 
                           s(19) => s(19), s(18) => s(18), s(17) => s(17), 
                           s(16) => s(16), s(15) => s(15), s(14) => s(14), 
                           s(13) => s(13), s(12) => s(12), s(11) => s(11), 
                           s(10) => s(10), s(9) => s(9), s(8) => s(8), s(7) => 
                           s(7), s(6) => s(6), s(5) => s(5), s(4) => s(4), s(3)
                           => s(3), s(2) => s(2), s(1) => s(1), s(0) => s(0), 
                           cout => cout);

end SYN_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FullAdder_0 is

   port( ci, a, b : in std_logic;  s, co : out std_logic);

end FullAdder_0;

architecture SYN_full_adder_arch of FullAdder_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => b, B => n1, Z => s);
   U2 : INV_X1 port map( A => n2, ZN => co);
   U3 : AOI22_X1 port map( A1 => ci, A2 => a, B1 => n1, B2 => b, ZN => n2);
   U4 : XOR2_X1 port map( A => a, B => ci, Z => n1);

end SYN_full_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderSumGenerator_DATA_SIZE64_SPARSITY4 is

   port( a, b : in std_logic_vector (63 downto 0);  cin : in std_logic_vector 
         (15 downto 0);  sum : out std_logic_vector (63 downto 0));

end AdderSumGenerator_DATA_SIZE64_SPARSITY4;

architecture SYN_adder_sum_generator_arch of 
   AdderSumGenerator_DATA_SIZE64_SPARSITY4 is

   component AdderCarrySelect_DATA_SIZE4_17
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_18
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_19
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_20
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_21
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_22
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_23
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_24
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_25
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_26
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_27
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_28
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_29
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_30
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_31
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_32
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;

begin
   
   ACSi_0 : AdderCarrySelect_DATA_SIZE4_32 port map( a(3) => a(3), a(2) => a(2)
                           , a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), sel => cin(0), 
                           sum(3) => sum(3), sum(2) => sum(2), sum(1) => sum(1)
                           , sum(0) => sum(0));
   ACSi_1 : AdderCarrySelect_DATA_SIZE4_31 port map( a(3) => a(7), a(2) => a(6)
                           , a(1) => a(5), a(0) => a(4), b(3) => b(7), b(2) => 
                           b(6), b(1) => b(5), b(0) => b(4), sel => cin(1), 
                           sum(3) => sum(7), sum(2) => sum(6), sum(1) => sum(5)
                           , sum(0) => sum(4));
   ACSi_2 : AdderCarrySelect_DATA_SIZE4_30 port map( a(3) => a(11), a(2) => 
                           a(10), a(1) => a(9), a(0) => a(8), b(3) => b(11), 
                           b(2) => b(10), b(1) => b(9), b(0) => b(8), sel => 
                           cin(2), sum(3) => sum(11), sum(2) => sum(10), sum(1)
                           => sum(9), sum(0) => sum(8));
   ACSi_3 : AdderCarrySelect_DATA_SIZE4_29 port map( a(3) => a(15), a(2) => 
                           a(14), a(1) => a(13), a(0) => a(12), b(3) => b(15), 
                           b(2) => b(14), b(1) => b(13), b(0) => b(12), sel => 
                           cin(3), sum(3) => sum(15), sum(2) => sum(14), sum(1)
                           => sum(13), sum(0) => sum(12));
   ACSi_4 : AdderCarrySelect_DATA_SIZE4_28 port map( a(3) => a(19), a(2) => 
                           a(18), a(1) => a(17), a(0) => a(16), b(3) => b(19), 
                           b(2) => b(18), b(1) => b(17), b(0) => b(16), sel => 
                           cin(4), sum(3) => sum(19), sum(2) => sum(18), sum(1)
                           => sum(17), sum(0) => sum(16));
   ACSi_5 : AdderCarrySelect_DATA_SIZE4_27 port map( a(3) => a(23), a(2) => 
                           a(22), a(1) => a(21), a(0) => a(20), b(3) => b(23), 
                           b(2) => b(22), b(1) => b(21), b(0) => b(20), sel => 
                           cin(5), sum(3) => sum(23), sum(2) => sum(22), sum(1)
                           => sum(21), sum(0) => sum(20));
   ACSi_6 : AdderCarrySelect_DATA_SIZE4_26 port map( a(3) => a(27), a(2) => 
                           a(26), a(1) => a(25), a(0) => a(24), b(3) => b(27), 
                           b(2) => b(26), b(1) => b(25), b(0) => b(24), sel => 
                           cin(6), sum(3) => sum(27), sum(2) => sum(26), sum(1)
                           => sum(25), sum(0) => sum(24));
   ACSi_7 : AdderCarrySelect_DATA_SIZE4_25 port map( a(3) => a(31), a(2) => 
                           a(30), a(1) => a(29), a(0) => a(28), b(3) => b(31), 
                           b(2) => b(30), b(1) => b(29), b(0) => b(28), sel => 
                           cin(7), sum(3) => sum(31), sum(2) => sum(30), sum(1)
                           => sum(29), sum(0) => sum(28));
   ACSi_8 : AdderCarrySelect_DATA_SIZE4_24 port map( a(3) => a(35), a(2) => 
                           a(34), a(1) => a(33), a(0) => a(32), b(3) => b(35), 
                           b(2) => b(34), b(1) => b(33), b(0) => b(32), sel => 
                           cin(8), sum(3) => sum(35), sum(2) => sum(34), sum(1)
                           => sum(33), sum(0) => sum(32));
   ACSi_9 : AdderCarrySelect_DATA_SIZE4_23 port map( a(3) => a(39), a(2) => 
                           a(38), a(1) => a(37), a(0) => a(36), b(3) => b(39), 
                           b(2) => b(38), b(1) => b(37), b(0) => b(36), sel => 
                           cin(9), sum(3) => sum(39), sum(2) => sum(38), sum(1)
                           => sum(37), sum(0) => sum(36));
   ACSi_10 : AdderCarrySelect_DATA_SIZE4_22 port map( a(3) => a(43), a(2) => 
                           a(42), a(1) => a(41), a(0) => a(40), b(3) => b(43), 
                           b(2) => b(42), b(1) => b(41), b(0) => b(40), sel => 
                           cin(10), sum(3) => sum(43), sum(2) => sum(42), 
                           sum(1) => sum(41), sum(0) => sum(40));
   ACSi_11 : AdderCarrySelect_DATA_SIZE4_21 port map( a(3) => a(47), a(2) => 
                           a(46), a(1) => a(45), a(0) => a(44), b(3) => b(47), 
                           b(2) => b(46), b(1) => b(45), b(0) => b(44), sel => 
                           cin(11), sum(3) => sum(47), sum(2) => sum(46), 
                           sum(1) => sum(45), sum(0) => sum(44));
   ACSi_12 : AdderCarrySelect_DATA_SIZE4_20 port map( a(3) => a(51), a(2) => 
                           a(50), a(1) => a(49), a(0) => a(48), b(3) => b(51), 
                           b(2) => b(50), b(1) => b(49), b(0) => b(48), sel => 
                           cin(12), sum(3) => sum(51), sum(2) => sum(50), 
                           sum(1) => sum(49), sum(0) => sum(48));
   ACSi_13 : AdderCarrySelect_DATA_SIZE4_19 port map( a(3) => a(55), a(2) => 
                           a(54), a(1) => a(53), a(0) => a(52), b(3) => b(55), 
                           b(2) => b(54), b(1) => b(53), b(0) => b(52), sel => 
                           cin(13), sum(3) => sum(55), sum(2) => sum(54), 
                           sum(1) => sum(53), sum(0) => sum(52));
   ACSi_14 : AdderCarrySelect_DATA_SIZE4_18 port map( a(3) => a(59), a(2) => 
                           a(58), a(1) => a(57), a(0) => a(56), b(3) => b(59), 
                           b(2) => b(58), b(1) => b(57), b(0) => b(56), sel => 
                           cin(14), sum(3) => sum(59), sum(2) => sum(58), 
                           sum(1) => sum(57), sum(0) => sum(56));
   ACSi_15 : AdderCarrySelect_DATA_SIZE4_17 port map( a(3) => a(63), a(2) => 
                           a(62), a(1) => a(61), a(0) => a(60), b(3) => b(63), 
                           b(2) => b(62), b(1) => b(61), b(0) => b(60), sel => 
                           cin(15), sum(3) => sum(63), sum(2) => sum(62), 
                           sum(1) => sum(61), sum(0) => sum(60));

end SYN_adder_sum_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4CarryGenerator_DATA_SIZE64_SPARSITY4 is

   port( a, b : in std_logic_vector (63 downto 0);  cin : in std_logic;  cout :
         out std_logic_vector (15 downto 0));

end P4CarryGenerator_DATA_SIZE64_SPARSITY4;

architecture SYN_p4_carry_generator_arch of 
   P4CarryGenerator_DATA_SIZE64_SPARSITY4 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal cout_15_port, cout_14_port, cout_13_port, cout_12_port, cout_11_port,
      cout_10_port, cout_9_port, cout_8_port, cout_7_port, cout_6_port, 
      cout_5_port, cout_4_port, cout_3_port, cout_2_port, cout_1_port, 
      cout_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      n210, n211, n212, n213, n214, n215, n216 : std_logic;

begin
   cout <= ( cout_15_port, cout_14_port, cout_13_port, cout_12_port, 
      cout_11_port, cout_10_port, cout_9_port, cout_8_port, cout_7_port, 
      cout_6_port, cout_5_port, cout_4_port, cout_3_port, cout_2_port, 
      cout_1_port, cout_0_port );
   
   U1 : OAI21_X1 port map( B1 => n1, B2 => n2, A => n3, ZN => cout_9_port);
   U2 : OAI21_X1 port map( B1 => n4, B2 => n2, A => n5, ZN => cout_8_port);
   U3 : INV_X1 port map( A => n2, ZN => cout_7_port);
   U4 : OAI22_X1 port map( A1 => n6, A2 => n7, B1 => n8, B2 => n9, ZN => 
                           cout_15_port);
   U5 : AOI22_X1 port map( A1 => b(62), A2 => n10, B1 => a(62), B2 => n11, ZN 
                           => n9);
   U6 : OR2_X1 port map( A1 => n11, A2 => a(62), ZN => n10);
   U7 : OAI21_X1 port map( B1 => n12, B2 => n13, A => n14, ZN => n11);
   U8 : OAI21_X1 port map( B1 => b(61), B2 => a(61), A => n15, ZN => n14);
   U9 : INV_X1 port map( A => n16, ZN => n15);
   U10 : AOI21_X1 port map( B1 => cout_14_port, B2 => a(60), A => n17, ZN => 
                           n16);
   U11 : INV_X1 port map( A => n18, ZN => n17);
   U12 : OAI21_X1 port map( B1 => a(60), B2 => cout_14_port, A => b(60), ZN => 
                           n18);
   U13 : INV_X1 port map( A => b(61), ZN => n13);
   U14 : INV_X1 port map( A => a(61), ZN => n12);
   U15 : NOR2_X1 port map( A1 => b(63), A2 => a(63), ZN => n8);
   U16 : INV_X1 port map( A => b(63), ZN => n7);
   U17 : INV_X1 port map( A => a(63), ZN => n6);
   U18 : OAI21_X1 port map( B1 => n19, B2 => n20, A => n21, ZN => cout_14_port)
                           ;
   U19 : OAI21_X1 port map( B1 => a(59), B2 => n22, A => b(59), ZN => n21);
   U20 : INV_X1 port map( A => n19, ZN => n22);
   U21 : INV_X1 port map( A => a(59), ZN => n20);
   U22 : AOI21_X1 port map( B1 => a(58), B2 => b(58), A => n23, ZN => n19);
   U23 : INV_X1 port map( A => n24, ZN => n23);
   U24 : OAI22_X1 port map( A1 => n25, A2 => n26, B1 => a(58), B2 => b(58), ZN 
                           => n24);
   U25 : NOR2_X1 port map( A1 => n27, A2 => n28, ZN => n26);
   U26 : AOI22_X1 port map( A1 => n27, A2 => n28, B1 => n29, B2 => n30, ZN => 
                           n25);
   U27 : OAI21_X1 port map( B1 => a(56), B2 => cout_13_port, A => b(56), ZN => 
                           n30);
   U28 : NAND2_X1 port map( A1 => a(56), A2 => cout_13_port, ZN => n29);
   U29 : INV_X1 port map( A => b(57), ZN => n28);
   U30 : INV_X1 port map( A => a(57), ZN => n27);
   U31 : OAI22_X1 port map( A1 => n31, A2 => n32, B1 => n33, B2 => n34, ZN => 
                           cout_13_port);
   U32 : AOI22_X1 port map( A1 => b(54), A2 => n35, B1 => a(54), B2 => n36, ZN 
                           => n34);
   U33 : OR2_X1 port map( A1 => n36, A2 => a(54), ZN => n35);
   U34 : OAI21_X1 port map( B1 => n37, B2 => n38, A => n39, ZN => n36);
   U35 : OAI21_X1 port map( B1 => b(53), B2 => a(53), A => n40, ZN => n39);
   U36 : OAI21_X1 port map( B1 => n41, B2 => n42, A => n43, ZN => n40);
   U37 : OAI21_X1 port map( B1 => a(52), B2 => cout_12_port, A => b(52), ZN => 
                           n43);
   U38 : INV_X1 port map( A => a(52), ZN => n42);
   U39 : INV_X1 port map( A => cout_12_port, ZN => n41);
   U40 : INV_X1 port map( A => b(53), ZN => n38);
   U41 : INV_X1 port map( A => a(53), ZN => n37);
   U42 : NOR2_X1 port map( A1 => b(55), A2 => a(55), ZN => n33);
   U43 : INV_X1 port map( A => b(55), ZN => n32);
   U44 : INV_X1 port map( A => a(55), ZN => n31);
   U45 : OAI211_X1 port map( C1 => n44, C2 => n45, A => n46, B => n47, ZN => 
                           cout_12_port);
   U46 : OAI211_X1 port map( C1 => b(51), C2 => a(51), A => cout_11_port, B => 
                           n48, ZN => n47);
   U47 : AOI221_X1 port map( B1 => n49, B2 => n50, C1 => n51, C2 => n52, A => 
                           n53, ZN => n48);
   U48 : OAI21_X1 port map( B1 => n54, B2 => a(51), A => b(51), ZN => n46);
   U49 : INV_X1 port map( A => a(51), ZN => n45);
   U50 : INV_X1 port map( A => n54, ZN => n44);
   U51 : AOI21_X1 port map( B1 => n49, B2 => n55, A => n56, ZN => n54);
   U52 : INV_X1 port map( A => n57, ZN => n56);
   U53 : OAI21_X1 port map( B1 => n55, B2 => n49, A => n50, ZN => n57);
   U54 : INV_X1 port map( A => b(50), ZN => n50);
   U55 : AOI21_X1 port map( B1 => a(49), B2 => b(49), A => n58, ZN => n55);
   U56 : NOR3_X1 port map( A1 => n51, A2 => n53, A3 => n52, ZN => n58);
   U57 : INV_X1 port map( A => b(48), ZN => n52);
   U58 : NOR2_X1 port map( A1 => b(49), A2 => a(49), ZN => n53);
   U59 : INV_X1 port map( A => a(48), ZN => n51);
   U60 : INV_X1 port map( A => a(50), ZN => n49);
   U61 : INV_X1 port map( A => n59, ZN => cout_11_port);
   U62 : OAI22_X1 port map( A1 => a(47), A2 => n60, B1 => b(47), B2 => n61, ZN 
                           => n59);
   U63 : AND2_X1 port map( A1 => n60, A2 => a(47), ZN => n61);
   U64 : INV_X1 port map( A => n62, ZN => n60);
   U65 : OAI22_X1 port map( A1 => a(46), A2 => n63, B1 => b(46), B2 => n64, ZN 
                           => n62);
   U66 : AND2_X1 port map( A1 => n63, A2 => a(46), ZN => n64);
   U67 : OAI21_X1 port map( B1 => n65, B2 => n66, A => n67, ZN => n63);
   U68 : OAI21_X1 port map( B1 => a(45), B2 => b(45), A => n68, ZN => n67);
   U69 : OAI21_X1 port map( B1 => n69, B2 => n70, A => n71, ZN => n68);
   U70 : OAI21_X1 port map( B1 => a(44), B2 => cout_10_port, A => b(44), ZN => 
                           n71);
   U71 : INV_X1 port map( A => a(44), ZN => n70);
   U72 : INV_X1 port map( A => cout_10_port, ZN => n69);
   U73 : INV_X1 port map( A => b(45), ZN => n66);
   U74 : INV_X1 port map( A => a(45), ZN => n65);
   U75 : OAI211_X1 port map( C1 => n72, C2 => n73, A => n74, B => n75, ZN => 
                           cout_10_port);
   U76 : OAI221_X1 port map( B1 => b(43), B2 => a(43), C1 => n76, C2 => n77, A 
                           => n78, ZN => n75);
   U77 : AOI221_X1 port map( B1 => n79, B2 => n80, C1 => n81, C2 => n82, A => 
                           n83, ZN => n78);
   U78 : INV_X1 port map( A => n3, ZN => n77);
   U79 : OAI22_X1 port map( A1 => a(39), A2 => n84, B1 => b(39), B2 => n85, ZN 
                           => n3);
   U80 : AND2_X1 port map( A1 => n84, A2 => a(39), ZN => n85);
   U81 : AOI21_X1 port map( B1 => n86, B2 => n87, A => n88, ZN => n84);
   U82 : AOI21_X1 port map( B1 => n89, B2 => a(38), A => b(38), ZN => n88);
   U83 : INV_X1 port map( A => n87, ZN => n89);
   U84 : AOI21_X1 port map( B1 => n90, B2 => a(37), A => n91, ZN => n87);
   U85 : INV_X1 port map( A => n92, ZN => n91);
   U86 : OAI21_X1 port map( B1 => n90, B2 => a(37), A => b(37), ZN => n92);
   U87 : AOI21_X1 port map( B1 => n93, B2 => n5, A => n94, ZN => n90);
   U88 : AOI21_X1 port map( B1 => n95, B2 => a(36), A => b(36), ZN => n94);
   U89 : INV_X1 port map( A => n95, ZN => n5);
   U90 : AOI21_X1 port map( B1 => n96, B2 => n97, A => n98, ZN => n95);
   U91 : AOI21_X1 port map( B1 => n99, B2 => a(35), A => b(35), ZN => n98);
   U92 : INV_X1 port map( A => n97, ZN => n99);
   U93 : OAI21_X1 port map( B1 => a(34), B2 => n100, A => n101, ZN => n97);
   U94 : INV_X1 port map( A => n102, ZN => n101);
   U95 : AOI21_X1 port map( B1 => n100, B2 => a(34), A => b(34), ZN => n102);
   U96 : OAI21_X1 port map( B1 => n103, B2 => n104, A => n105, ZN => n100);
   U97 : NAND3_X1 port map( A1 => a(32), A2 => n106, A3 => b(32), ZN => n105);
   U98 : INV_X1 port map( A => a(35), ZN => n96);
   U99 : INV_X1 port map( A => a(36), ZN => n93);
   U100 : INV_X1 port map( A => a(38), ZN => n86);
   U101 : NOR2_X1 port map( A1 => n1, A2 => n2, ZN => n76);
   U102 : OAI22_X1 port map( A1 => a(31), A2 => n107, B1 => b(31), B2 => n108, 
                           ZN => n2);
   U103 : AND2_X1 port map( A1 => n107, A2 => a(31), ZN => n108);
   U104 : INV_X1 port map( A => n109, ZN => n107);
   U105 : OAI22_X1 port map( A1 => a(30), A2 => n110, B1 => b(30), B2 => n111, 
                           ZN => n109);
   U106 : AND2_X1 port map( A1 => n110, A2 => a(30), ZN => n111);
   U107 : OAI21_X1 port map( B1 => n112, B2 => n113, A => n114, ZN => n110);
   U108 : OAI21_X1 port map( B1 => b(29), B2 => a(29), A => n115, ZN => n114);
   U109 : INV_X1 port map( A => n116, ZN => n115);
   U110 : AOI21_X1 port map( B1 => cout_6_port, B2 => a(28), A => n117, ZN => 
                           n116);
   U111 : INV_X1 port map( A => n118, ZN => n117);
   U112 : OAI21_X1 port map( B1 => a(28), B2 => cout_6_port, A => b(28), ZN => 
                           n118);
   U113 : OAI21_X1 port map( B1 => n119, B2 => n120, A => n121, ZN => 
                           cout_6_port);
   U114 : OAI21_X1 port map( B1 => a(27), B2 => n122, A => b(27), ZN => n121);
   U115 : INV_X1 port map( A => n119, ZN => n122);
   U116 : INV_X1 port map( A => a(27), ZN => n120);
   U117 : AOI21_X1 port map( B1 => a(26), B2 => b(26), A => n123, ZN => n119);
   U118 : INV_X1 port map( A => n124, ZN => n123);
   U119 : OAI22_X1 port map( A1 => n125, A2 => n126, B1 => a(26), B2 => b(26), 
                           ZN => n124);
   U120 : NOR2_X1 port map( A1 => n127, A2 => n128, ZN => n126);
   U121 : AOI22_X1 port map( A1 => n127, A2 => n128, B1 => n129, B2 => n130, ZN
                           => n125);
   U122 : OAI21_X1 port map( B1 => a(24), B2 => cout_5_port, A => b(24), ZN => 
                           n130);
   U123 : NAND2_X1 port map( A1 => a(24), A2 => cout_5_port, ZN => n129);
   U124 : OAI22_X1 port map( A1 => n131, A2 => n132, B1 => n133, B2 => n134, ZN
                           => cout_5_port);
   U125 : AOI22_X1 port map( A1 => b(22), A2 => n135, B1 => a(22), B2 => n136, 
                           ZN => n134);
   U126 : OR2_X1 port map( A1 => n136, A2 => a(22), ZN => n135);
   U127 : OAI21_X1 port map( B1 => n137, B2 => n138, A => n139, ZN => n136);
   U128 : OAI21_X1 port map( B1 => b(21), B2 => a(21), A => n140, ZN => n139);
   U129 : OAI21_X1 port map( B1 => n141, B2 => n142, A => n143, ZN => n140);
   U130 : OAI21_X1 port map( B1 => a(20), B2 => cout_4_port, A => b(20), ZN => 
                           n143);
   U131 : INV_X1 port map( A => a(20), ZN => n142);
   U132 : INV_X1 port map( A => cout_4_port, ZN => n141);
   U133 : OAI211_X1 port map( C1 => n144, C2 => n145, A => n146, B => n147, ZN 
                           => cout_4_port);
   U134 : OAI21_X1 port map( B1 => n148, B2 => a(19), A => b(19), ZN => n147);
   U135 : OAI211_X1 port map( C1 => b(19), C2 => a(19), A => cout_3_port, B => 
                           n149, ZN => n146);
   U136 : AOI221_X1 port map( B1 => n150, B2 => n151, C1 => n152, C2 => n153, A
                           => n154, ZN => n149);
   U137 : INV_X1 port map( A => n155, ZN => cout_3_port);
   U138 : OAI22_X1 port map( A1 => a(15), A2 => n156, B1 => b(15), B2 => n157, 
                           ZN => n155);
   U139 : AND2_X1 port map( A1 => n156, A2 => a(15), ZN => n157);
   U140 : INV_X1 port map( A => n158, ZN => n156);
   U141 : OAI22_X1 port map( A1 => a(14), A2 => n159, B1 => b(14), B2 => n160, 
                           ZN => n158);
   U142 : AND2_X1 port map( A1 => n159, A2 => a(14), ZN => n160);
   U143 : OAI21_X1 port map( B1 => n161, B2 => n162, A => n163, ZN => n159);
   U144 : OAI21_X1 port map( B1 => b(13), B2 => a(13), A => n164, ZN => n163);
   U145 : INV_X1 port map( A => n165, ZN => n164);
   U146 : AOI21_X1 port map( B1 => cout_2_port, B2 => a(12), A => n166, ZN => 
                           n165);
   U147 : INV_X1 port map( A => n167, ZN => n166);
   U148 : OAI21_X1 port map( B1 => a(12), B2 => cout_2_port, A => b(12), ZN => 
                           n167);
   U149 : OAI21_X1 port map( B1 => n168, B2 => n169, A => n170, ZN => 
                           cout_2_port);
   U150 : OAI21_X1 port map( B1 => a(11), B2 => n171, A => b(11), ZN => n170);
   U151 : INV_X1 port map( A => n168, ZN => n171);
   U152 : INV_X1 port map( A => a(11), ZN => n169);
   U153 : AOI21_X1 port map( B1 => a(10), B2 => b(10), A => n172, ZN => n168);
   U154 : INV_X1 port map( A => n173, ZN => n172);
   U155 : OAI22_X1 port map( A1 => n174, A2 => n175, B1 => a(10), B2 => b(10), 
                           ZN => n173);
   U156 : NOR2_X1 port map( A1 => n176, A2 => n177, ZN => n175);
   U157 : AOI22_X1 port map( A1 => n176, A2 => n177, B1 => n178, B2 => n179, ZN
                           => n174);
   U158 : OAI21_X1 port map( B1 => a(8), B2 => cout_1_port, A => b(8), ZN => 
                           n179);
   U159 : NAND2_X1 port map( A1 => a(8), A2 => cout_1_port, ZN => n178);
   U160 : OAI21_X1 port map( B1 => n180, B2 => n181, A => n182, ZN => 
                           cout_1_port);
   U161 : OAI21_X1 port map( B1 => b(7), B2 => a(7), A => n183, ZN => n182);
   U162 : OAI21_X1 port map( B1 => n184, B2 => n185, A => n186, ZN => n183);
   U163 : OAI21_X1 port map( B1 => a(6), B2 => n187, A => b(6), ZN => n186);
   U164 : INV_X1 port map( A => n184, ZN => n187);
   U165 : INV_X1 port map( A => a(6), ZN => n185);
   U166 : AOI22_X1 port map( A1 => a(5), A2 => b(5), B1 => n188, B2 => n189, ZN
                           => n184);
   U167 : INV_X1 port map( A => n190, ZN => n189);
   U168 : AOI22_X1 port map( A1 => b(4), A2 => n191, B1 => a(4), B2 => 
                           cout_0_port, ZN => n190);
   U169 : OR2_X1 port map( A1 => a(4), A2 => cout_0_port, ZN => n191);
   U170 : OR2_X1 port map( A1 => b(5), A2 => a(5), ZN => n188);
   U171 : INV_X1 port map( A => b(7), ZN => n181);
   U172 : INV_X1 port map( A => a(7), ZN => n180);
   U173 : INV_X1 port map( A => b(9), ZN => n177);
   U174 : INV_X1 port map( A => a(9), ZN => n176);
   U175 : INV_X1 port map( A => b(13), ZN => n162);
   U176 : INV_X1 port map( A => a(13), ZN => n161);
   U177 : INV_X1 port map( A => a(19), ZN => n145);
   U178 : INV_X1 port map( A => n148, ZN => n144);
   U179 : AOI21_X1 port map( B1 => n150, B2 => n192, A => n193, ZN => n148);
   U180 : INV_X1 port map( A => n194, ZN => n193);
   U181 : OAI21_X1 port map( B1 => n192, B2 => n150, A => n151, ZN => n194);
   U182 : INV_X1 port map( A => b(18), ZN => n151);
   U183 : AOI21_X1 port map( B1 => a(17), B2 => b(17), A => n195, ZN => n192);
   U184 : NOR3_X1 port map( A1 => n152, A2 => n154, A3 => n153, ZN => n195);
   U185 : INV_X1 port map( A => b(16), ZN => n153);
   U186 : NOR2_X1 port map( A1 => b(17), A2 => a(17), ZN => n154);
   U187 : INV_X1 port map( A => a(16), ZN => n152);
   U188 : INV_X1 port map( A => a(18), ZN => n150);
   U189 : INV_X1 port map( A => b(21), ZN => n138);
   U190 : INV_X1 port map( A => a(21), ZN => n137);
   U191 : NOR2_X1 port map( A1 => b(23), A2 => a(23), ZN => n133);
   U192 : INV_X1 port map( A => b(23), ZN => n132);
   U193 : INV_X1 port map( A => a(23), ZN => n131);
   U194 : INV_X1 port map( A => b(25), ZN => n128);
   U195 : INV_X1 port map( A => a(25), ZN => n127);
   U196 : INV_X1 port map( A => b(29), ZN => n113);
   U197 : INV_X1 port map( A => a(29), ZN => n112);
   U198 : OAI211_X1 port map( C1 => b(39), C2 => a(39), A => n196, B => n197, 
                           ZN => n1);
   U199 : INV_X1 port map( A => n198, ZN => n197);
   U200 : OAI222_X1 port map( A1 => a(38), A2 => b(38), B1 => a(36), B2 => 
                           b(36), C1 => a(37), C2 => b(37), ZN => n198);
   U201 : INV_X1 port map( A => n4, ZN => n196);
   U202 : OAI211_X1 port map( C1 => b(32), C2 => a(32), A => n106, B => n199, 
                           ZN => n4);
   U203 : INV_X1 port map( A => n200, ZN => n199);
   U204 : OAI22_X1 port map( A1 => a(34), A2 => b(34), B1 => a(35), B2 => b(35)
                           , ZN => n200);
   U205 : NAND2_X1 port map( A1 => n104, A2 => n103, ZN => n106);
   U206 : INV_X1 port map( A => a(33), ZN => n103);
   U207 : INV_X1 port map( A => b(33), ZN => n104);
   U208 : OAI21_X1 port map( B1 => n201, B2 => a(43), A => b(43), ZN => n74);
   U209 : INV_X1 port map( A => a(43), ZN => n73);
   U210 : INV_X1 port map( A => n201, ZN => n72);
   U211 : AOI21_X1 port map( B1 => n79, B2 => n202, A => n203, ZN => n201);
   U212 : INV_X1 port map( A => n204, ZN => n203);
   U213 : OAI21_X1 port map( B1 => n202, B2 => n79, A => n80, ZN => n204);
   U214 : INV_X1 port map( A => b(42), ZN => n80);
   U215 : AOI21_X1 port map( B1 => a(41), B2 => b(41), A => n205, ZN => n202);
   U216 : NOR3_X1 port map( A1 => n81, A2 => n83, A3 => n82, ZN => n205);
   U217 : INV_X1 port map( A => b(40), ZN => n82);
   U218 : NOR2_X1 port map( A1 => b(41), A2 => a(41), ZN => n83);
   U219 : INV_X1 port map( A => a(40), ZN => n81);
   U220 : INV_X1 port map( A => a(42), ZN => n79);
   U221 : INV_X1 port map( A => n206, ZN => cout_0_port);
   U222 : OAI22_X1 port map( A1 => a(3), A2 => n207, B1 => b(3), B2 => n208, ZN
                           => n206);
   U223 : AND2_X1 port map( A1 => n207, A2 => a(3), ZN => n208);
   U224 : INV_X1 port map( A => n209, ZN => n207);
   U225 : OAI22_X1 port map( A1 => a(2), A2 => n210, B1 => b(2), B2 => n211, ZN
                           => n209);
   U226 : AND2_X1 port map( A1 => n210, A2 => a(2), ZN => n211);
   U227 : INV_X1 port map( A => n212, ZN => n210);
   U228 : AOI22_X1 port map( A1 => a(1), A2 => b(1), B1 => n213, B2 => n214, ZN
                           => n212);
   U229 : INV_X1 port map( A => n215, ZN => n214);
   U230 : AOI22_X1 port map( A1 => cin, A2 => n216, B1 => b(0), B2 => a(0), ZN 
                           => n215);
   U231 : OR2_X1 port map( A1 => b(0), A2 => a(0), ZN => n216);
   U232 : OR2_X1 port map( A1 => b(1), A2 => a(1), ZN => n213);

end SYN_p4_carry_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderSumGenerator_DATA_SIZE16_SPARSITY4 is

   port( a, b : in std_logic_vector (15 downto 0);  cin : in std_logic_vector 
         (3 downto 0);  sum : out std_logic_vector (15 downto 0));

end AdderSumGenerator_DATA_SIZE16_SPARSITY4;

architecture SYN_adder_sum_generator_arch of 
   AdderSumGenerator_DATA_SIZE16_SPARSITY4 is

   component AdderCarrySelect_DATA_SIZE4_57
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_58
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_59
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_60
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;

begin
   
   ACSi_0 : AdderCarrySelect_DATA_SIZE4_60 port map( a(3) => a(3), a(2) => a(2)
                           , a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), sel => cin(0), 
                           sum(3) => sum(3), sum(2) => sum(2), sum(1) => sum(1)
                           , sum(0) => sum(0));
   ACSi_1 : AdderCarrySelect_DATA_SIZE4_59 port map( a(3) => a(7), a(2) => a(6)
                           , a(1) => a(5), a(0) => a(4), b(3) => b(7), b(2) => 
                           b(6), b(1) => b(5), b(0) => b(4), sel => cin(1), 
                           sum(3) => sum(7), sum(2) => sum(6), sum(1) => sum(5)
                           , sum(0) => sum(4));
   ACSi_2 : AdderCarrySelect_DATA_SIZE4_58 port map( a(3) => a(11), a(2) => 
                           a(10), a(1) => a(9), a(0) => a(8), b(3) => b(11), 
                           b(2) => b(10), b(1) => b(9), b(0) => b(8), sel => 
                           cin(2), sum(3) => sum(11), sum(2) => sum(10), sum(1)
                           => sum(9), sum(0) => sum(8));
   ACSi_3 : AdderCarrySelect_DATA_SIZE4_57 port map( a(3) => a(15), a(2) => 
                           a(14), a(1) => a(13), a(0) => a(12), b(3) => b(15), 
                           b(2) => b(14), b(1) => b(13), b(0) => b(12), sel => 
                           cin(3), sum(3) => sum(15), sum(2) => sum(14), sum(1)
                           => sum(13), sum(0) => sum(12));

end SYN_adder_sum_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4CarryGenerator_DATA_SIZE16_SPARSITY4 is

   port( a, b : in std_logic_vector (15 downto 0);  cin : in std_logic;  cout :
         out std_logic_vector (3 downto 0));

end P4CarryGenerator_DATA_SIZE16_SPARSITY4;

architecture SYN_p4_carry_generator_arch of 
   P4CarryGenerator_DATA_SIZE16_SPARSITY4 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal cout_3_port, cout_2_port, cout_1_port, cout_0_port, n1, n2, n3, n4, 
      n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20
      , n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, 
      n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48 : 
      std_logic;

begin
   cout <= ( cout_3_port, cout_2_port, cout_1_port, cout_0_port );
   
   U1 : OAI22_X1 port map( A1 => n1, A2 => n2, B1 => n3, B2 => n4, ZN => 
                           cout_3_port);
   U2 : AOI22_X1 port map( A1 => b(14), A2 => n5, B1 => a(14), B2 => n6, ZN => 
                           n4);
   U3 : OR2_X1 port map( A1 => n6, A2 => a(14), ZN => n5);
   U4 : OAI21_X1 port map( B1 => n7, B2 => n8, A => n9, ZN => n6);
   U5 : OAI21_X1 port map( B1 => b(13), B2 => a(13), A => n10, ZN => n9);
   U6 : INV_X1 port map( A => n11, ZN => n10);
   U7 : AOI21_X1 port map( B1 => cout_2_port, B2 => a(12), A => n12, ZN => n11)
                           ;
   U8 : INV_X1 port map( A => n13, ZN => n12);
   U9 : OAI21_X1 port map( B1 => a(12), B2 => cout_2_port, A => b(12), ZN => 
                           n13);
   U10 : INV_X1 port map( A => b(13), ZN => n8);
   U11 : INV_X1 port map( A => a(13), ZN => n7);
   U12 : NOR2_X1 port map( A1 => b(15), A2 => a(15), ZN => n3);
   U13 : INV_X1 port map( A => b(15), ZN => n2);
   U14 : INV_X1 port map( A => a(15), ZN => n1);
   U15 : OAI21_X1 port map( B1 => n14, B2 => n15, A => n16, ZN => cout_2_port);
   U16 : OAI21_X1 port map( B1 => a(11), B2 => n17, A => b(11), ZN => n16);
   U17 : INV_X1 port map( A => n14, ZN => n17);
   U18 : INV_X1 port map( A => a(11), ZN => n15);
   U19 : AOI21_X1 port map( B1 => a(10), B2 => b(10), A => n18, ZN => n14);
   U20 : INV_X1 port map( A => n19, ZN => n18);
   U21 : OAI22_X1 port map( A1 => n20, A2 => n21, B1 => a(10), B2 => b(10), ZN 
                           => n19);
   U22 : NOR2_X1 port map( A1 => n22, A2 => n23, ZN => n21);
   U23 : AOI22_X1 port map( A1 => n22, A2 => n23, B1 => n24, B2 => n25, ZN => 
                           n20);
   U24 : OAI21_X1 port map( B1 => a(8), B2 => cout_1_port, A => b(8), ZN => n25
                           );
   U25 : NAND2_X1 port map( A1 => a(8), A2 => cout_1_port, ZN => n24);
   U26 : INV_X1 port map( A => b(9), ZN => n23);
   U27 : INV_X1 port map( A => a(9), ZN => n22);
   U28 : OAI21_X1 port map( B1 => n26, B2 => n27, A => n28, ZN => cout_1_port);
   U29 : OAI21_X1 port map( B1 => b(7), B2 => a(7), A => n29, ZN => n28);
   U30 : OAI21_X1 port map( B1 => n30, B2 => n31, A => n32, ZN => n29);
   U31 : OAI21_X1 port map( B1 => a(6), B2 => n33, A => b(6), ZN => n32);
   U32 : INV_X1 port map( A => n30, ZN => n33);
   U33 : INV_X1 port map( A => a(6), ZN => n31);
   U34 : AOI22_X1 port map( A1 => a(5), A2 => b(5), B1 => n34, B2 => n35, ZN =>
                           n30);
   U35 : INV_X1 port map( A => n36, ZN => n35);
   U36 : AOI22_X1 port map( A1 => b(4), A2 => n37, B1 => a(4), B2 => 
                           cout_0_port, ZN => n36);
   U37 : OR2_X1 port map( A1 => a(4), A2 => cout_0_port, ZN => n37);
   U38 : OR2_X1 port map( A1 => b(5), A2 => a(5), ZN => n34);
   U39 : INV_X1 port map( A => b(7), ZN => n27);
   U40 : INV_X1 port map( A => a(7), ZN => n26);
   U41 : INV_X1 port map( A => n38, ZN => cout_0_port);
   U42 : OAI22_X1 port map( A1 => a(3), A2 => n39, B1 => b(3), B2 => n40, ZN =>
                           n38);
   U43 : AND2_X1 port map( A1 => n39, A2 => a(3), ZN => n40);
   U44 : INV_X1 port map( A => n41, ZN => n39);
   U45 : OAI22_X1 port map( A1 => a(2), A2 => n42, B1 => b(2), B2 => n43, ZN =>
                           n41);
   U46 : AND2_X1 port map( A1 => n42, A2 => a(2), ZN => n43);
   U47 : INV_X1 port map( A => n44, ZN => n42);
   U48 : AOI22_X1 port map( A1 => a(1), A2 => b(1), B1 => n45, B2 => n46, ZN =>
                           n44);
   U49 : INV_X1 port map( A => n47, ZN => n46);
   U50 : AOI22_X1 port map( A1 => cin, A2 => n48, B1 => b(0), B2 => a(0), ZN =>
                           n47);
   U51 : OR2_X1 port map( A1 => b(0), A2 => a(0), ZN => n48);
   U52 : OR2_X1 port map( A1 => b(1), A2 => a(1), ZN => n45);

end SYN_p4_carry_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE4_0 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);  
         dout : out std_logic_vector (3 downto 0));

end Mux_DATA_SIZE4_0;

architecture SYN_mux_arch of Mux_DATA_SIZE4_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U2 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U3 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U4 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Rca_DATA_SIZE4_0 is

   port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : out 
         std_logic_vector (3 downto 0);  co : out std_logic);

end Rca_DATA_SIZE4_0;

architecture SYN_rca_arch of Rca_DATA_SIZE4_0 is

   component FullAdder_669
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_670
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_671
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   component FullAdder_0
      port( ci, a, b : in std_logic;  s, co : out std_logic);
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   FA1_0 : FullAdder_0 port map( ci => ci, a => a(0), b => b(0), s => s(0), co 
                           => carry_1_port);
   FA3_1 : FullAdder_671 port map( ci => carry_1_port, a => a(1), b => b(1), s 
                           => s(1), co => carry_2_port);
   FA3_2 : FullAdder_670 port map( ci => carry_2_port, a => a(2), b => b(2), s 
                           => s(2), co => carry_3_port);
   FA3_3 : FullAdder_669 port map( ci => carry_3_port, a => a(3), b => b(3), s 
                           => s(3), co => co);

end SYN_rca_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4Adder_DATA_SIZE64_SPARSITY4 is

   port( cin : in std_logic;  a, b : in std_logic_vector (63 downto 0);  s : 
         out std_logic_vector (63 downto 0);  cout : out std_logic);

end P4Adder_DATA_SIZE64_SPARSITY4;

architecture SYN_p4_adder_arch of P4Adder_DATA_SIZE64_SPARSITY4 is

   component AdderSumGenerator_DATA_SIZE64_SPARSITY4
      port( a, b : in std_logic_vector (63 downto 0);  cin : in 
            std_logic_vector (15 downto 0);  sum : out std_logic_vector (63 
            downto 0));
   end component;
   
   component P4CarryGenerator_DATA_SIZE64_SPARSITY4
      port( a, b : in std_logic_vector (63 downto 0);  cin : in std_logic;  
            cout : out std_logic_vector (15 downto 0));
   end component;
   
   signal carry_15_port, carry_14_port, carry_13_port, carry_12_port, 
      carry_11_port, carry_10_port, carry_9_port, carry_8_port, carry_7_port, 
      carry_6_port, carry_5_port, carry_4_port, carry_3_port, carry_2_port, 
      carry_1_port : std_logic;

begin
   
   CG0 : P4CarryGenerator_DATA_SIZE64_SPARSITY4 port map( a(63) => a(63), a(62)
                           => a(62), a(61) => a(61), a(60) => a(60), a(59) => 
                           a(59), a(58) => a(58), a(57) => a(57), a(56) => 
                           a(56), a(55) => a(55), a(54) => a(54), a(53) => 
                           a(53), a(52) => a(52), a(51) => a(51), a(50) => 
                           a(50), a(49) => a(49), a(48) => a(48), a(47) => 
                           a(47), a(46) => a(46), a(45) => a(45), a(44) => 
                           a(44), a(43) => a(43), a(42) => a(42), a(41) => 
                           a(41), a(40) => a(40), a(39) => a(39), a(38) => 
                           a(38), a(37) => a(37), a(36) => a(36), a(35) => 
                           a(35), a(34) => a(34), a(33) => a(33), a(32) => 
                           a(32), a(31) => a(31), a(30) => a(30), a(29) => 
                           a(29), a(28) => a(28), a(27) => a(27), a(26) => 
                           a(26), a(25) => a(25), a(24) => a(24), a(23) => 
                           a(23), a(22) => a(22), a(21) => a(21), a(20) => 
                           a(20), a(19) => a(19), a(18) => a(18), a(17) => 
                           a(17), a(16) => a(16), a(15) => a(15), a(14) => 
                           a(14), a(13) => a(13), a(12) => a(12), a(11) => 
                           a(11), a(10) => a(10), a(9) => a(9), a(8) => a(8), 
                           a(7) => a(7), a(6) => a(6), a(5) => a(5), a(4) => 
                           a(4), a(3) => a(3), a(2) => a(2), a(1) => a(1), a(0)
                           => a(0), b(63) => b(63), b(62) => b(62), b(61) => 
                           b(61), b(60) => b(60), b(59) => b(59), b(58) => 
                           b(58), b(57) => b(57), b(56) => b(56), b(55) => 
                           b(55), b(54) => b(54), b(53) => b(53), b(52) => 
                           b(52), b(51) => b(51), b(50) => b(50), b(49) => 
                           b(49), b(48) => b(48), b(47) => b(47), b(46) => 
                           b(46), b(45) => b(45), b(44) => b(44), b(43) => 
                           b(43), b(42) => b(42), b(41) => b(41), b(40) => 
                           b(40), b(39) => b(39), b(38) => b(38), b(37) => 
                           b(37), b(36) => b(36), b(35) => b(35), b(34) => 
                           b(34), b(33) => b(33), b(32) => b(32), b(31) => 
                           b(31), b(30) => b(30), b(29) => b(29), b(28) => 
                           b(28), b(27) => b(27), b(26) => b(26), b(25) => 
                           b(25), b(24) => b(24), b(23) => b(23), b(22) => 
                           b(22), b(21) => b(21), b(20) => b(20), b(19) => 
                           b(19), b(18) => b(18), b(17) => b(17), b(16) => 
                           b(16), b(15) => b(15), b(14) => b(14), b(13) => 
                           b(13), b(12) => b(12), b(11) => b(11), b(10) => 
                           b(10), b(9) => b(9), b(8) => b(8), b(7) => b(7), 
                           b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3) => 
                           b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), cin 
                           => cin, cout(15) => cout, cout(14) => carry_15_port,
                           cout(13) => carry_14_port, cout(12) => carry_13_port
                           , cout(11) => carry_12_port, cout(10) => 
                           carry_11_port, cout(9) => carry_10_port, cout(8) => 
                           carry_9_port, cout(7) => carry_8_port, cout(6) => 
                           carry_7_port, cout(5) => carry_6_port, cout(4) => 
                           carry_5_port, cout(3) => carry_4_port, cout(2) => 
                           carry_3_port, cout(1) => carry_2_port, cout(0) => 
                           carry_1_port);
   SG0 : AdderSumGenerator_DATA_SIZE64_SPARSITY4 port map( a(63) => a(63), 
                           a(62) => a(62), a(61) => a(61), a(60) => a(60), 
                           a(59) => a(59), a(58) => a(58), a(57) => a(57), 
                           a(56) => a(56), a(55) => a(55), a(54) => a(54), 
                           a(53) => a(53), a(52) => a(52), a(51) => a(51), 
                           a(50) => a(50), a(49) => a(49), a(48) => a(48), 
                           a(47) => a(47), a(46) => a(46), a(45) => a(45), 
                           a(44) => a(44), a(43) => a(43), a(42) => a(42), 
                           a(41) => a(41), a(40) => a(40), a(39) => a(39), 
                           a(38) => a(38), a(37) => a(37), a(36) => a(36), 
                           a(35) => a(35), a(34) => a(34), a(33) => a(33), 
                           a(32) => a(32), a(31) => a(31), a(30) => a(30), 
                           a(29) => a(29), a(28) => a(28), a(27) => a(27), 
                           a(26) => a(26), a(25) => a(25), a(24) => a(24), 
                           a(23) => a(23), a(22) => a(22), a(21) => a(21), 
                           a(20) => a(20), a(19) => a(19), a(18) => a(18), 
                           a(17) => a(17), a(16) => a(16), a(15) => a(15), 
                           a(14) => a(14), a(13) => a(13), a(12) => a(12), 
                           a(11) => a(11), a(10) => a(10), a(9) => a(9), a(8) 
                           => a(8), a(7) => a(7), a(6) => a(6), a(5) => a(5), 
                           a(4) => a(4), a(3) => a(3), a(2) => a(2), a(1) => 
                           a(1), a(0) => a(0), b(63) => b(63), b(62) => b(62), 
                           b(61) => b(61), b(60) => b(60), b(59) => b(59), 
                           b(58) => b(58), b(57) => b(57), b(56) => b(56), 
                           b(55) => b(55), b(54) => b(54), b(53) => b(53), 
                           b(52) => b(52), b(51) => b(51), b(50) => b(50), 
                           b(49) => b(49), b(48) => b(48), b(47) => b(47), 
                           b(46) => b(46), b(45) => b(45), b(44) => b(44), 
                           b(43) => b(43), b(42) => b(42), b(41) => b(41), 
                           b(40) => b(40), b(39) => b(39), b(38) => b(38), 
                           b(37) => b(37), b(36) => b(36), b(35) => b(35), 
                           b(34) => b(34), b(33) => b(33), b(32) => b(32), 
                           b(31) => b(31), b(30) => b(30), b(29) => b(29), 
                           b(28) => b(28), b(27) => b(27), b(26) => b(26), 
                           b(25) => b(25), b(24) => b(24), b(23) => b(23), 
                           b(22) => b(22), b(21) => b(21), b(20) => b(20), 
                           b(19) => b(19), b(18) => b(18), b(17) => b(17), 
                           b(16) => b(16), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           cin(15) => carry_15_port, cin(14) => carry_14_port, 
                           cin(13) => carry_13_port, cin(12) => carry_12_port, 
                           cin(11) => carry_11_port, cin(10) => carry_10_port, 
                           cin(9) => carry_9_port, cin(8) => carry_8_port, 
                           cin(7) => carry_7_port, cin(6) => carry_6_port, 
                           cin(5) => carry_5_port, cin(4) => carry_4_port, 
                           cin(3) => carry_3_port, cin(2) => carry_2_port, 
                           cin(1) => carry_1_port, cin(0) => cin, sum(63) => 
                           s(63), sum(62) => s(62), sum(61) => s(61), sum(60) 
                           => s(60), sum(59) => s(59), sum(58) => s(58), 
                           sum(57) => s(57), sum(56) => s(56), sum(55) => s(55)
                           , sum(54) => s(54), sum(53) => s(53), sum(52) => 
                           s(52), sum(51) => s(51), sum(50) => s(50), sum(49) 
                           => s(49), sum(48) => s(48), sum(47) => s(47), 
                           sum(46) => s(46), sum(45) => s(45), sum(44) => s(44)
                           , sum(43) => s(43), sum(42) => s(42), sum(41) => 
                           s(41), sum(40) => s(40), sum(39) => s(39), sum(38) 
                           => s(38), sum(37) => s(37), sum(36) => s(36), 
                           sum(35) => s(35), sum(34) => s(34), sum(33) => s(33)
                           , sum(32) => s(32), sum(31) => s(31), sum(30) => 
                           s(30), sum(29) => s(29), sum(28) => s(28), sum(27) 
                           => s(27), sum(26) => s(26), sum(25) => s(25), 
                           sum(24) => s(24), sum(23) => s(23), sum(22) => s(22)
                           , sum(21) => s(21), sum(20) => s(20), sum(19) => 
                           s(19), sum(18) => s(18), sum(17) => s(17), sum(16) 
                           => s(16), sum(15) => s(15), sum(14) => s(14), 
                           sum(13) => s(13), sum(12) => s(12), sum(11) => s(11)
                           , sum(10) => s(10), sum(9) => s(9), sum(8) => s(8), 
                           sum(7) => s(7), sum(6) => s(6), sum(5) => s(5), 
                           sum(4) => s(4), sum(3) => s(3), sum(2) => s(2), 
                           sum(1) => s(1), sum(0) => s(0));

end SYN_p4_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4Adder_DATA_SIZE16_SPARSITY4 is

   port( cin : in std_logic;  a, b : in std_logic_vector (15 downto 0);  s : 
         out std_logic_vector (15 downto 0);  cout : out std_logic);

end P4Adder_DATA_SIZE16_SPARSITY4;

architecture SYN_p4_adder_arch of P4Adder_DATA_SIZE16_SPARSITY4 is

   component AdderSumGenerator_DATA_SIZE16_SPARSITY4
      port( a, b : in std_logic_vector (15 downto 0);  cin : in 
            std_logic_vector (3 downto 0);  sum : out std_logic_vector (15 
            downto 0));
   end component;
   
   component P4CarryGenerator_DATA_SIZE16_SPARSITY4
      port( a, b : in std_logic_vector (15 downto 0);  cin : in std_logic;  
            cout : out std_logic_vector (3 downto 0));
   end component;
   
   signal carry_3_port, carry_2_port, carry_1_port : std_logic;

begin
   
   CG0 : P4CarryGenerator_DATA_SIZE16_SPARSITY4 port map( a(15) => a(15), a(14)
                           => a(14), a(13) => a(13), a(12) => a(12), a(11) => 
                           a(11), a(10) => a(10), a(9) => a(9), a(8) => a(8), 
                           a(7) => a(7), a(6) => a(6), a(5) => a(5), a(4) => 
                           a(4), a(3) => a(3), a(2) => a(2), a(1) => a(1), a(0)
                           => a(0), b(15) => b(15), b(14) => b(14), b(13) => 
                           b(13), b(12) => b(12), b(11) => b(11), b(10) => 
                           b(10), b(9) => b(9), b(8) => b(8), b(7) => b(7), 
                           b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3) => 
                           b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), cin 
                           => cin, cout(3) => cout, cout(2) => carry_3_port, 
                           cout(1) => carry_2_port, cout(0) => carry_1_port);
   SG0 : AdderSumGenerator_DATA_SIZE16_SPARSITY4 port map( a(15) => a(15), 
                           a(14) => a(14), a(13) => a(13), a(12) => a(12), 
                           a(11) => a(11), a(10) => a(10), a(9) => a(9), a(8) 
                           => a(8), a(7) => a(7), a(6) => a(6), a(5) => a(5), 
                           a(4) => a(4), a(3) => a(3), a(2) => a(2), a(1) => 
                           a(1), a(0) => a(0), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           cin(3) => carry_3_port, cin(2) => carry_2_port, 
                           cin(1) => carry_1_port, cin(0) => cin, sum(15) => 
                           s(15), sum(14) => s(14), sum(13) => s(13), sum(12) 
                           => s(12), sum(11) => s(11), sum(10) => s(10), sum(9)
                           => s(9), sum(8) => s(8), sum(7) => s(7), sum(6) => 
                           s(6), sum(5) => s(5), sum(4) => s(4), sum(3) => s(3)
                           , sum(2) => s(2), sum(1) => s(1), sum(0) => s(0));

end SYN_p4_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderCarrySelect_DATA_SIZE4_0 is

   port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum : 
         out std_logic_vector (3 downto 0));

end AdderCarrySelect_DATA_SIZE4_0;

architecture SYN_adder_carry_select_arch of AdderCarrySelect_DATA_SIZE4_0 is

   component Mux_DATA_SIZE4_0
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (3 downto 0);
            dout : out std_logic_vector (3 downto 0));
   end component;
   
   component Rca_DATA_SIZE4_167
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   component Rca_DATA_SIZE4_0
      port( ci : in std_logic;  a, b : in std_logic_vector (3 downto 0);  s : 
            out std_logic_vector (3 downto 0);  co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sum0_3_port, sum0_2_port, sum0_1_port, 
      sum0_0_port, sum1_3_port, sum1_2_port, sum1_1_port, sum1_0_port, net4592,
      net4593 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA0 : Rca_DATA_SIZE4_0 port map( ci => X_Logic0_port, a(3) => a(3), a(2) =>
                           a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2)
                           => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum0_3_port, s(2) => sum0_2_port, s(1) => 
                           sum0_1_port, s(0) => sum0_0_port, co => net4593);
   RCA1 : Rca_DATA_SIZE4_167 port map( ci => X_Logic1_port, a(3) => a(3), a(2) 
                           => a(2), a(1) => a(1), a(0) => a(0), b(3) => b(3), 
                           b(2) => b(2), b(1) => b(1), b(0) => b(0), s(3) => 
                           sum1_3_port, s(2) => sum1_2_port, s(1) => 
                           sum1_1_port, s(0) => sum1_0_port, co => net4592);
   MUX0 : Mux_DATA_SIZE4_0 port map( sel => sel, din0(3) => sum0_3_port, 
                           din0(2) => sum0_2_port, din0(1) => sum0_1_port, 
                           din0(0) => sum0_0_port, din1(3) => sum1_3_port, 
                           din1(2) => sum1_2_port, din1(1) => sum1_1_port, 
                           din1(0) => sum1_0_port, dout(3) => sum(3), dout(2) 
                           => sum(2), dout(1) => sum(1), dout(0) => sum(0));

end SYN_adder_carry_select_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Adder_DATA_SIZE64 is

   port( cin : in std_logic;  a, b : in std_logic_vector (63 downto 0);  s : 
         out std_logic_vector (63 downto 0);  cout : out std_logic);

end Adder_DATA_SIZE64;

architecture SYN_adder_arch of Adder_DATA_SIZE64 is

   component P4Adder_DATA_SIZE64_SPARSITY4
      port( cin : in std_logic;  a, b : in std_logic_vector (63 downto 0);  s :
            out std_logic_vector (63 downto 0);  cout : out std_logic);
   end component;

begin
   
   ADDER0 : P4Adder_DATA_SIZE64_SPARSITY4 port map( cin => cin, a(63) => a(63),
                           a(62) => a(62), a(61) => a(61), a(60) => a(60), 
                           a(59) => a(59), a(58) => a(58), a(57) => a(57), 
                           a(56) => a(56), a(55) => a(55), a(54) => a(54), 
                           a(53) => a(53), a(52) => a(52), a(51) => a(51), 
                           a(50) => a(50), a(49) => a(49), a(48) => a(48), 
                           a(47) => a(47), a(46) => a(46), a(45) => a(45), 
                           a(44) => a(44), a(43) => a(43), a(42) => a(42), 
                           a(41) => a(41), a(40) => a(40), a(39) => a(39), 
                           a(38) => a(38), a(37) => a(37), a(36) => a(36), 
                           a(35) => a(35), a(34) => a(34), a(33) => a(33), 
                           a(32) => a(32), a(31) => a(31), a(30) => a(30), 
                           a(29) => a(29), a(28) => a(28), a(27) => a(27), 
                           a(26) => a(26), a(25) => a(25), a(24) => a(24), 
                           a(23) => a(23), a(22) => a(22), a(21) => a(21), 
                           a(20) => a(20), a(19) => a(19), a(18) => a(18), 
                           a(17) => a(17), a(16) => a(16), a(15) => a(15), 
                           a(14) => a(14), a(13) => a(13), a(12) => a(12), 
                           a(11) => a(11), a(10) => a(10), a(9) => a(9), a(8) 
                           => a(8), a(7) => a(7), a(6) => a(6), a(5) => a(5), 
                           a(4) => a(4), a(3) => a(3), a(2) => a(2), a(1) => 
                           a(1), a(0) => a(0), b(63) => b(63), b(62) => b(62), 
                           b(61) => b(61), b(60) => b(60), b(59) => b(59), 
                           b(58) => b(58), b(57) => b(57), b(56) => b(56), 
                           b(55) => b(55), b(54) => b(54), b(53) => b(53), 
                           b(52) => b(52), b(51) => b(51), b(50) => b(50), 
                           b(49) => b(49), b(48) => b(48), b(47) => b(47), 
                           b(46) => b(46), b(45) => b(45), b(44) => b(44), 
                           b(43) => b(43), b(42) => b(42), b(41) => b(41), 
                           b(40) => b(40), b(39) => b(39), b(38) => b(38), 
                           b(37) => b(37), b(36) => b(36), b(35) => b(35), 
                           b(34) => b(34), b(33) => b(33), b(32) => b(32), 
                           b(31) => b(31), b(30) => b(30), b(29) => b(29), 
                           b(28) => b(28), b(27) => b(27), b(26) => b(26), 
                           b(25) => b(25), b(24) => b(24), b(23) => b(23), 
                           b(22) => b(22), b(21) => b(21), b(20) => b(20), 
                           b(19) => b(19), b(18) => b(18), b(17) => b(17), 
                           b(16) => b(16), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           s(63) => s(63), s(62) => s(62), s(61) => s(61), 
                           s(60) => s(60), s(59) => s(59), s(58) => s(58), 
                           s(57) => s(57), s(56) => s(56), s(55) => s(55), 
                           s(54) => s(54), s(53) => s(53), s(52) => s(52), 
                           s(51) => s(51), s(50) => s(50), s(49) => s(49), 
                           s(48) => s(48), s(47) => s(47), s(46) => s(46), 
                           s(45) => s(45), s(44) => s(44), s(43) => s(43), 
                           s(42) => s(42), s(41) => s(41), s(40) => s(40), 
                           s(39) => s(39), s(38) => s(38), s(37) => s(37), 
                           s(36) => s(36), s(35) => s(35), s(34) => s(34), 
                           s(33) => s(33), s(32) => s(32), s(31) => s(31), 
                           s(30) => s(30), s(29) => s(29), s(28) => s(28), 
                           s(27) => s(27), s(26) => s(26), s(25) => s(25), 
                           s(24) => s(24), s(23) => s(23), s(22) => s(22), 
                           s(21) => s(21), s(20) => s(20), s(19) => s(19), 
                           s(18) => s(18), s(17) => s(17), s(16) => s(16), 
                           s(15) => s(15), s(14) => s(14), s(13) => s(13), 
                           s(12) => s(12), s(11) => s(11), s(10) => s(10), s(9)
                           => s(9), s(8) => s(8), s(7) => s(7), s(6) => s(6), 
                           s(5) => s(5), s(4) => s(4), s(3) => s(3), s(2) => 
                           s(2), s(1) => s(1), s(0) => s(0), cout => cout);

end SYN_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity BoothEncoder is

   port( din : in std_logic_vector (2 downto 0);  sel : out std_logic_vector (2
         downto 0));

end BoothEncoder;

architecture SYN_booth_encoder_arch of BoothEncoder is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n8, n2, n3, n4, n5, n6, n7 : std_logic;

begin
   
   U3 : OAI21_X1 port map( B1 => din(1), B2 => n5, A => n3, ZN => n8);
   U4 : MUX2_X2 port map( A => n6, B => n7, S => din(1), Z => sel(0));
   U5 : CLKBUF_X2 port map( A => n8, Z => sel(1));
   U6 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => sel(2));
   U7 : MUX2_X1 port map( A => n4, B => din(2), S => din(1), Z => n2);
   U8 : INV_X1 port map( A => din(2), ZN => n5);
   U9 : NOR2_X1 port map( A1 => din(2), A2 => n4, ZN => n7);
   U10 : INV_X1 port map( A => n3, ZN => n6);
   U11 : NAND2_X1 port map( A1 => din(2), A2 => n4, ZN => n3);
   U12 : INV_X1 port map( A => din(0), ZN => n4);

end SYN_booth_encoder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Adder_DATA_SIZE16 is

   port( cin : in std_logic;  a, b : in std_logic_vector (15 downto 0);  s : 
         out std_logic_vector (15 downto 0);  cout : out std_logic);

end Adder_DATA_SIZE16;

architecture SYN_adder_arch of Adder_DATA_SIZE16 is

   component P4Adder_DATA_SIZE16_SPARSITY4
      port( cin : in std_logic;  a, b : in std_logic_vector (15 downto 0);  s :
            out std_logic_vector (15 downto 0);  cout : out std_logic);
   end component;

begin
   
   ADDER0 : P4Adder_DATA_SIZE16_SPARSITY4 port map( cin => cin, a(15) => a(15),
                           a(14) => a(14), a(13) => a(13), a(12) => a(12), 
                           a(11) => a(11), a(10) => a(10), a(9) => a(9), a(8) 
                           => a(8), a(7) => a(7), a(6) => a(6), a(5) => a(5), 
                           a(4) => a(4), a(3) => a(3), a(2) => a(2), a(1) => 
                           a(1), a(0) => a(0), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           s(15) => s(15), s(14) => s(14), s(13) => s(13), 
                           s(12) => s(12), s(11) => s(11), s(10) => s(10), s(9)
                           => s(9), s(8) => s(8), s(7) => s(7), s(6) => s(6), 
                           s(5) => s(5), s(4) => s(4), s(3) => s(3), s(2) => 
                           s(2), s(1) => s(1), s(0) => s(0), cout => cout);

end SYN_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AdderSumGenerator_DATA_SIZE32_SPARSITY4_0 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic_vector 
         (7 downto 0);  sum : out std_logic_vector (31 downto 0));

end AdderSumGenerator_DATA_SIZE32_SPARSITY4_0;

architecture SYN_adder_sum_generator_arch of 
   AdderSumGenerator_DATA_SIZE32_SPARSITY4_0 is

   component AdderCarrySelect_DATA_SIZE4_77
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_78
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_79
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_80
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_81
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_82
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_83
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;
   
   component AdderCarrySelect_DATA_SIZE4_0
      port( a, b : in std_logic_vector (3 downto 0);  sel : in std_logic;  sum 
            : out std_logic_vector (3 downto 0));
   end component;

begin
   
   ACSi_0 : AdderCarrySelect_DATA_SIZE4_0 port map( a(3) => a(3), a(2) => a(2),
                           a(1) => a(1), a(0) => a(0), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), sel => cin(0), 
                           sum(3) => sum(3), sum(2) => sum(2), sum(1) => sum(1)
                           , sum(0) => sum(0));
   ACSi_1 : AdderCarrySelect_DATA_SIZE4_83 port map( a(3) => a(7), a(2) => a(6)
                           , a(1) => a(5), a(0) => a(4), b(3) => b(7), b(2) => 
                           b(6), b(1) => b(5), b(0) => b(4), sel => cin(1), 
                           sum(3) => sum(7), sum(2) => sum(6), sum(1) => sum(5)
                           , sum(0) => sum(4));
   ACSi_2 : AdderCarrySelect_DATA_SIZE4_82 port map( a(3) => a(11), a(2) => 
                           a(10), a(1) => a(9), a(0) => a(8), b(3) => b(11), 
                           b(2) => b(10), b(1) => b(9), b(0) => b(8), sel => 
                           cin(2), sum(3) => sum(11), sum(2) => sum(10), sum(1)
                           => sum(9), sum(0) => sum(8));
   ACSi_3 : AdderCarrySelect_DATA_SIZE4_81 port map( a(3) => a(15), a(2) => 
                           a(14), a(1) => a(13), a(0) => a(12), b(3) => b(15), 
                           b(2) => b(14), b(1) => b(13), b(0) => b(12), sel => 
                           cin(3), sum(3) => sum(15), sum(2) => sum(14), sum(1)
                           => sum(13), sum(0) => sum(12));
   ACSi_4 : AdderCarrySelect_DATA_SIZE4_80 port map( a(3) => a(19), a(2) => 
                           a(18), a(1) => a(17), a(0) => a(16), b(3) => b(19), 
                           b(2) => b(18), b(1) => b(17), b(0) => b(16), sel => 
                           cin(4), sum(3) => sum(19), sum(2) => sum(18), sum(1)
                           => sum(17), sum(0) => sum(16));
   ACSi_5 : AdderCarrySelect_DATA_SIZE4_79 port map( a(3) => a(23), a(2) => 
                           a(22), a(1) => a(21), a(0) => a(20), b(3) => b(23), 
                           b(2) => b(22), b(1) => b(21), b(0) => b(20), sel => 
                           cin(5), sum(3) => sum(23), sum(2) => sum(22), sum(1)
                           => sum(21), sum(0) => sum(20));
   ACSi_6 : AdderCarrySelect_DATA_SIZE4_78 port map( a(3) => a(27), a(2) => 
                           a(26), a(1) => a(25), a(0) => a(24), b(3) => b(27), 
                           b(2) => b(26), b(1) => b(25), b(0) => b(24), sel => 
                           cin(6), sum(3) => sum(27), sum(2) => sum(26), sum(1)
                           => sum(25), sum(0) => sum(24));
   ACSi_7 : AdderCarrySelect_DATA_SIZE4_77 port map( a(3) => a(31), a(2) => 
                           a(30), a(1) => a(29), a(0) => a(28), b(3) => b(31), 
                           b(2) => b(30), b(1) => b(29), b(0) => b(28), sel => 
                           cin(7), sum(3) => sum(31), sum(2) => sum(30), sum(1)
                           => sum(29), sum(0) => sum(28));

end SYN_adder_sum_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4CarryGenerator_DATA_SIZE32_SPARSITY4_0 is

   port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  cout :
         out std_logic_vector (7 downto 0));

end P4CarryGenerator_DATA_SIZE32_SPARSITY4_0;

architecture SYN_p4_carry_generator_arch of 
   P4CarryGenerator_DATA_SIZE32_SPARSITY4_0 is

   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal cout_7_port, cout_6_port, cout_5_port, cout_4_port, cout_3_port, 
      cout_2_port, cout_1_port, cout_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9
      , n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, 
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, 
      n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96
      , n97, n98, n99, n100, n101 : std_logic;

begin
   cout <= ( cout_7_port, cout_6_port, cout_5_port, cout_4_port, cout_3_port, 
      cout_2_port, cout_1_port, cout_0_port );
   
   U1 : OAI22_X1 port map( A1 => n1, A2 => n2, B1 => n3, B2 => n4, ZN => 
                           cout_7_port);
   U2 : AOI22_X1 port map( A1 => b(30), A2 => n5, B1 => a(30), B2 => n6, ZN => 
                           n4);
   U3 : OR2_X1 port map( A1 => n6, A2 => a(30), ZN => n5);
   U4 : OAI21_X1 port map( B1 => n7, B2 => n8, A => n9, ZN => n6);
   U5 : OAI21_X1 port map( B1 => b(29), B2 => a(29), A => n10, ZN => n9);
   U6 : INV_X1 port map( A => n11, ZN => n10);
   U7 : AOI21_X1 port map( B1 => cout_6_port, B2 => a(28), A => n12, ZN => n11)
                           ;
   U8 : INV_X1 port map( A => n13, ZN => n12);
   U9 : OAI21_X1 port map( B1 => a(28), B2 => cout_6_port, A => b(28), ZN => 
                           n13);
   U10 : INV_X1 port map( A => b(29), ZN => n8);
   U11 : INV_X1 port map( A => a(29), ZN => n7);
   U12 : NOR2_X1 port map( A1 => b(31), A2 => a(31), ZN => n3);
   U13 : INV_X1 port map( A => b(31), ZN => n2);
   U14 : INV_X1 port map( A => a(31), ZN => n1);
   U15 : OAI21_X1 port map( B1 => n14, B2 => n15, A => n16, ZN => cout_6_port);
   U16 : OAI21_X1 port map( B1 => a(27), B2 => n17, A => b(27), ZN => n16);
   U17 : INV_X1 port map( A => n14, ZN => n17);
   U18 : INV_X1 port map( A => a(27), ZN => n15);
   U19 : AOI21_X1 port map( B1 => a(26), B2 => b(26), A => n18, ZN => n14);
   U20 : INV_X1 port map( A => n19, ZN => n18);
   U21 : OAI22_X1 port map( A1 => n20, A2 => n21, B1 => a(26), B2 => b(26), ZN 
                           => n19);
   U22 : NOR2_X1 port map( A1 => n22, A2 => n23, ZN => n21);
   U23 : AOI22_X1 port map( A1 => n22, A2 => n23, B1 => n24, B2 => n25, ZN => 
                           n20);
   U24 : OAI21_X1 port map( B1 => a(24), B2 => cout_5_port, A => b(24), ZN => 
                           n25);
   U25 : NAND2_X1 port map( A1 => a(24), A2 => cout_5_port, ZN => n24);
   U26 : INV_X1 port map( A => b(25), ZN => n23);
   U27 : INV_X1 port map( A => a(25), ZN => n22);
   U28 : OAI22_X1 port map( A1 => n26, A2 => n27, B1 => n28, B2 => n29, ZN => 
                           cout_5_port);
   U29 : AOI22_X1 port map( A1 => b(22), A2 => n30, B1 => a(22), B2 => n31, ZN 
                           => n29);
   U30 : OR2_X1 port map( A1 => n31, A2 => a(22), ZN => n30);
   U31 : OAI21_X1 port map( B1 => n32, B2 => n33, A => n34, ZN => n31);
   U32 : OAI21_X1 port map( B1 => b(21), B2 => a(21), A => n35, ZN => n34);
   U33 : OAI21_X1 port map( B1 => n36, B2 => n37, A => n38, ZN => n35);
   U34 : OAI21_X1 port map( B1 => a(20), B2 => cout_4_port, A => b(20), ZN => 
                           n38);
   U35 : INV_X1 port map( A => a(20), ZN => n37);
   U36 : INV_X1 port map( A => cout_4_port, ZN => n36);
   U37 : INV_X1 port map( A => b(21), ZN => n33);
   U38 : INV_X1 port map( A => a(21), ZN => n32);
   U39 : NOR2_X1 port map( A1 => b(23), A2 => a(23), ZN => n28);
   U40 : INV_X1 port map( A => b(23), ZN => n27);
   U41 : INV_X1 port map( A => a(23), ZN => n26);
   U42 : OAI211_X1 port map( C1 => n39, C2 => n40, A => n41, B => n42, ZN => 
                           cout_4_port);
   U43 : OAI211_X1 port map( C1 => b(19), C2 => a(19), A => cout_3_port, B => 
                           n43, ZN => n42);
   U44 : AOI221_X1 port map( B1 => n44, B2 => n45, C1 => n46, C2 => n47, A => 
                           n48, ZN => n43);
   U45 : OAI21_X1 port map( B1 => n49, B2 => a(19), A => b(19), ZN => n41);
   U46 : INV_X1 port map( A => a(19), ZN => n40);
   U47 : INV_X1 port map( A => n49, ZN => n39);
   U48 : AOI21_X1 port map( B1 => n44, B2 => n50, A => n51, ZN => n49);
   U49 : INV_X1 port map( A => n52, ZN => n51);
   U50 : OAI21_X1 port map( B1 => n50, B2 => n44, A => n45, ZN => n52);
   U51 : INV_X1 port map( A => b(18), ZN => n45);
   U52 : AOI21_X1 port map( B1 => a(17), B2 => b(17), A => n53, ZN => n50);
   U53 : NOR3_X1 port map( A1 => n46, A2 => n48, A3 => n47, ZN => n53);
   U54 : INV_X1 port map( A => b(16), ZN => n47);
   U55 : NOR2_X1 port map( A1 => b(17), A2 => a(17), ZN => n48);
   U56 : INV_X1 port map( A => a(16), ZN => n46);
   U57 : INV_X1 port map( A => a(18), ZN => n44);
   U58 : INV_X1 port map( A => n54, ZN => cout_3_port);
   U59 : OAI22_X1 port map( A1 => a(15), A2 => n55, B1 => b(15), B2 => n56, ZN 
                           => n54);
   U60 : AND2_X1 port map( A1 => n55, A2 => a(15), ZN => n56);
   U61 : INV_X1 port map( A => n57, ZN => n55);
   U62 : OAI22_X1 port map( A1 => a(14), A2 => n58, B1 => b(14), B2 => n59, ZN 
                           => n57);
   U63 : AND2_X1 port map( A1 => n58, A2 => a(14), ZN => n59);
   U64 : OAI21_X1 port map( B1 => n60, B2 => n61, A => n62, ZN => n58);
   U65 : OAI21_X1 port map( B1 => b(13), B2 => a(13), A => n63, ZN => n62);
   U66 : INV_X1 port map( A => n64, ZN => n63);
   U67 : AOI21_X1 port map( B1 => cout_2_port, B2 => a(12), A => n65, ZN => n64
                           );
   U68 : INV_X1 port map( A => n66, ZN => n65);
   U69 : OAI21_X1 port map( B1 => a(12), B2 => cout_2_port, A => b(12), ZN => 
                           n66);
   U70 : INV_X1 port map( A => b(13), ZN => n61);
   U71 : INV_X1 port map( A => a(13), ZN => n60);
   U72 : OAI21_X1 port map( B1 => n67, B2 => n68, A => n69, ZN => cout_2_port);
   U73 : OAI21_X1 port map( B1 => a(11), B2 => n70, A => b(11), ZN => n69);
   U74 : INV_X1 port map( A => n67, ZN => n70);
   U75 : INV_X1 port map( A => a(11), ZN => n68);
   U76 : AOI21_X1 port map( B1 => a(10), B2 => b(10), A => n71, ZN => n67);
   U77 : INV_X1 port map( A => n72, ZN => n71);
   U78 : OAI22_X1 port map( A1 => n73, A2 => n74, B1 => a(10), B2 => b(10), ZN 
                           => n72);
   U79 : NOR2_X1 port map( A1 => n75, A2 => n76, ZN => n74);
   U80 : AOI22_X1 port map( A1 => n75, A2 => n76, B1 => n77, B2 => n78, ZN => 
                           n73);
   U81 : OAI21_X1 port map( B1 => a(8), B2 => cout_1_port, A => b(8), ZN => n78
                           );
   U82 : NAND2_X1 port map( A1 => a(8), A2 => cout_1_port, ZN => n77);
   U83 : INV_X1 port map( A => b(9), ZN => n76);
   U84 : INV_X1 port map( A => a(9), ZN => n75);
   U85 : OAI21_X1 port map( B1 => n79, B2 => n80, A => n81, ZN => cout_1_port);
   U86 : OAI21_X1 port map( B1 => b(7), B2 => a(7), A => n82, ZN => n81);
   U87 : OAI21_X1 port map( B1 => n83, B2 => n84, A => n85, ZN => n82);
   U88 : OAI21_X1 port map( B1 => a(6), B2 => n86, A => b(6), ZN => n85);
   U89 : INV_X1 port map( A => n83, ZN => n86);
   U90 : INV_X1 port map( A => a(6), ZN => n84);
   U91 : AOI22_X1 port map( A1 => a(5), A2 => b(5), B1 => n87, B2 => n88, ZN =>
                           n83);
   U92 : INV_X1 port map( A => n89, ZN => n88);
   U93 : AOI22_X1 port map( A1 => b(4), A2 => n90, B1 => a(4), B2 => 
                           cout_0_port, ZN => n89);
   U94 : OR2_X1 port map( A1 => a(4), A2 => cout_0_port, ZN => n90);
   U95 : OR2_X1 port map( A1 => b(5), A2 => a(5), ZN => n87);
   U96 : INV_X1 port map( A => b(7), ZN => n80);
   U97 : INV_X1 port map( A => a(7), ZN => n79);
   U98 : INV_X1 port map( A => n91, ZN => cout_0_port);
   U99 : OAI22_X1 port map( A1 => a(3), A2 => n92, B1 => b(3), B2 => n93, ZN =>
                           n91);
   U100 : AND2_X1 port map( A1 => n92, A2 => a(3), ZN => n93);
   U101 : INV_X1 port map( A => n94, ZN => n92);
   U102 : OAI22_X1 port map( A1 => a(2), A2 => n95, B1 => b(2), B2 => n96, ZN 
                           => n94);
   U103 : AND2_X1 port map( A1 => n95, A2 => a(2), ZN => n96);
   U104 : INV_X1 port map( A => n97, ZN => n95);
   U105 : AOI22_X1 port map( A1 => a(1), A2 => b(1), B1 => n98, B2 => n99, ZN 
                           => n97);
   U106 : INV_X1 port map( A => n100, ZN => n99);
   U107 : AOI22_X1 port map( A1 => cin, A2 => n101, B1 => b(0), B2 => a(0), ZN 
                           => n100);
   U108 : OR2_X1 port map( A1 => b(0), A2 => a(0), ZN => n101);
   U109 : OR2_X1 port map( A1 => b(1), A2 => a(1), ZN => n98);

end SYN_p4_carry_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Sipo_DATA_SIZE32 is

   port( rst, en, clk, din : in std_logic;  dout : out std_logic_vector (31 
         downto 0));

end Sipo_DATA_SIZE32;

architecture SYN_sipo_arch of Sipo_DATA_SIZE32 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal dout_31_port, dout_30_port, dout_29_port, dout_28_port, dout_27_port,
      dout_26_port, dout_25_port, dout_24_port, dout_23_port, dout_22_port, 
      dout_21_port, dout_20_port, dout_19_port, dout_18_port, dout_17_port, 
      dout_16_port, dout_15_port, dout_14_port, dout_13_port, dout_12_port, 
      dout_11_port, dout_10_port, dout_9_port, dout_8_port, dout_7_port, 
      dout_6_port, dout_5_port, dout_4_port, dout_3_port, dout_2_port, 
      dout_1_port, dout_0_port, n101, n102, n103, n104, n105, n106, n107, n108,
      n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, 
      n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, 
      n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, 
      n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, 
      n157, n158, n159, n160, n161, n162, n163, n1, n2, n3, n4, n5, n6, n7, n8,
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67
      , n68, n69, n70, net108809, net108810, net108811, net108812, net108813, 
      net108814, net108815, net108816, net108817, net108818, net108819, 
      net108820, net108821, net108822, net108823, net108824, net108825, 
      net108826, net108827, net108828, net108829, net108830, net108831, 
      net108832, net108833, net108834, net108835, net108836, net108837, 
      net108838, net108839, net108840 : std_logic;

begin
   dout <= ( dout_31_port, dout_30_port, dout_29_port, dout_28_port, 
      dout_27_port, dout_26_port, dout_25_port, dout_24_port, dout_23_port, 
      dout_22_port, dout_21_port, dout_20_port, dout_19_port, dout_18_port, 
      dout_17_port, dout_16_port, dout_15_port, dout_14_port, dout_13_port, 
      dout_12_port, dout_11_port, dout_10_port, dout_9_port, dout_8_port, 
      dout_7_port, dout_6_port, dout_5_port, dout_4_port, dout_3_port, 
      dout_2_port, dout_1_port, dout_0_port );
   
   dout_reg_0_inst : DFFR_X1 port map( D => n163, CK => clk, RN => rst, Q => 
                           dout_0_port, QN => net108840);
   data_reg_1_inst : DFF_X1 port map( D => n162, CK => clk, Q => n1, QN => n70)
                           ;
   dout_reg_1_inst : DFFR_X1 port map( D => n161, CK => clk, RN => rst, Q => 
                           dout_1_port, QN => net108839);
   data_reg_2_inst : DFF_X1 port map( D => n160, CK => clk, Q => n2, QN => n69)
                           ;
   dout_reg_2_inst : DFFR_X1 port map( D => n159, CK => clk, RN => rst, Q => 
                           dout_2_port, QN => net108838);
   data_reg_3_inst : DFF_X1 port map( D => n158, CK => clk, Q => n3, QN => n68)
                           ;
   dout_reg_3_inst : DFFR_X1 port map( D => n157, CK => clk, RN => rst, Q => 
                           dout_3_port, QN => net108837);
   data_reg_4_inst : DFF_X1 port map( D => n156, CK => clk, Q => n4, QN => n67)
                           ;
   dout_reg_4_inst : DFFR_X1 port map( D => n155, CK => clk, RN => rst, Q => 
                           dout_4_port, QN => net108836);
   data_reg_5_inst : DFF_X1 port map( D => n154, CK => clk, Q => n5, QN => n66)
                           ;
   dout_reg_5_inst : DFFR_X1 port map( D => n153, CK => clk, RN => rst, Q => 
                           dout_5_port, QN => net108835);
   data_reg_6_inst : DFF_X1 port map( D => n152, CK => clk, Q => n6, QN => n65)
                           ;
   dout_reg_6_inst : DFFR_X1 port map( D => n151, CK => clk, RN => rst, Q => 
                           dout_6_port, QN => net108834);
   data_reg_7_inst : DFF_X1 port map( D => n150, CK => clk, Q => n7, QN => n64)
                           ;
   dout_reg_7_inst : DFFR_X1 port map( D => n149, CK => clk, RN => rst, Q => 
                           dout_7_port, QN => net108833);
   data_reg_8_inst : DFF_X1 port map( D => n148, CK => clk, Q => n8, QN => n63)
                           ;
   dout_reg_8_inst : DFFR_X1 port map( D => n147, CK => clk, RN => rst, Q => 
                           dout_8_port, QN => net108832);
   data_reg_9_inst : DFF_X1 port map( D => n146, CK => clk, Q => n9, QN => n62)
                           ;
   dout_reg_9_inst : DFFR_X1 port map( D => n145, CK => clk, RN => rst, Q => 
                           dout_9_port, QN => net108831);
   data_reg_10_inst : DFF_X1 port map( D => n144, CK => clk, Q => n10, QN => 
                           n61);
   dout_reg_10_inst : DFFR_X1 port map( D => n143, CK => clk, RN => rst, Q => 
                           dout_10_port, QN => net108830);
   data_reg_11_inst : DFF_X1 port map( D => n142, CK => clk, Q => n11, QN => 
                           n60);
   dout_reg_11_inst : DFFR_X1 port map( D => n141, CK => clk, RN => rst, Q => 
                           dout_11_port, QN => net108829);
   data_reg_12_inst : DFF_X1 port map( D => n140, CK => clk, Q => n12, QN => 
                           n59);
   dout_reg_12_inst : DFFR_X1 port map( D => n139, CK => clk, RN => rst, Q => 
                           dout_12_port, QN => net108828);
   data_reg_13_inst : DFF_X1 port map( D => n138, CK => clk, Q => n13, QN => 
                           n58);
   dout_reg_13_inst : DFFR_X1 port map( D => n137, CK => clk, RN => rst, Q => 
                           dout_13_port, QN => net108827);
   data_reg_14_inst : DFF_X1 port map( D => n136, CK => clk, Q => n14, QN => 
                           n57);
   dout_reg_14_inst : DFFR_X1 port map( D => n135, CK => clk, RN => rst, Q => 
                           dout_14_port, QN => net108826);
   data_reg_15_inst : DFF_X1 port map( D => n134, CK => clk, Q => n15, QN => 
                           n56);
   dout_reg_15_inst : DFFR_X1 port map( D => n133, CK => clk, RN => rst, Q => 
                           dout_15_port, QN => net108825);
   data_reg_16_inst : DFF_X1 port map( D => n132, CK => clk, Q => n16, QN => 
                           n55);
   dout_reg_16_inst : DFFR_X1 port map( D => n131, CK => clk, RN => rst, Q => 
                           dout_16_port, QN => net108824);
   data_reg_17_inst : DFF_X1 port map( D => n130, CK => clk, Q => n17, QN => 
                           n54);
   dout_reg_17_inst : DFFR_X1 port map( D => n129, CK => clk, RN => rst, Q => 
                           dout_17_port, QN => net108823);
   data_reg_18_inst : DFF_X1 port map( D => n128, CK => clk, Q => n18, QN => 
                           n53);
   dout_reg_18_inst : DFFR_X1 port map( D => n127, CK => clk, RN => rst, Q => 
                           dout_18_port, QN => net108822);
   data_reg_19_inst : DFF_X1 port map( D => n126, CK => clk, Q => n19, QN => 
                           n52);
   dout_reg_19_inst : DFFR_X1 port map( D => n125, CK => clk, RN => rst, Q => 
                           dout_19_port, QN => net108821);
   data_reg_20_inst : DFF_X1 port map( D => n124, CK => clk, Q => n20, QN => 
                           n51);
   dout_reg_20_inst : DFFR_X1 port map( D => n123, CK => clk, RN => rst, Q => 
                           dout_20_port, QN => net108820);
   data_reg_21_inst : DFF_X1 port map( D => n122, CK => clk, Q => n21, QN => 
                           n50);
   dout_reg_21_inst : DFFR_X1 port map( D => n121, CK => clk, RN => rst, Q => 
                           dout_21_port, QN => net108819);
   data_reg_22_inst : DFF_X1 port map( D => n120, CK => clk, Q => n22, QN => 
                           n49);
   dout_reg_22_inst : DFFR_X1 port map( D => n119, CK => clk, RN => rst, Q => 
                           dout_22_port, QN => net108818);
   data_reg_23_inst : DFF_X1 port map( D => n118, CK => clk, Q => n23, QN => 
                           n48);
   dout_reg_23_inst : DFFR_X1 port map( D => n117, CK => clk, RN => rst, Q => 
                           dout_23_port, QN => net108817);
   data_reg_24_inst : DFF_X1 port map( D => n116, CK => clk, Q => n24, QN => 
                           n47);
   dout_reg_24_inst : DFFR_X1 port map( D => n115, CK => clk, RN => rst, Q => 
                           dout_24_port, QN => net108816);
   data_reg_25_inst : DFF_X1 port map( D => n114, CK => clk, Q => n25, QN => 
                           n46);
   dout_reg_25_inst : DFFR_X1 port map( D => n113, CK => clk, RN => rst, Q => 
                           dout_25_port, QN => net108815);
   data_reg_26_inst : DFF_X1 port map( D => n112, CK => clk, Q => n26, QN => 
                           n45);
   dout_reg_26_inst : DFFR_X1 port map( D => n111, CK => clk, RN => rst, Q => 
                           dout_26_port, QN => net108814);
   data_reg_27_inst : DFF_X1 port map( D => n110, CK => clk, Q => n27, QN => 
                           n44);
   dout_reg_27_inst : DFFR_X1 port map( D => n109, CK => clk, RN => rst, Q => 
                           dout_27_port, QN => net108813);
   data_reg_28_inst : DFF_X1 port map( D => n108, CK => clk, Q => n28, QN => 
                           n43);
   dout_reg_28_inst : DFFR_X1 port map( D => n107, CK => clk, RN => rst, Q => 
                           dout_28_port, QN => net108812);
   data_reg_29_inst : DFF_X1 port map( D => n106, CK => clk, Q => n29, QN => 
                           n42);
   dout_reg_29_inst : DFFR_X1 port map( D => n105, CK => clk, RN => rst, Q => 
                           dout_29_port, QN => net108811);
   data_reg_30_inst : DFF_X1 port map( D => n104, CK => clk, Q => n30, QN => 
                           n41);
   dout_reg_30_inst : DFFR_X1 port map( D => n103, CK => clk, RN => rst, Q => 
                           dout_30_port, QN => net108810);
   data_reg_31_inst : DFF_X1 port map( D => n102, CK => clk, Q => n31, QN => 
                           n40);
   dout_reg_31_inst : DFFR_X1 port map( D => n101, CK => clk, RN => rst, Q => 
                           dout_31_port, QN => net108809);
   U3 : NAND2_X2 port map( A1 => rst, A2 => n37, ZN => n39);
   U4 : NAND2_X2 port map( A1 => rst, A2 => n34, ZN => n37);
   U5 : BUF_X1 port map( A => n35, Z => n32);
   U6 : BUF_X1 port map( A => n35, Z => n33);
   U7 : BUF_X1 port map( A => n35, Z => n34);
   U8 : INV_X1 port map( A => en, ZN => n35);
   U9 : MUX2_X1 port map( A => n36, B => dout_0_port, S => n33, Z => n163);
   U10 : AND2_X1 port map( A1 => din, A2 => rst, ZN => n36);
   U11 : OAI22_X1 port map( A1 => n70, A2 => n37, B1 => n38, B2 => n39, ZN => 
                           n162);
   U12 : INV_X1 port map( A => din, ZN => n38);
   U13 : MUX2_X1 port map( A => n1, B => dout_1_port, S => n32, Z => n161);
   U14 : OAI22_X1 port map( A1 => n69, A2 => n37, B1 => n70, B2 => n39, ZN => 
                           n160);
   U15 : MUX2_X1 port map( A => n2, B => dout_2_port, S => n32, Z => n159);
   U16 : OAI22_X1 port map( A1 => n68, A2 => n37, B1 => n69, B2 => n39, ZN => 
                           n158);
   U17 : MUX2_X1 port map( A => n3, B => dout_3_port, S => n32, Z => n157);
   U18 : OAI22_X1 port map( A1 => n67, A2 => n37, B1 => n68, B2 => n39, ZN => 
                           n156);
   U19 : MUX2_X1 port map( A => n4, B => dout_4_port, S => n32, Z => n155);
   U20 : OAI22_X1 port map( A1 => n66, A2 => n37, B1 => n67, B2 => n39, ZN => 
                           n154);
   U21 : MUX2_X1 port map( A => n5, B => dout_5_port, S => n32, Z => n153);
   U22 : OAI22_X1 port map( A1 => n65, A2 => n37, B1 => n66, B2 => n39, ZN => 
                           n152);
   U23 : MUX2_X1 port map( A => n6, B => dout_6_port, S => n32, Z => n151);
   U24 : OAI22_X1 port map( A1 => n64, A2 => n37, B1 => n65, B2 => n39, ZN => 
                           n150);
   U25 : MUX2_X1 port map( A => n7, B => dout_7_port, S => n32, Z => n149);
   U26 : OAI22_X1 port map( A1 => n63, A2 => n37, B1 => n64, B2 => n39, ZN => 
                           n148);
   U27 : MUX2_X1 port map( A => n8, B => dout_8_port, S => n32, Z => n147);
   U28 : OAI22_X1 port map( A1 => n62, A2 => n37, B1 => n63, B2 => n39, ZN => 
                           n146);
   U29 : MUX2_X1 port map( A => n9, B => dout_9_port, S => n32, Z => n145);
   U30 : OAI22_X1 port map( A1 => n61, A2 => n37, B1 => n62, B2 => n39, ZN => 
                           n144);
   U31 : MUX2_X1 port map( A => n10, B => dout_10_port, S => n32, Z => n143);
   U32 : OAI22_X1 port map( A1 => n60, A2 => n37, B1 => n61, B2 => n39, ZN => 
                           n142);
   U33 : MUX2_X1 port map( A => n11, B => dout_11_port, S => n32, Z => n141);
   U34 : OAI22_X1 port map( A1 => n59, A2 => n37, B1 => n60, B2 => n39, ZN => 
                           n140);
   U35 : MUX2_X1 port map( A => n12, B => dout_12_port, S => n33, Z => n139);
   U36 : OAI22_X1 port map( A1 => n58, A2 => n37, B1 => n59, B2 => n39, ZN => 
                           n138);
   U37 : MUX2_X1 port map( A => n13, B => dout_13_port, S => n33, Z => n137);
   U38 : OAI22_X1 port map( A1 => n57, A2 => n37, B1 => n58, B2 => n39, ZN => 
                           n136);
   U39 : MUX2_X1 port map( A => n14, B => dout_14_port, S => n33, Z => n135);
   U40 : OAI22_X1 port map( A1 => n56, A2 => n37, B1 => n57, B2 => n39, ZN => 
                           n134);
   U41 : MUX2_X1 port map( A => n15, B => dout_15_port, S => n33, Z => n133);
   U42 : OAI22_X1 port map( A1 => n55, A2 => n37, B1 => n56, B2 => n39, ZN => 
                           n132);
   U43 : MUX2_X1 port map( A => n16, B => dout_16_port, S => n33, Z => n131);
   U44 : OAI22_X1 port map( A1 => n54, A2 => n37, B1 => n55, B2 => n39, ZN => 
                           n130);
   U45 : MUX2_X1 port map( A => n17, B => dout_17_port, S => n33, Z => n129);
   U46 : OAI22_X1 port map( A1 => n53, A2 => n37, B1 => n54, B2 => n39, ZN => 
                           n128);
   U47 : MUX2_X1 port map( A => n18, B => dout_18_port, S => n33, Z => n127);
   U48 : OAI22_X1 port map( A1 => n52, A2 => n37, B1 => n53, B2 => n39, ZN => 
                           n126);
   U49 : MUX2_X1 port map( A => n19, B => dout_19_port, S => n33, Z => n125);
   U50 : OAI22_X1 port map( A1 => n51, A2 => n37, B1 => n52, B2 => n39, ZN => 
                           n124);
   U51 : MUX2_X1 port map( A => n20, B => dout_20_port, S => n33, Z => n123);
   U52 : OAI22_X1 port map( A1 => n50, A2 => n37, B1 => n51, B2 => n39, ZN => 
                           n122);
   U53 : MUX2_X1 port map( A => n21, B => dout_21_port, S => n33, Z => n121);
   U54 : OAI22_X1 port map( A1 => n49, A2 => n37, B1 => n50, B2 => n39, ZN => 
                           n120);
   U55 : MUX2_X1 port map( A => n22, B => dout_22_port, S => n33, Z => n119);
   U56 : OAI22_X1 port map( A1 => n48, A2 => n37, B1 => n49, B2 => n39, ZN => 
                           n118);
   U57 : MUX2_X1 port map( A => n23, B => dout_23_port, S => n34, Z => n117);
   U58 : OAI22_X1 port map( A1 => n47, A2 => n37, B1 => n48, B2 => n39, ZN => 
                           n116);
   U59 : MUX2_X1 port map( A => n24, B => dout_24_port, S => n34, Z => n115);
   U60 : OAI22_X1 port map( A1 => n46, A2 => n37, B1 => n47, B2 => n39, ZN => 
                           n114);
   U61 : MUX2_X1 port map( A => n25, B => dout_25_port, S => n34, Z => n113);
   U62 : OAI22_X1 port map( A1 => n45, A2 => n37, B1 => n46, B2 => n39, ZN => 
                           n112);
   U63 : MUX2_X1 port map( A => n26, B => dout_26_port, S => n34, Z => n111);
   U64 : OAI22_X1 port map( A1 => n44, A2 => n37, B1 => n45, B2 => n39, ZN => 
                           n110);
   U65 : MUX2_X1 port map( A => n27, B => dout_27_port, S => n34, Z => n109);
   U66 : OAI22_X1 port map( A1 => n43, A2 => n37, B1 => n44, B2 => n39, ZN => 
                           n108);
   U67 : MUX2_X1 port map( A => n28, B => dout_28_port, S => n34, Z => n107);
   U68 : OAI22_X1 port map( A1 => n42, A2 => n37, B1 => n43, B2 => n39, ZN => 
                           n106);
   U69 : MUX2_X1 port map( A => n29, B => dout_29_port, S => n34, Z => n105);
   U70 : OAI22_X1 port map( A1 => n41, A2 => n37, B1 => n42, B2 => n39, ZN => 
                           n104);
   U71 : MUX2_X1 port map( A => n30, B => dout_30_port, S => n34, Z => n103);
   U72 : OAI22_X1 port map( A1 => n40, A2 => n37, B1 => n41, B2 => n39, ZN => 
                           n102);
   U73 : MUX2_X1 port map( A => n31, B => dout_31_port, S => n32, Z => n101);

end SYN_sipo_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE64 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (63 downto 0);
         dout : out std_logic_vector (63 downto 0));

end Reg_DATA_SIZE64;

architecture SYN_reg_arch of Reg_DATA_SIZE64 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal dout_63_port, dout_62_port, dout_61_port, dout_60_port, dout_59_port,
      dout_58_port, dout_57_port, dout_56_port, dout_55_port, dout_54_port, 
      dout_53_port, dout_52_port, dout_51_port, dout_50_port, dout_49_port, 
      dout_48_port, dout_47_port, dout_46_port, dout_45_port, dout_44_port, 
      dout_43_port, dout_42_port, dout_41_port, dout_40_port, dout_39_port, 
      dout_38_port, dout_37_port, dout_36_port, dout_35_port, dout_34_port, 
      dout_33_port, dout_32_port, dout_31_port, dout_30_port, dout_29_port, 
      dout_28_port, dout_27_port, dout_26_port, dout_25_port, dout_24_port, 
      dout_23_port, dout_22_port, dout_21_port, dout_20_port, dout_19_port, 
      dout_18_port, dout_17_port, dout_16_port, dout_15_port, dout_14_port, 
      dout_13_port, dout_12_port, dout_11_port, dout_10_port, dout_9_port, 
      dout_8_port, dout_7_port, dout_6_port, dout_5_port, dout_4_port, 
      dout_3_port, dout_2_port, dout_1_port, dout_0_port, n129, n130, n131, 
      n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, 
      n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, 
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n1, n2, n3, n4, n5, n6, net108745, net108746, net108747, net108748,
      net108749, net108750, net108751, net108752, net108753, net108754, 
      net108755, net108756, net108757, net108758, net108759, net108760, 
      net108761, net108762, net108763, net108764, net108765, net108766, 
      net108767, net108768, net108769, net108770, net108771, net108772, 
      net108773, net108774, net108775, net108776, net108777, net108778, 
      net108779, net108780, net108781, net108782, net108783, net108784, 
      net108785, net108786, net108787, net108788, net108789, net108790, 
      net108791, net108792, net108793, net108794, net108795, net108796, 
      net108797, net108798, net108799, net108800, net108801, net108802, 
      net108803, net108804, net108805, net108806, net108807, net108808 : 
      std_logic;

begin
   dout <= ( dout_63_port, dout_62_port, dout_61_port, dout_60_port, 
      dout_59_port, dout_58_port, dout_57_port, dout_56_port, dout_55_port, 
      dout_54_port, dout_53_port, dout_52_port, dout_51_port, dout_50_port, 
      dout_49_port, dout_48_port, dout_47_port, dout_46_port, dout_45_port, 
      dout_44_port, dout_43_port, dout_42_port, dout_41_port, dout_40_port, 
      dout_39_port, dout_38_port, dout_37_port, dout_36_port, dout_35_port, 
      dout_34_port, dout_33_port, dout_32_port, dout_31_port, dout_30_port, 
      dout_29_port, dout_28_port, dout_27_port, dout_26_port, dout_25_port, 
      dout_24_port, dout_23_port, dout_22_port, dout_21_port, dout_20_port, 
      dout_19_port, dout_18_port, dout_17_port, dout_16_port, dout_15_port, 
      dout_14_port, dout_13_port, dout_12_port, dout_11_port, dout_10_port, 
      dout_9_port, dout_8_port, dout_7_port, dout_6_port, dout_5_port, 
      dout_4_port, dout_3_port, dout_2_port, dout_1_port, dout_0_port );
   
   dout_reg_63_inst : DFFR_X1 port map( D => n192, CK => clk, RN => rst, Q => 
                           dout_63_port, QN => net108808);
   dout_reg_62_inst : DFFR_X1 port map( D => n191, CK => clk, RN => rst, Q => 
                           dout_62_port, QN => net108807);
   dout_reg_61_inst : DFFR_X1 port map( D => n190, CK => clk, RN => rst, Q => 
                           dout_61_port, QN => net108806);
   dout_reg_60_inst : DFFR_X1 port map( D => n189, CK => clk, RN => rst, Q => 
                           dout_60_port, QN => net108805);
   dout_reg_59_inst : DFFR_X1 port map( D => n188, CK => clk, RN => rst, Q => 
                           dout_59_port, QN => net108804);
   dout_reg_58_inst : DFFR_X1 port map( D => n187, CK => clk, RN => rst, Q => 
                           dout_58_port, QN => net108803);
   dout_reg_57_inst : DFFR_X1 port map( D => n186, CK => clk, RN => rst, Q => 
                           dout_57_port, QN => net108802);
   dout_reg_56_inst : DFFR_X1 port map( D => n185, CK => clk, RN => rst, Q => 
                           dout_56_port, QN => net108801);
   dout_reg_55_inst : DFFR_X1 port map( D => n184, CK => clk, RN => rst, Q => 
                           dout_55_port, QN => net108800);
   dout_reg_54_inst : DFFR_X1 port map( D => n183, CK => clk, RN => rst, Q => 
                           dout_54_port, QN => net108799);
   dout_reg_53_inst : DFFR_X1 port map( D => n182, CK => clk, RN => rst, Q => 
                           dout_53_port, QN => net108798);
   dout_reg_52_inst : DFFR_X1 port map( D => n181, CK => clk, RN => rst, Q => 
                           dout_52_port, QN => net108797);
   dout_reg_51_inst : DFFR_X1 port map( D => n180, CK => clk, RN => rst, Q => 
                           dout_51_port, QN => net108796);
   dout_reg_50_inst : DFFR_X1 port map( D => n179, CK => clk, RN => rst, Q => 
                           dout_50_port, QN => net108795);
   dout_reg_49_inst : DFFR_X1 port map( D => n178, CK => clk, RN => rst, Q => 
                           dout_49_port, QN => net108794);
   dout_reg_48_inst : DFFR_X1 port map( D => n177, CK => clk, RN => rst, Q => 
                           dout_48_port, QN => net108793);
   dout_reg_47_inst : DFFR_X1 port map( D => n176, CK => clk, RN => rst, Q => 
                           dout_47_port, QN => net108792);
   dout_reg_46_inst : DFFR_X1 port map( D => n175, CK => clk, RN => rst, Q => 
                           dout_46_port, QN => net108791);
   dout_reg_45_inst : DFFR_X1 port map( D => n174, CK => clk, RN => rst, Q => 
                           dout_45_port, QN => net108790);
   dout_reg_44_inst : DFFR_X1 port map( D => n173, CK => clk, RN => rst, Q => 
                           dout_44_port, QN => net108789);
   dout_reg_43_inst : DFFR_X1 port map( D => n172, CK => clk, RN => rst, Q => 
                           dout_43_port, QN => net108788);
   dout_reg_42_inst : DFFR_X1 port map( D => n171, CK => clk, RN => rst, Q => 
                           dout_42_port, QN => net108787);
   dout_reg_41_inst : DFFR_X1 port map( D => n170, CK => clk, RN => rst, Q => 
                           dout_41_port, QN => net108786);
   dout_reg_40_inst : DFFR_X1 port map( D => n169, CK => clk, RN => rst, Q => 
                           dout_40_port, QN => net108785);
   dout_reg_39_inst : DFFR_X1 port map( D => n168, CK => clk, RN => rst, Q => 
                           dout_39_port, QN => net108784);
   dout_reg_38_inst : DFFR_X1 port map( D => n167, CK => clk, RN => rst, Q => 
                           dout_38_port, QN => net108783);
   dout_reg_37_inst : DFFR_X1 port map( D => n166, CK => clk, RN => rst, Q => 
                           dout_37_port, QN => net108782);
   dout_reg_36_inst : DFFR_X1 port map( D => n165, CK => clk, RN => rst, Q => 
                           dout_36_port, QN => net108781);
   dout_reg_35_inst : DFFR_X1 port map( D => n164, CK => clk, RN => rst, Q => 
                           dout_35_port, QN => net108780);
   dout_reg_34_inst : DFFR_X1 port map( D => n163, CK => clk, RN => rst, Q => 
                           dout_34_port, QN => net108779);
   dout_reg_33_inst : DFFR_X1 port map( D => n162, CK => clk, RN => rst, Q => 
                           dout_33_port, QN => net108778);
   dout_reg_32_inst : DFFR_X1 port map( D => n161, CK => clk, RN => rst, Q => 
                           dout_32_port, QN => net108777);
   dout_reg_31_inst : DFFR_X1 port map( D => n160, CK => clk, RN => rst, Q => 
                           dout_31_port, QN => net108776);
   dout_reg_30_inst : DFFR_X1 port map( D => n159, CK => clk, RN => rst, Q => 
                           dout_30_port, QN => net108775);
   dout_reg_29_inst : DFFR_X1 port map( D => n158, CK => clk, RN => rst, Q => 
                           dout_29_port, QN => net108774);
   dout_reg_28_inst : DFFR_X1 port map( D => n157, CK => clk, RN => rst, Q => 
                           dout_28_port, QN => net108773);
   dout_reg_27_inst : DFFR_X1 port map( D => n156, CK => clk, RN => rst, Q => 
                           dout_27_port, QN => net108772);
   dout_reg_26_inst : DFFR_X1 port map( D => n155, CK => clk, RN => rst, Q => 
                           dout_26_port, QN => net108771);
   dout_reg_25_inst : DFFR_X1 port map( D => n154, CK => clk, RN => rst, Q => 
                           dout_25_port, QN => net108770);
   dout_reg_24_inst : DFFR_X1 port map( D => n153, CK => clk, RN => rst, Q => 
                           dout_24_port, QN => net108769);
   dout_reg_23_inst : DFFR_X1 port map( D => n152, CK => clk, RN => rst, Q => 
                           dout_23_port, QN => net108768);
   dout_reg_22_inst : DFFR_X1 port map( D => n151, CK => clk, RN => rst, Q => 
                           dout_22_port, QN => net108767);
   dout_reg_21_inst : DFFR_X1 port map( D => n150, CK => clk, RN => rst, Q => 
                           dout_21_port, QN => net108766);
   dout_reg_20_inst : DFFR_X1 port map( D => n149, CK => clk, RN => rst, Q => 
                           dout_20_port, QN => net108765);
   dout_reg_19_inst : DFFR_X1 port map( D => n148, CK => clk, RN => rst, Q => 
                           dout_19_port, QN => net108764);
   dout_reg_18_inst : DFFR_X1 port map( D => n147, CK => clk, RN => rst, Q => 
                           dout_18_port, QN => net108763);
   dout_reg_17_inst : DFFR_X1 port map( D => n146, CK => clk, RN => rst, Q => 
                           dout_17_port, QN => net108762);
   dout_reg_16_inst : DFFR_X1 port map( D => n145, CK => clk, RN => rst, Q => 
                           dout_16_port, QN => net108761);
   dout_reg_15_inst : DFFR_X1 port map( D => n144, CK => clk, RN => rst, Q => 
                           dout_15_port, QN => net108760);
   dout_reg_14_inst : DFFR_X1 port map( D => n143, CK => clk, RN => rst, Q => 
                           dout_14_port, QN => net108759);
   dout_reg_13_inst : DFFR_X1 port map( D => n142, CK => clk, RN => rst, Q => 
                           dout_13_port, QN => net108758);
   dout_reg_12_inst : DFFR_X1 port map( D => n141, CK => clk, RN => rst, Q => 
                           dout_12_port, QN => net108757);
   dout_reg_11_inst : DFFR_X1 port map( D => n140, CK => clk, RN => rst, Q => 
                           dout_11_port, QN => net108756);
   dout_reg_10_inst : DFFR_X1 port map( D => n139, CK => clk, RN => rst, Q => 
                           dout_10_port, QN => net108755);
   dout_reg_9_inst : DFFR_X1 port map( D => n138, CK => clk, RN => rst, Q => 
                           dout_9_port, QN => net108754);
   dout_reg_8_inst : DFFR_X1 port map( D => n137, CK => clk, RN => rst, Q => 
                           dout_8_port, QN => net108753);
   dout_reg_7_inst : DFFR_X1 port map( D => n136, CK => clk, RN => rst, Q => 
                           dout_7_port, QN => net108752);
   dout_reg_6_inst : DFFR_X1 port map( D => n135, CK => clk, RN => rst, Q => 
                           dout_6_port, QN => net108751);
   dout_reg_5_inst : DFFR_X1 port map( D => n134, CK => clk, RN => rst, Q => 
                           dout_5_port, QN => net108750);
   dout_reg_4_inst : DFFR_X1 port map( D => n133, CK => clk, RN => rst, Q => 
                           dout_4_port, QN => net108749);
   dout_reg_3_inst : DFFR_X1 port map( D => n132, CK => clk, RN => rst, Q => 
                           dout_3_port, QN => net108748);
   dout_reg_2_inst : DFFR_X1 port map( D => n131, CK => clk, RN => rst, Q => 
                           dout_2_port, QN => net108747);
   dout_reg_1_inst : DFFR_X1 port map( D => n130, CK => clk, RN => rst, Q => 
                           dout_1_port, QN => net108746);
   dout_reg_0_inst : DFFR_X1 port map( D => n129, CK => clk, RN => rst, Q => 
                           dout_0_port, QN => net108745);
   U2 : CLKBUF_X1 port map( A => en, Z => n1);
   U3 : CLKBUF_X1 port map( A => en, Z => n2);
   U4 : CLKBUF_X1 port map( A => en, Z => n3);
   U5 : CLKBUF_X1 port map( A => en, Z => n4);
   U6 : CLKBUF_X1 port map( A => en, Z => n5);
   U7 : CLKBUF_X1 port map( A => en, Z => n6);
   U8 : MUX2_X1 port map( A => dout_63_port, B => din(63), S => n1, Z => n192);
   U9 : MUX2_X1 port map( A => dout_62_port, B => din(62), S => n1, Z => n191);
   U10 : MUX2_X1 port map( A => dout_61_port, B => din(61), S => n1, Z => n190)
                           ;
   U11 : MUX2_X1 port map( A => dout_60_port, B => din(60), S => n1, Z => n189)
                           ;
   U12 : MUX2_X1 port map( A => dout_59_port, B => din(59), S => n1, Z => n188)
                           ;
   U13 : MUX2_X1 port map( A => dout_58_port, B => din(58), S => n1, Z => n187)
                           ;
   U14 : MUX2_X1 port map( A => dout_57_port, B => din(57), S => n1, Z => n186)
                           ;
   U15 : MUX2_X1 port map( A => dout_56_port, B => din(56), S => n1, Z => n185)
                           ;
   U16 : MUX2_X1 port map( A => dout_55_port, B => din(55), S => n1, Z => n184)
                           ;
   U17 : MUX2_X1 port map( A => dout_54_port, B => din(54), S => n1, Z => n183)
                           ;
   U18 : MUX2_X1 port map( A => dout_53_port, B => din(53), S => n1, Z => n182)
                           ;
   U19 : MUX2_X1 port map( A => dout_52_port, B => din(52), S => n1, Z => n181)
                           ;
   U20 : MUX2_X1 port map( A => dout_51_port, B => din(51), S => n2, Z => n180)
                           ;
   U21 : MUX2_X1 port map( A => dout_50_port, B => din(50), S => n2, Z => n179)
                           ;
   U22 : MUX2_X1 port map( A => dout_49_port, B => din(49), S => n2, Z => n178)
                           ;
   U23 : MUX2_X1 port map( A => dout_48_port, B => din(48), S => n2, Z => n177)
                           ;
   U24 : MUX2_X1 port map( A => dout_47_port, B => din(47), S => n2, Z => n176)
                           ;
   U25 : MUX2_X1 port map( A => dout_46_port, B => din(46), S => n2, Z => n175)
                           ;
   U26 : MUX2_X1 port map( A => dout_45_port, B => din(45), S => n2, Z => n174)
                           ;
   U27 : MUX2_X1 port map( A => dout_44_port, B => din(44), S => n2, Z => n173)
                           ;
   U28 : MUX2_X1 port map( A => dout_43_port, B => din(43), S => n2, Z => n172)
                           ;
   U29 : MUX2_X1 port map( A => dout_42_port, B => din(42), S => n2, Z => n171)
                           ;
   U30 : MUX2_X1 port map( A => dout_41_port, B => din(41), S => n2, Z => n170)
                           ;
   U31 : MUX2_X1 port map( A => dout_40_port, B => din(40), S => n2, Z => n169)
                           ;
   U32 : MUX2_X1 port map( A => dout_39_port, B => din(39), S => n3, Z => n168)
                           ;
   U33 : MUX2_X1 port map( A => dout_38_port, B => din(38), S => n3, Z => n167)
                           ;
   U34 : MUX2_X1 port map( A => dout_37_port, B => din(37), S => n3, Z => n166)
                           ;
   U35 : MUX2_X1 port map( A => dout_36_port, B => din(36), S => n3, Z => n165)
                           ;
   U36 : MUX2_X1 port map( A => dout_35_port, B => din(35), S => n3, Z => n164)
                           ;
   U37 : MUX2_X1 port map( A => dout_34_port, B => din(34), S => n3, Z => n163)
                           ;
   U38 : MUX2_X1 port map( A => dout_33_port, B => din(33), S => n3, Z => n162)
                           ;
   U39 : MUX2_X1 port map( A => dout_32_port, B => din(32), S => n3, Z => n161)
                           ;
   U40 : MUX2_X1 port map( A => dout_31_port, B => din(31), S => n3, Z => n160)
                           ;
   U41 : MUX2_X1 port map( A => dout_30_port, B => din(30), S => n3, Z => n159)
                           ;
   U42 : MUX2_X1 port map( A => dout_29_port, B => din(29), S => n3, Z => n158)
                           ;
   U43 : MUX2_X1 port map( A => dout_28_port, B => din(28), S => n3, Z => n157)
                           ;
   U44 : MUX2_X1 port map( A => dout_27_port, B => din(27), S => n4, Z => n156)
                           ;
   U45 : MUX2_X1 port map( A => dout_26_port, B => din(26), S => n4, Z => n155)
                           ;
   U46 : MUX2_X1 port map( A => dout_25_port, B => din(25), S => n4, Z => n154)
                           ;
   U47 : MUX2_X1 port map( A => dout_24_port, B => din(24), S => n4, Z => n153)
                           ;
   U48 : MUX2_X1 port map( A => dout_23_port, B => din(23), S => n4, Z => n152)
                           ;
   U49 : MUX2_X1 port map( A => dout_22_port, B => din(22), S => n4, Z => n151)
                           ;
   U50 : MUX2_X1 port map( A => dout_21_port, B => din(21), S => n4, Z => n150)
                           ;
   U51 : MUX2_X1 port map( A => dout_20_port, B => din(20), S => n4, Z => n149)
                           ;
   U52 : MUX2_X1 port map( A => dout_19_port, B => din(19), S => n4, Z => n148)
                           ;
   U53 : MUX2_X1 port map( A => dout_18_port, B => din(18), S => n4, Z => n147)
                           ;
   U54 : MUX2_X1 port map( A => dout_17_port, B => din(17), S => n4, Z => n146)
                           ;
   U55 : MUX2_X1 port map( A => dout_16_port, B => din(16), S => n4, Z => n145)
                           ;
   U56 : MUX2_X1 port map( A => dout_15_port, B => din(15), S => n5, Z => n144)
                           ;
   U57 : MUX2_X1 port map( A => dout_14_port, B => din(14), S => n5, Z => n143)
                           ;
   U58 : MUX2_X1 port map( A => dout_13_port, B => din(13), S => n5, Z => n142)
                           ;
   U59 : MUX2_X1 port map( A => dout_12_port, B => din(12), S => n5, Z => n141)
                           ;
   U60 : MUX2_X1 port map( A => dout_11_port, B => din(11), S => n5, Z => n140)
                           ;
   U61 : MUX2_X1 port map( A => dout_10_port, B => din(10), S => n5, Z => n139)
                           ;
   U62 : MUX2_X1 port map( A => dout_9_port, B => din(9), S => n5, Z => n138);
   U63 : MUX2_X1 port map( A => dout_8_port, B => din(8), S => n5, Z => n137);
   U64 : MUX2_X1 port map( A => dout_7_port, B => din(7), S => n5, Z => n136);
   U65 : MUX2_X1 port map( A => dout_6_port, B => din(6), S => n5, Z => n135);
   U66 : MUX2_X1 port map( A => dout_5_port, B => din(5), S => n5, Z => n134);
   U67 : MUX2_X1 port map( A => dout_4_port, B => din(4), S => n5, Z => n133);
   U68 : MUX2_X1 port map( A => dout_3_port, B => din(3), S => n6, Z => n132);
   U69 : MUX2_X1 port map( A => dout_2_port, B => din(2), S => n6, Z => n131);
   U70 : MUX2_X1 port map( A => dout_1_port, B => din(1), S => n6, Z => n130);
   U71 : MUX2_X1 port map( A => dout_0_port, B => din(0), S => n6, Z => n129);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AddSub_DATA_SIZE64 is

   port( as : in std_logic;  a, b : in std_logic_vector (63 downto 0);  re : 
         out std_logic_vector (63 downto 0);  cout : out std_logic);

end AddSub_DATA_SIZE64;

architecture SYN_add_sub_arch of AddSub_DATA_SIZE64 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component Adder_DATA_SIZE64
      port( cin : in std_logic;  a, b : in std_logic_vector (63 downto 0);  s :
            out std_logic_vector (63 downto 0);  cout : out std_logic);
   end component;
   
   signal b_new_63_port, b_new_62_port, b_new_61_port, b_new_60_port, 
      b_new_59_port, b_new_58_port, b_new_57_port, b_new_56_port, b_new_55_port
      , b_new_54_port, b_new_53_port, b_new_52_port, b_new_51_port, 
      b_new_50_port, b_new_49_port, b_new_48_port, b_new_47_port, b_new_46_port
      , b_new_45_port, b_new_44_port, b_new_43_port, b_new_42_port, 
      b_new_41_port, b_new_40_port, b_new_39_port, b_new_38_port, b_new_37_port
      , b_new_36_port, b_new_35_port, b_new_34_port, b_new_33_port, 
      b_new_32_port, b_new_31_port, b_new_30_port, b_new_29_port, b_new_28_port
      , b_new_27_port, b_new_26_port, b_new_25_port, b_new_24_port, 
      b_new_23_port, b_new_22_port, b_new_21_port, b_new_20_port, b_new_19_port
      , b_new_18_port, b_new_17_port, b_new_16_port, b_new_15_port, 
      b_new_14_port, b_new_13_port, b_new_12_port, b_new_11_port, b_new_10_port
      , b_new_9_port, b_new_8_port, b_new_7_port, b_new_6_port, b_new_5_port, 
      b_new_4_port, b_new_3_port, b_new_2_port, b_new_1_port, b_new_0_port : 
      std_logic;

begin
   
   ADDER0 : Adder_DATA_SIZE64 port map( cin => as, a(63) => a(63), a(62) => 
                           a(62), a(61) => a(61), a(60) => a(60), a(59) => 
                           a(59), a(58) => a(58), a(57) => a(57), a(56) => 
                           a(56), a(55) => a(55), a(54) => a(54), a(53) => 
                           a(53), a(52) => a(52), a(51) => a(51), a(50) => 
                           a(50), a(49) => a(49), a(48) => a(48), a(47) => 
                           a(47), a(46) => a(46), a(45) => a(45), a(44) => 
                           a(44), a(43) => a(43), a(42) => a(42), a(41) => 
                           a(41), a(40) => a(40), a(39) => a(39), a(38) => 
                           a(38), a(37) => a(37), a(36) => a(36), a(35) => 
                           a(35), a(34) => a(34), a(33) => a(33), a(32) => 
                           a(32), a(31) => a(31), a(30) => a(30), a(29) => 
                           a(29), a(28) => a(28), a(27) => a(27), a(26) => 
                           a(26), a(25) => a(25), a(24) => a(24), a(23) => 
                           a(23), a(22) => a(22), a(21) => a(21), a(20) => 
                           a(20), a(19) => a(19), a(18) => a(18), a(17) => 
                           a(17), a(16) => a(16), a(15) => a(15), a(14) => 
                           a(14), a(13) => a(13), a(12) => a(12), a(11) => 
                           a(11), a(10) => a(10), a(9) => a(9), a(8) => a(8), 
                           a(7) => a(7), a(6) => a(6), a(5) => a(5), a(4) => 
                           a(4), a(3) => a(3), a(2) => a(2), a(1) => a(1), a(0)
                           => a(0), b(63) => b_new_63_port, b(62) => 
                           b_new_62_port, b(61) => b_new_61_port, b(60) => 
                           b_new_60_port, b(59) => b_new_59_port, b(58) => 
                           b_new_58_port, b(57) => b_new_57_port, b(56) => 
                           b_new_56_port, b(55) => b_new_55_port, b(54) => 
                           b_new_54_port, b(53) => b_new_53_port, b(52) => 
                           b_new_52_port, b(51) => b_new_51_port, b(50) => 
                           b_new_50_port, b(49) => b_new_49_port, b(48) => 
                           b_new_48_port, b(47) => b_new_47_port, b(46) => 
                           b_new_46_port, b(45) => b_new_45_port, b(44) => 
                           b_new_44_port, b(43) => b_new_43_port, b(42) => 
                           b_new_42_port, b(41) => b_new_41_port, b(40) => 
                           b_new_40_port, b(39) => b_new_39_port, b(38) => 
                           b_new_38_port, b(37) => b_new_37_port, b(36) => 
                           b_new_36_port, b(35) => b_new_35_port, b(34) => 
                           b_new_34_port, b(33) => b_new_33_port, b(32) => 
                           b_new_32_port, b(31) => b_new_31_port, b(30) => 
                           b_new_30_port, b(29) => b_new_29_port, b(28) => 
                           b_new_28_port, b(27) => b_new_27_port, b(26) => 
                           b_new_26_port, b(25) => b_new_25_port, b(24) => 
                           b_new_24_port, b(23) => b_new_23_port, b(22) => 
                           b_new_22_port, b(21) => b_new_21_port, b(20) => 
                           b_new_20_port, b(19) => b_new_19_port, b(18) => 
                           b_new_18_port, b(17) => b_new_17_port, b(16) => 
                           b_new_16_port, b(15) => b_new_15_port, b(14) => 
                           b_new_14_port, b(13) => b_new_13_port, b(12) => 
                           b_new_12_port, b(11) => b_new_11_port, b(10) => 
                           b_new_10_port, b(9) => b_new_9_port, b(8) => 
                           b_new_8_port, b(7) => b_new_7_port, b(6) => 
                           b_new_6_port, b(5) => b_new_5_port, b(4) => 
                           b_new_4_port, b(3) => b_new_3_port, b(2) => 
                           b_new_2_port, b(1) => b_new_1_port, b(0) => 
                           b_new_0_port, s(63) => re(63), s(62) => re(62), 
                           s(61) => re(61), s(60) => re(60), s(59) => re(59), 
                           s(58) => re(58), s(57) => re(57), s(56) => re(56), 
                           s(55) => re(55), s(54) => re(54), s(53) => re(53), 
                           s(52) => re(52), s(51) => re(51), s(50) => re(50), 
                           s(49) => re(49), s(48) => re(48), s(47) => re(47), 
                           s(46) => re(46), s(45) => re(45), s(44) => re(44), 
                           s(43) => re(43), s(42) => re(42), s(41) => re(41), 
                           s(40) => re(40), s(39) => re(39), s(38) => re(38), 
                           s(37) => re(37), s(36) => re(36), s(35) => re(35), 
                           s(34) => re(34), s(33) => re(33), s(32) => re(32), 
                           s(31) => re(31), s(30) => re(30), s(29) => re(29), 
                           s(28) => re(28), s(27) => re(27), s(26) => re(26), 
                           s(25) => re(25), s(24) => re(24), s(23) => re(23), 
                           s(22) => re(22), s(21) => re(21), s(20) => re(20), 
                           s(19) => re(19), s(18) => re(18), s(17) => re(17), 
                           s(16) => re(16), s(15) => re(15), s(14) => re(14), 
                           s(13) => re(13), s(12) => re(12), s(11) => re(11), 
                           s(10) => re(10), s(9) => re(9), s(8) => re(8), s(7) 
                           => re(7), s(6) => re(6), s(5) => re(5), s(4) => 
                           re(4), s(3) => re(3), s(2) => re(2), s(1) => re(1), 
                           s(0) => re(0), cout => cout);
   U1 : XOR2_X1 port map( A => b(9), B => as, Z => b_new_9_port);
   U2 : XOR2_X1 port map( A => b(8), B => as, Z => b_new_8_port);
   U3 : XOR2_X1 port map( A => b(7), B => as, Z => b_new_7_port);
   U4 : XOR2_X1 port map( A => b(6), B => as, Z => b_new_6_port);
   U5 : XOR2_X1 port map( A => b(63), B => as, Z => b_new_63_port);
   U6 : XOR2_X1 port map( A => b(62), B => as, Z => b_new_62_port);
   U7 : XOR2_X1 port map( A => b(61), B => as, Z => b_new_61_port);
   U8 : XOR2_X1 port map( A => b(60), B => as, Z => b_new_60_port);
   U9 : XOR2_X1 port map( A => b(5), B => as, Z => b_new_5_port);
   U10 : XOR2_X1 port map( A => b(59), B => as, Z => b_new_59_port);
   U11 : XOR2_X1 port map( A => b(58), B => as, Z => b_new_58_port);
   U12 : XOR2_X1 port map( A => b(57), B => as, Z => b_new_57_port);
   U13 : XOR2_X1 port map( A => b(56), B => as, Z => b_new_56_port);
   U14 : XOR2_X1 port map( A => b(55), B => as, Z => b_new_55_port);
   U15 : XOR2_X1 port map( A => b(54), B => as, Z => b_new_54_port);
   U16 : XOR2_X1 port map( A => b(53), B => as, Z => b_new_53_port);
   U17 : XOR2_X1 port map( A => b(52), B => as, Z => b_new_52_port);
   U18 : XOR2_X1 port map( A => b(51), B => as, Z => b_new_51_port);
   U19 : XOR2_X1 port map( A => b(50), B => as, Z => b_new_50_port);
   U20 : XOR2_X1 port map( A => b(4), B => as, Z => b_new_4_port);
   U21 : XOR2_X1 port map( A => b(49), B => as, Z => b_new_49_port);
   U22 : XOR2_X1 port map( A => b(48), B => as, Z => b_new_48_port);
   U23 : XOR2_X1 port map( A => b(47), B => as, Z => b_new_47_port);
   U24 : XOR2_X1 port map( A => b(46), B => as, Z => b_new_46_port);
   U25 : XOR2_X1 port map( A => b(45), B => as, Z => b_new_45_port);
   U26 : XOR2_X1 port map( A => b(44), B => as, Z => b_new_44_port);
   U27 : XOR2_X1 port map( A => b(43), B => as, Z => b_new_43_port);
   U28 : XOR2_X1 port map( A => b(42), B => as, Z => b_new_42_port);
   U29 : XOR2_X1 port map( A => b(41), B => as, Z => b_new_41_port);
   U30 : XOR2_X1 port map( A => b(40), B => as, Z => b_new_40_port);
   U31 : XOR2_X1 port map( A => b(3), B => as, Z => b_new_3_port);
   U32 : XOR2_X1 port map( A => b(39), B => as, Z => b_new_39_port);
   U33 : XOR2_X1 port map( A => b(38), B => as, Z => b_new_38_port);
   U34 : XOR2_X1 port map( A => b(37), B => as, Z => b_new_37_port);
   U35 : XOR2_X1 port map( A => b(36), B => as, Z => b_new_36_port);
   U36 : XOR2_X1 port map( A => b(35), B => as, Z => b_new_35_port);
   U37 : XOR2_X1 port map( A => b(34), B => as, Z => b_new_34_port);
   U38 : XOR2_X1 port map( A => b(33), B => as, Z => b_new_33_port);
   U39 : XOR2_X1 port map( A => b(32), B => as, Z => b_new_32_port);
   U40 : XOR2_X1 port map( A => b(31), B => as, Z => b_new_31_port);
   U41 : XOR2_X1 port map( A => b(30), B => as, Z => b_new_30_port);
   U42 : XOR2_X1 port map( A => b(2), B => as, Z => b_new_2_port);
   U43 : XOR2_X1 port map( A => b(29), B => as, Z => b_new_29_port);
   U44 : XOR2_X1 port map( A => b(28), B => as, Z => b_new_28_port);
   U45 : XOR2_X1 port map( A => b(27), B => as, Z => b_new_27_port);
   U46 : XOR2_X1 port map( A => b(26), B => as, Z => b_new_26_port);
   U47 : XOR2_X1 port map( A => b(25), B => as, Z => b_new_25_port);
   U48 : XOR2_X1 port map( A => b(24), B => as, Z => b_new_24_port);
   U49 : XOR2_X1 port map( A => b(23), B => as, Z => b_new_23_port);
   U50 : XOR2_X1 port map( A => b(22), B => as, Z => b_new_22_port);
   U51 : XOR2_X1 port map( A => b(21), B => as, Z => b_new_21_port);
   U52 : XOR2_X1 port map( A => b(20), B => as, Z => b_new_20_port);
   U53 : XOR2_X1 port map( A => b(1), B => as, Z => b_new_1_port);
   U54 : XOR2_X1 port map( A => b(19), B => as, Z => b_new_19_port);
   U55 : XOR2_X1 port map( A => b(18), B => as, Z => b_new_18_port);
   U56 : XOR2_X1 port map( A => b(17), B => as, Z => b_new_17_port);
   U57 : XOR2_X1 port map( A => b(16), B => as, Z => b_new_16_port);
   U58 : XOR2_X1 port map( A => b(15), B => as, Z => b_new_15_port);
   U59 : XOR2_X1 port map( A => b(14), B => as, Z => b_new_14_port);
   U60 : XOR2_X1 port map( A => b(13), B => as, Z => b_new_13_port);
   U61 : XOR2_X1 port map( A => b(12), B => as, Z => b_new_12_port);
   U62 : XOR2_X1 port map( A => b(11), B => as, Z => b_new_11_port);
   U63 : XOR2_X1 port map( A => b(10), B => as, Z => b_new_10_port);
   U64 : XOR2_X1 port map( A => b(0), B => as, Z => b_new_0_port);

end SYN_add_sub_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE64 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (63 downto 0);  
         dout : out std_logic_vector (63 downto 0));

end Mux_DATA_SIZE64;

architecture SYN_mux_arch of Mux_DATA_SIZE64 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(9), B => din1(9), S => sel, Z => dout(9));
   U2 : MUX2_X1 port map( A => din0(8), B => din1(8), S => sel, Z => dout(8));
   U3 : MUX2_X1 port map( A => din0(7), B => din1(7), S => sel, Z => dout(7));
   U4 : MUX2_X1 port map( A => din0(6), B => din1(6), S => sel, Z => dout(6));
   U5 : MUX2_X1 port map( A => din0(63), B => din1(63), S => sel, Z => dout(63)
                           );
   U6 : MUX2_X1 port map( A => din0(62), B => din1(62), S => sel, Z => dout(62)
                           );
   U7 : MUX2_X1 port map( A => din0(61), B => din1(61), S => sel, Z => dout(61)
                           );
   U8 : MUX2_X1 port map( A => din0(60), B => din1(60), S => sel, Z => dout(60)
                           );
   U9 : MUX2_X1 port map( A => din0(5), B => din1(5), S => sel, Z => dout(5));
   U10 : MUX2_X1 port map( A => din0(59), B => din1(59), S => sel, Z => 
                           dout(59));
   U11 : MUX2_X1 port map( A => din0(58), B => din1(58), S => sel, Z => 
                           dout(58));
   U12 : MUX2_X1 port map( A => din0(57), B => din1(57), S => sel, Z => 
                           dout(57));
   U13 : MUX2_X1 port map( A => din0(56), B => din1(56), S => sel, Z => 
                           dout(56));
   U14 : MUX2_X1 port map( A => din0(55), B => din1(55), S => sel, Z => 
                           dout(55));
   U15 : MUX2_X1 port map( A => din0(54), B => din1(54), S => sel, Z => 
                           dout(54));
   U16 : MUX2_X1 port map( A => din0(53), B => din1(53), S => sel, Z => 
                           dout(53));
   U17 : MUX2_X1 port map( A => din0(52), B => din1(52), S => sel, Z => 
                           dout(52));
   U18 : MUX2_X1 port map( A => din0(51), B => din1(51), S => sel, Z => 
                           dout(51));
   U19 : MUX2_X1 port map( A => din0(50), B => din1(50), S => sel, Z => 
                           dout(50));
   U20 : MUX2_X1 port map( A => din0(4), B => din1(4), S => sel, Z => dout(4));
   U21 : MUX2_X1 port map( A => din0(49), B => din1(49), S => sel, Z => 
                           dout(49));
   U22 : MUX2_X1 port map( A => din0(48), B => din1(48), S => sel, Z => 
                           dout(48));
   U23 : MUX2_X1 port map( A => din0(47), B => din1(47), S => sel, Z => 
                           dout(47));
   U24 : MUX2_X1 port map( A => din0(46), B => din1(46), S => sel, Z => 
                           dout(46));
   U25 : MUX2_X1 port map( A => din0(45), B => din1(45), S => sel, Z => 
                           dout(45));
   U26 : MUX2_X1 port map( A => din0(44), B => din1(44), S => sel, Z => 
                           dout(44));
   U27 : MUX2_X1 port map( A => din0(43), B => din1(43), S => sel, Z => 
                           dout(43));
   U28 : MUX2_X1 port map( A => din0(42), B => din1(42), S => sel, Z => 
                           dout(42));
   U29 : MUX2_X1 port map( A => din0(41), B => din1(41), S => sel, Z => 
                           dout(41));
   U30 : MUX2_X1 port map( A => din0(40), B => din1(40), S => sel, Z => 
                           dout(40));
   U31 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U32 : MUX2_X1 port map( A => din0(39), B => din1(39), S => sel, Z => 
                           dout(39));
   U33 : MUX2_X1 port map( A => din0(38), B => din1(38), S => sel, Z => 
                           dout(38));
   U34 : MUX2_X1 port map( A => din0(37), B => din1(37), S => sel, Z => 
                           dout(37));
   U35 : MUX2_X1 port map( A => din0(36), B => din1(36), S => sel, Z => 
                           dout(36));
   U36 : MUX2_X1 port map( A => din0(35), B => din1(35), S => sel, Z => 
                           dout(35));
   U37 : MUX2_X1 port map( A => din0(34), B => din1(34), S => sel, Z => 
                           dout(34));
   U38 : MUX2_X1 port map( A => din0(33), B => din1(33), S => sel, Z => 
                           dout(33));
   U39 : MUX2_X1 port map( A => din0(32), B => din1(32), S => sel, Z => 
                           dout(32));
   U40 : MUX2_X1 port map( A => din0(31), B => din1(31), S => sel, Z => 
                           dout(31));
   U41 : MUX2_X1 port map( A => din0(30), B => din1(30), S => sel, Z => 
                           dout(30));
   U42 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U43 : MUX2_X1 port map( A => din0(29), B => din1(29), S => sel, Z => 
                           dout(29));
   U44 : MUX2_X1 port map( A => din0(28), B => din1(28), S => sel, Z => 
                           dout(28));
   U45 : MUX2_X1 port map( A => din0(27), B => din1(27), S => sel, Z => 
                           dout(27));
   U46 : MUX2_X1 port map( A => din0(26), B => din1(26), S => sel, Z => 
                           dout(26));
   U47 : MUX2_X1 port map( A => din0(25), B => din1(25), S => sel, Z => 
                           dout(25));
   U48 : MUX2_X1 port map( A => din0(24), B => din1(24), S => sel, Z => 
                           dout(24));
   U49 : MUX2_X1 port map( A => din0(23), B => din1(23), S => sel, Z => 
                           dout(23));
   U50 : MUX2_X1 port map( A => din0(22), B => din1(22), S => sel, Z => 
                           dout(22));
   U51 : MUX2_X1 port map( A => din0(21), B => din1(21), S => sel, Z => 
                           dout(21));
   U52 : MUX2_X1 port map( A => din0(20), B => din1(20), S => sel, Z => 
                           dout(20));
   U53 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U54 : MUX2_X1 port map( A => din0(19), B => din1(19), S => sel, Z => 
                           dout(19));
   U55 : MUX2_X1 port map( A => din0(18), B => din1(18), S => sel, Z => 
                           dout(18));
   U56 : MUX2_X1 port map( A => din0(17), B => din1(17), S => sel, Z => 
                           dout(17));
   U57 : MUX2_X1 port map( A => din0(16), B => din1(16), S => sel, Z => 
                           dout(16));
   U58 : MUX2_X1 port map( A => din0(15), B => din1(15), S => sel, Z => 
                           dout(15));
   U59 : MUX2_X1 port map( A => din0(14), B => din1(14), S => sel, Z => 
                           dout(14));
   U60 : MUX2_X1 port map( A => din0(13), B => din1(13), S => sel, Z => 
                           dout(13));
   U61 : MUX2_X1 port map( A => din0(12), B => din1(12), S => sel, Z => 
                           dout(12));
   U62 : MUX2_X1 port map( A => din0(11), B => din1(11), S => sel, Z => 
                           dout(11));
   U63 : MUX2_X1 port map( A => din0(10), B => din1(10), S => sel, Z => 
                           dout(10));
   U64 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity AddSub_DATA_SIZE32_0 is

   port( as : in std_logic;  a, b : in std_logic_vector (31 downto 0);  re : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end AddSub_DATA_SIZE32_0;

architecture SYN_add_sub_arch of AddSub_DATA_SIZE32_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component Adder_DATA_SIZE32_4
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;
   
   signal b_new_31_port, b_new_30_port, b_new_29_port, b_new_28_port, 
      b_new_27_port, b_new_26_port, b_new_25_port, b_new_24_port, b_new_23_port
      , b_new_22_port, b_new_21_port, b_new_20_port, b_new_19_port, 
      b_new_18_port, b_new_17_port, b_new_16_port, b_new_15_port, b_new_14_port
      , b_new_13_port, b_new_12_port, b_new_11_port, b_new_10_port, 
      b_new_9_port, b_new_8_port, b_new_7_port, b_new_6_port, b_new_5_port, 
      b_new_4_port, b_new_3_port, b_new_2_port, b_new_1_port, b_new_0_port : 
      std_logic;

begin
   
   ADDER0 : Adder_DATA_SIZE32_4 port map( cin => as, a(31) => a(31), a(30) => 
                           a(30), a(29) => a(29), a(28) => a(28), a(27) => 
                           a(27), a(26) => a(26), a(25) => a(25), a(24) => 
                           a(24), a(23) => a(23), a(22) => a(22), a(21) => 
                           a(21), a(20) => a(20), a(19) => a(19), a(18) => 
                           a(18), a(17) => a(17), a(16) => a(16), a(15) => 
                           a(15), a(14) => a(14), a(13) => a(13), a(12) => 
                           a(12), a(11) => a(11), a(10) => a(10), a(9) => a(9),
                           a(8) => a(8), a(7) => a(7), a(6) => a(6), a(5) => 
                           a(5), a(4) => a(4), a(3) => a(3), a(2) => a(2), a(1)
                           => a(1), a(0) => a(0), b(31) => b_new_31_port, b(30)
                           => b_new_30_port, b(29) => b_new_29_port, b(28) => 
                           b_new_28_port, b(27) => b_new_27_port, b(26) => 
                           b_new_26_port, b(25) => b_new_25_port, b(24) => 
                           b_new_24_port, b(23) => b_new_23_port, b(22) => 
                           b_new_22_port, b(21) => b_new_21_port, b(20) => 
                           b_new_20_port, b(19) => b_new_19_port, b(18) => 
                           b_new_18_port, b(17) => b_new_17_port, b(16) => 
                           b_new_16_port, b(15) => b_new_15_port, b(14) => 
                           b_new_14_port, b(13) => b_new_13_port, b(12) => 
                           b_new_12_port, b(11) => b_new_11_port, b(10) => 
                           b_new_10_port, b(9) => b_new_9_port, b(8) => 
                           b_new_8_port, b(7) => b_new_7_port, b(6) => 
                           b_new_6_port, b(5) => b_new_5_port, b(4) => 
                           b_new_4_port, b(3) => b_new_3_port, b(2) => 
                           b_new_2_port, b(1) => b_new_1_port, b(0) => 
                           b_new_0_port, s(31) => re(31), s(30) => re(30), 
                           s(29) => re(29), s(28) => re(28), s(27) => re(27), 
                           s(26) => re(26), s(25) => re(25), s(24) => re(24), 
                           s(23) => re(23), s(22) => re(22), s(21) => re(21), 
                           s(20) => re(20), s(19) => re(19), s(18) => re(18), 
                           s(17) => re(17), s(16) => re(16), s(15) => re(15), 
                           s(14) => re(14), s(13) => re(13), s(12) => re(12), 
                           s(11) => re(11), s(10) => re(10), s(9) => re(9), 
                           s(8) => re(8), s(7) => re(7), s(6) => re(6), s(5) =>
                           re(5), s(4) => re(4), s(3) => re(3), s(2) => re(2), 
                           s(1) => re(1), s(0) => re(0), cout => cout);
   U1 : XOR2_X1 port map( A => b(9), B => as, Z => b_new_9_port);
   U2 : XOR2_X1 port map( A => b(8), B => as, Z => b_new_8_port);
   U3 : XOR2_X1 port map( A => b(7), B => as, Z => b_new_7_port);
   U4 : XOR2_X1 port map( A => b(6), B => as, Z => b_new_6_port);
   U5 : XOR2_X1 port map( A => b(5), B => as, Z => b_new_5_port);
   U6 : XOR2_X1 port map( A => b(4), B => as, Z => b_new_4_port);
   U7 : XOR2_X1 port map( A => b(3), B => as, Z => b_new_3_port);
   U8 : XOR2_X1 port map( A => b(31), B => as, Z => b_new_31_port);
   U9 : XOR2_X1 port map( A => b(30), B => as, Z => b_new_30_port);
   U10 : XOR2_X1 port map( A => b(2), B => as, Z => b_new_2_port);
   U11 : XOR2_X1 port map( A => b(29), B => as, Z => b_new_29_port);
   U12 : XOR2_X1 port map( A => b(28), B => as, Z => b_new_28_port);
   U13 : XOR2_X1 port map( A => b(27), B => as, Z => b_new_27_port);
   U14 : XOR2_X1 port map( A => b(26), B => as, Z => b_new_26_port);
   U15 : XOR2_X1 port map( A => b(25), B => as, Z => b_new_25_port);
   U16 : XOR2_X1 port map( A => b(24), B => as, Z => b_new_24_port);
   U17 : XOR2_X1 port map( A => b(23), B => as, Z => b_new_23_port);
   U18 : XOR2_X1 port map( A => b(22), B => as, Z => b_new_22_port);
   U19 : XOR2_X1 port map( A => b(21), B => as, Z => b_new_21_port);
   U20 : XOR2_X1 port map( A => b(20), B => as, Z => b_new_20_port);
   U21 : XOR2_X1 port map( A => b(1), B => as, Z => b_new_1_port);
   U22 : XOR2_X1 port map( A => b(19), B => as, Z => b_new_19_port);
   U23 : XOR2_X1 port map( A => b(18), B => as, Z => b_new_18_port);
   U24 : XOR2_X1 port map( A => b(17), B => as, Z => b_new_17_port);
   U25 : XOR2_X1 port map( A => b(16), B => as, Z => b_new_16_port);
   U26 : XOR2_X1 port map( A => b(15), B => as, Z => b_new_15_port);
   U27 : XOR2_X1 port map( A => b(14), B => as, Z => b_new_14_port);
   U28 : XOR2_X1 port map( A => b(13), B => as, Z => b_new_13_port);
   U29 : XOR2_X1 port map( A => b(12), B => as, Z => b_new_12_port);
   U30 : XOR2_X1 port map( A => b(11), B => as, Z => b_new_11_port);
   U31 : XOR2_X1 port map( A => b(10), B => as, Z => b_new_10_port);
   U32 : XOR2_X1 port map( A => b(0), B => as, Z => b_new_0_port);

end SYN_add_sub_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity BoothMul_DATA_SIZE16_STAGE10 is

   port( rst, clk, en, lock, sign : in std_logic;  a, b : in std_logic_vector 
         (15 downto 0);  o : out std_logic_vector (31 downto 0));

end BoothMul_DATA_SIZE16_STAGE10;

architecture SYN_booth_mul_arch of BoothMul_DATA_SIZE16_STAGE10 is

   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X4
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BoothMul_DATA_SIZE16_STAGE10_DW01_inc_0
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component Adder_DATA_SIZE32_5
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;
   
   component Reg_DATA_SIZE32_1
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 
            0);  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component AddSub_DATA_SIZE32_1
      port( as : in std_logic;  a, b : in std_logic_vector (31 downto 0);  re :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;
   
   component Mux_DATA_SIZE32_1
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0)
            ;  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component BoothEncoder
      port( din : in std_logic_vector (2 downto 0);  sel : out std_logic_vector
            (2 downto 0));
   end component;
   
   component Adder_DATA_SIZE16
      port( cin : in std_logic;  a, b : in std_logic_vector (15 downto 0);  s :
            out std_logic_vector (15 downto 0);  cout : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic0_port, e_a_31_port, e_a_30_port, e_a_29_port, e_a_28_port, 
      e_a_27_port, e_a_26_port, e_a_25_port, e_a_24_port, e_a_23_port, 
      e_a_22_port, e_a_21_port, e_a_20_port, e_a_19_port, e_a_18_port, 
      e_a_17_port, e_a_16_port, e_a_15_port, e_a_14_port, e_a_13_port, 
      e_a_12_port, e_a_11_port, e_a_10_port, e_a_9_port, e_a_8_port, e_a_7_port
      , e_a_6_port, e_a_5_port, e_a_4_port, e_a_3_port, e_a_2_port, e_a_1_port,
      e_a_0_port, e_b_16_port, e_b_15_port, e_b_14_port, e_b_13_port, 
      e_b_12_port, e_b_11_port, e_b_10_port, e_b_9_port, e_b_8_port, e_b_7_port
      , e_b_6_port, e_b_5_port, e_b_4_port, e_b_3_port, e_b_2_port, e_b_1_port,
      e_b_0_port, adj_final_mod_31_port, adj_final_mod_30_port, 
      adj_final_mod_29_port, adj_final_mod_28_port, adj_final_mod_27_port, 
      adj_final_mod_26_port, adj_final_mod_25_port, adj_final_mod_24_port, 
      adj_final_mod_23_port, adj_final_mod_22_port, adj_final_mod_21_port, 
      adj_final_mod_20_port, adj_final_mod_19_port, adj_final_mod_18_port, 
      adj_final_mod_17_port, adj_final_mod_16_port, adj_final_mod_15_port, 
      adj_final_mod_14_port, adj_final_mod_13_port, adj_final_mod_12_port, 
      adj_final_mod_11_port, adj_final_mod_10_port, adj_final_mod_9_port, 
      adj_final_mod_8_port, adj_final_mod_7_port, adj_final_mod_6_port, 
      adj_final_mod_5_port, adj_final_mod_4_port, adj_final_mod_3_port, 
      adj_final_mod_2_port, adj_final_mod_1_port, adj_final_mod_0_port, N9, N10
      , N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, 
      N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39
      , N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, 
      N54, N55, N56, N57, adj_sum_15_port, adj_sum_14_port, adj_sum_13_port, 
      adj_sum_12_port, adj_sum_11_port, adj_sum_10_port, adj_sum_9_port, 
      adj_sum_8_port, adj_sum_7_port, adj_sum_6_port, adj_sum_5_port, 
      adj_sum_4_port, adj_sum_3_port, adj_sum_2_port, adj_sum_1_port, 
      adj_sum_0_port, adj_cout, sel_2_port, sel_1_port, sel_0_port, 
      mux_out_31_port, mux_out_30_port, mux_out_29_port, mux_out_28_port, 
      mux_out_27_port, mux_out_26_port, mux_out_25_port, mux_out_24_port, 
      mux_out_23_port, mux_out_22_port, mux_out_21_port, mux_out_20_port, 
      mux_out_19_port, mux_out_18_port, mux_out_17_port, mux_out_16_port, 
      mux_out_15_port, mux_out_14_port, mux_out_13_port, mux_out_12_port, 
      mux_out_11_port, mux_out_10_port, mux_out_9_port, mux_out_8_port, 
      mux_out_7_port, mux_out_6_port, mux_out_5_port, mux_out_4_port, 
      mux_out_3_port, mux_out_2_port, mux_out_1_port, mux_out_0_port, 
      zero_out_31_port, zero_out_30_port, zero_out_29_port, zero_out_28_port, 
      zero_out_27_port, zero_out_26_port, zero_out_25_port, zero_out_24_port, 
      zero_out_23_port, zero_out_22_port, zero_out_21_port, zero_out_20_port, 
      zero_out_19_port, zero_out_18_port, zero_out_17_port, zero_out_16_port, 
      zero_out_15_port, zero_out_14_port, zero_out_13_port, zero_out_12_port, 
      zero_out_11_port, zero_out_10_port, zero_out_9_port, zero_out_8_port, 
      zero_out_7_port, zero_out_6_port, zero_out_5_port, zero_out_4_port, 
      zero_out_3_port, zero_out_2_port, zero_out_1_port, zero_out_0_port, 
      add_out_reg_31_port, add_out_reg_30_port, add_out_reg_29_port, 
      add_out_reg_28_port, add_out_reg_27_port, add_out_reg_26_port, 
      add_out_reg_25_port, add_out_reg_24_port, add_out_reg_23_port, 
      add_out_reg_22_port, add_out_reg_21_port, add_out_reg_20_port, 
      add_out_reg_19_port, add_out_reg_18_port, add_out_reg_17_port, 
      add_out_reg_16_port, add_out_reg_15_port, add_out_reg_14_port, 
      add_out_reg_13_port, add_out_reg_12_port, add_out_reg_11_port, 
      add_out_reg_10_port, add_out_reg_9_port, add_out_reg_8_port, 
      add_out_reg_7_port, add_out_reg_6_port, add_out_reg_5_port, 
      add_out_reg_4_port, add_out_reg_3_port, add_out_reg_2_port, 
      add_out_reg_1_port, add_out_reg_0_port, add_out_31_port, add_out_30_port,
      add_out_29_port, add_out_28_port, add_out_27_port, add_out_26_port, 
      add_out_25_port, add_out_24_port, add_out_23_port, add_out_22_port, 
      add_out_21_port, add_out_20_port, add_out_19_port, add_out_18_port, 
      add_out_17_port, add_out_16_port, add_out_15_port, add_out_14_port, 
      add_out_13_port, add_out_12_port, add_out_11_port, add_out_10_port, 
      add_out_9_port, add_out_8_port, add_out_7_port, add_out_6_port, 
      add_out_5_port, add_out_4_port, add_out_3_port, add_out_2_port, 
      add_out_1_port, add_out_0_port, reg_rst, en_o, n_state_31_port, 
      n_state_30_port, n_state_29_port, n_state_28_port, n_state_27_port, 
      n_state_26_port, n_state_25_port, n_state_24_port, n_state_23_port, 
      n_state_22_port, n_state_21_port, n_state_20_port, n_state_19_port, 
      n_state_18_port, n_state_17_port, n_state_16_port, n_state_15_port, 
      n_state_14_port, n_state_13_port, n_state_12_port, n_state_11_port, 
      n_state_10_port, n_state_9_port, n_state_8_port, n_state_7_port, 
      n_state_6_port, n_state_5_port, n_state_4_port, n_state_3_port, 
      n_state_2_port, n_state_1_port, n_state_0_port, c_state_31_port, 
      c_state_30_port, c_state_29_port, c_state_28_port, c_state_27_port, 
      c_state_26_port, c_state_25_port, c_state_24_port, c_state_23_port, 
      c_state_22_port, c_state_21_port, c_state_20_port, c_state_19_port, 
      c_state_18_port, c_state_17_port, c_state_16_port, c_state_15_port, 
      c_state_14_port, c_state_13_port, c_state_12_port, c_state_11_port, 
      c_state_10_port, c_state_9_port, c_state_8_port, c_state_7_port, 
      c_state_6_port, c_state_5_port, c_state_4_port, c_state_3_port, 
      c_state_2_port, c_state_1_port, c_state_0_port, N70, N71, N72, N73, N74, 
      N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89
      , N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101, net4347, 
      net4348, n12_port, n13_port, n22_port, n23_port, n24_port, n28_port, 
      n29_port, n30_port, n31_port, n58, n65, n66, n67, n68, n69, n70_port, 
      n71_port, n72_port, n79_port, n80_port, n81_port, n82_port, n83_port, 
      n84_port, n85_port, n86_port, n87_port, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205, n206, n207, n208, n209, n210, n211, n1, n2, n3, n4, n5, n6, n7, n8,
      n9_port, n10_port, n11_port, n14_port, n15_port, n16_port, n17_port, 
      n18_port, n19_port, n20_port, n21_port, n25_port, n26_port, n27_port, 
      n32_port, n33_port, n34_port, n35_port, n36_port, n37_port, n38_port, 
      n39_port, n40_port, n41_port, n42_port, n43_port, n44_port, n45_port, 
      n46_port, n47_port, n48_port, n49_port, n50_port, n51_port, n52_port, 
      n53_port, n54_port, n55_port, n56_port, n57_port, n59, n60, n61, n62, n63
      , net108691, net108692, net108693, net108694, net108695, net108696, 
      net108697, net108698, net108699, net108700, net108701, net108702, 
      net108703, net108704, net108705, net108706, net108707, net108708, 
      net108709, net108710, net108711, net108712, net108713, net108714, 
      net108715, net108716, net108717, net108718, net108719, net108720, 
      net108721, net108722, net108723, net108724, net108725, net108726, 
      net108727, net108728, net108729, net108730, net108731, net108732, 
      net108733, net108734, net108735, net108736, net108737, net108738, 
      net108739, net108740, net108741, net108742, net108743, net108744 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   c_state_reg_0_inst : DFFR_X1 port map( D => n_state_0_port, CK => clk, RN =>
                           rst, Q => c_state_0_port, QN => n211);
   c_state_reg_10_inst : DFFR_X1 port map( D => n_state_10_port, CK => clk, RN 
                           => rst, Q => c_state_10_port, QN => n12_port);
   c_state_reg_1_inst : DFFR_X1 port map( D => n_state_1_port, CK => clk, RN =>
                           rst, Q => c_state_1_port, QN => n13_port);
   c_state_reg_2_inst : DFFR_X1 port map( D => n_state_2_port, CK => clk, RN =>
                           rst, Q => c_state_2_port, QN => n55_port);
   c_state_reg_3_inst : DFFR_X1 port map( D => n_state_3_port, CK => clk, RN =>
                           rst, Q => c_state_3_port, QN => n54_port);
   c_state_reg_4_inst : DFFR_X1 port map( D => n_state_4_port, CK => clk, RN =>
                           rst, Q => c_state_4_port, QN => n57_port);
   c_state_reg_5_inst : DFFR_X1 port map( D => n_state_5_port, CK => clk, RN =>
                           rst, Q => c_state_5_port, QN => n59);
   c_state_reg_6_inst : DFFR_X1 port map( D => n_state_6_port, CK => clk, RN =>
                           rst, Q => c_state_6_port, QN => net108744);
   c_state_reg_7_inst : DFFR_X1 port map( D => n_state_7_port, CK => clk, RN =>
                           rst, Q => c_state_7_port, QN => net108743);
   c_state_reg_8_inst : DFFR_X1 port map( D => n_state_8_port, CK => clk, RN =>
                           rst, Q => c_state_8_port, QN => net108742);
   c_state_reg_9_inst : DFFR_X1 port map( D => n_state_9_port, CK => clk, RN =>
                           rst, Q => c_state_9_port, QN => n56_port);
   c_state_reg_11_inst : DFFR_X1 port map( D => n_state_11_port, CK => clk, RN 
                           => rst, Q => c_state_11_port, QN => n22_port);
   c_state_reg_12_inst : DFFR_X1 port map( D => n_state_12_port, CK => clk, RN 
                           => rst, Q => c_state_12_port, QN => n23_port);
   c_state_reg_13_inst : DFFR_X1 port map( D => n_state_13_port, CK => clk, RN 
                           => rst, Q => c_state_13_port, QN => n24_port);
   c_state_reg_14_inst : DFFR_X1 port map( D => n_state_14_port, CK => clk, RN 
                           => rst, Q => c_state_14_port, QN => net108741);
   c_state_reg_15_inst : DFFR_X1 port map( D => n_state_15_port, CK => clk, RN 
                           => rst, Q => c_state_15_port, QN => net108740);
   c_state_reg_16_inst : DFFR_X1 port map( D => n_state_16_port, CK => clk, RN 
                           => rst, Q => c_state_16_port, QN => net108739);
   c_state_reg_17_inst : DFFR_X1 port map( D => n_state_17_port, CK => clk, RN 
                           => rst, Q => c_state_17_port, QN => n28_port);
   c_state_reg_18_inst : DFFR_X1 port map( D => n_state_18_port, CK => clk, RN 
                           => rst, Q => c_state_18_port, QN => n29_port);
   c_state_reg_19_inst : DFFR_X1 port map( D => n_state_19_port, CK => clk, RN 
                           => rst, Q => c_state_19_port, QN => n30_port);
   c_state_reg_20_inst : DFFR_X1 port map( D => n_state_20_port, CK => clk, RN 
                           => rst, Q => c_state_20_port, QN => n31_port);
   c_state_reg_21_inst : DFFR_X1 port map( D => n_state_21_port, CK => clk, RN 
                           => rst, Q => c_state_21_port, QN => net108738);
   c_state_reg_22_inst : DFFR_X1 port map( D => n_state_22_port, CK => clk, RN 
                           => rst, Q => c_state_22_port, QN => net108737);
   c_state_reg_23_inst : DFFR_X1 port map( D => n_state_23_port, CK => clk, RN 
                           => rst, Q => c_state_23_port, QN => net108736);
   c_state_reg_24_inst : DFFR_X1 port map( D => n_state_24_port, CK => clk, RN 
                           => rst, Q => c_state_24_port, QN => n62);
   c_state_reg_25_inst : DFFR_X1 port map( D => n_state_25_port, CK => clk, RN 
                           => rst, Q => c_state_25_port, QN => n63);
   c_state_reg_26_inst : DFFR_X1 port map( D => n_state_26_port, CK => clk, RN 
                           => rst, Q => c_state_26_port, QN => net108735);
   c_state_reg_27_inst : DFFR_X1 port map( D => n_state_27_port, CK => clk, RN 
                           => rst, Q => c_state_27_port, QN => net108734);
   c_state_reg_28_inst : DFFR_X1 port map( D => n_state_28_port, CK => clk, RN 
                           => rst, Q => c_state_28_port, QN => n60);
   c_state_reg_29_inst : DFFR_X1 port map( D => n_state_29_port, CK => clk, RN 
                           => rst, Q => c_state_29_port, QN => n61);
   c_state_reg_30_inst : DFFR_X1 port map( D => n_state_30_port, CK => clk, RN 
                           => rst, Q => c_state_30_port, QN => net108733);
   c_state_reg_31_inst : DFFR_X1 port map( D => n_state_31_port, CK => clk, RN 
                           => rst, Q => c_state_31_port, QN => n53_port);
   adj_final_mod_reg_31_inst : DFF_X1 port map( D => n210, CK => clk, Q => 
                           adj_final_mod_31_port, QN => n189);
   adj_final_mod_reg_30_inst : DFF_X1 port map( D => n209, CK => clk, Q => 
                           adj_final_mod_30_port, QN => n188);
   adj_final_mod_reg_29_inst : DFF_X1 port map( D => n208, CK => clk, Q => 
                           adj_final_mod_29_port, QN => net108732);
   adj_final_mod_reg_28_inst : DFF_X1 port map( D => n207, CK => clk, Q => 
                           adj_final_mod_28_port, QN => net108731);
   adj_final_mod_reg_27_inst : DFF_X1 port map( D => n206, CK => clk, Q => 
                           adj_final_mod_27_port, QN => net108730);
   adj_final_mod_reg_26_inst : DFF_X1 port map( D => n205, CK => clk, Q => 
                           adj_final_mod_26_port, QN => net108729);
   adj_final_mod_reg_25_inst : DFF_X1 port map( D => n204, CK => clk, Q => 
                           adj_final_mod_25_port, QN => net108728);
   adj_final_mod_reg_24_inst : DFF_X1 port map( D => n203, CK => clk, Q => 
                           adj_final_mod_24_port, QN => net108727);
   adj_final_mod_reg_23_inst : DFF_X1 port map( D => n202, CK => clk, Q => 
                           adj_final_mod_23_port, QN => net108726);
   adj_final_mod_reg_22_inst : DFF_X1 port map( D => n201, CK => clk, Q => 
                           adj_final_mod_22_port, QN => net108725);
   adj_final_mod_reg_21_inst : DFF_X1 port map( D => n200, CK => clk, Q => 
                           adj_final_mod_21_port, QN => net108724);
   adj_final_mod_reg_20_inst : DFF_X1 port map( D => n199, CK => clk, Q => 
                           adj_final_mod_20_port, QN => net108723);
   adj_final_mod_reg_19_inst : DFF_X1 port map( D => n198, CK => clk, Q => 
                           adj_final_mod_19_port, QN => net108722);
   adj_final_mod_reg_18_inst : DFF_X1 port map( D => n197, CK => clk, Q => 
                           adj_final_mod_18_port, QN => net108721);
   adj_final_mod_reg_17_inst : DFF_X1 port map( D => n196, CK => clk, Q => 
                           adj_final_mod_17_port, QN => net108720);
   adj_final_mod_reg_16_inst : DFF_X1 port map( D => n195, CK => clk, Q => 
                           adj_final_mod_16_port, QN => net108719);
   adj_final_mod_reg_15_inst : DFF_X1 port map( D => n194, CK => clk, Q => 
                           adj_final_mod_15_port, QN => net108718);
   e_a_reg_0_inst : DFF_X1 port map( D => N9, CK => clk, Q => e_a_0_port, QN =>
                           net108717);
   e_b_reg_16_inst : DFF_X1 port map( D => N57, CK => clk, Q => e_b_16_port, QN
                           => net108716);
   e_b_reg_15_inst : DFF_X1 port map( D => N56, CK => clk, Q => e_b_15_port, QN
                           => net108715);
   e_b_reg_14_inst : DFF_X1 port map( D => N55, CK => clk, Q => e_b_14_port, QN
                           => net108714);
   e_b_reg_13_inst : DFF_X1 port map( D => N54, CK => clk, Q => e_b_13_port, QN
                           => net108713);
   e_b_reg_12_inst : DFF_X1 port map( D => N53, CK => clk, Q => e_b_12_port, QN
                           => net108712);
   e_b_reg_11_inst : DFF_X1 port map( D => N52, CK => clk, Q => e_b_11_port, QN
                           => net108711);
   e_b_reg_10_inst : DFF_X1 port map( D => N51, CK => clk, Q => e_b_10_port, QN
                           => net108710);
   e_b_reg_9_inst : DFF_X1 port map( D => N50, CK => clk, Q => e_b_9_port, QN 
                           => net108709);
   e_b_reg_8_inst : DFF_X1 port map( D => N49, CK => clk, Q => e_b_8_port, QN 
                           => net108708);
   e_b_reg_7_inst : DFF_X1 port map( D => N48, CK => clk, Q => e_b_7_port, QN 
                           => net108707);
   e_b_reg_6_inst : DFF_X1 port map( D => N47, CK => clk, Q => e_b_6_port, QN 
                           => net108706);
   e_b_reg_5_inst : DFF_X1 port map( D => N46, CK => clk, Q => e_b_5_port, QN 
                           => net108705);
   e_b_reg_4_inst : DFF_X1 port map( D => N45, CK => clk, Q => e_b_4_port, QN 
                           => net108704);
   e_b_reg_3_inst : DFF_X1 port map( D => N44, CK => clk, Q => e_b_3_port, QN 
                           => net108703);
   e_b_reg_2_inst : DFF_X1 port map( D => N43, CK => clk, Q => e_b_2_port, QN 
                           => n58);
   e_b_reg_0_inst : DFF_X1 port map( D => N41, CK => clk, Q => e_b_0_port, QN 
                           => n193);
   e_b_reg_1_inst : DFF_X1 port map( D => N42, CK => clk, Q => e_b_1_port, QN 
                           => n192);
   e_a_reg_2_inst : DFF_X1 port map( D => N11, CK => clk, Q => e_a_2_port, QN 
                           => net108702);
   e_a_reg_4_inst : DFF_X1 port map( D => N13, CK => clk, Q => e_a_4_port, QN 
                           => net108701);
   e_a_reg_6_inst : DFF_X1 port map( D => N15, CK => clk, Q => e_a_6_port, QN 
                           => net108700);
   e_a_reg_8_inst : DFF_X1 port map( D => N17, CK => clk, Q => e_a_8_port, QN 
                           => net108699);
   e_a_reg_10_inst : DFF_X1 port map( D => N19, CK => clk, Q => e_a_10_port, QN
                           => net108698);
   e_a_reg_12_inst : DFF_X1 port map( D => N21, CK => clk, Q => e_a_12_port, QN
                           => net108697);
   e_a_reg_14_inst : DFF_X1 port map( D => N23, CK => clk, Q => e_a_14_port, QN
                           => n65);
   e_a_reg_16_inst : DFF_X1 port map( D => N25, CK => clk, Q => e_a_16_port, QN
                           => n66);
   e_a_reg_18_inst : DFF_X1 port map( D => N27, CK => clk, Q => e_a_18_port, QN
                           => n67);
   e_a_reg_20_inst : DFF_X1 port map( D => N29, CK => clk, Q => e_a_20_port, QN
                           => n68);
   e_a_reg_22_inst : DFF_X1 port map( D => N31, CK => clk, Q => e_a_22_port, QN
                           => n69);
   e_a_reg_24_inst : DFF_X1 port map( D => N33, CK => clk, Q => e_a_24_port, QN
                           => n70_port);
   e_a_reg_26_inst : DFF_X1 port map( D => N35, CK => clk, Q => e_a_26_port, QN
                           => n71_port);
   e_a_reg_28_inst : DFF_X1 port map( D => N37, CK => clk, Q => e_a_28_port, QN
                           => n72_port);
   e_a_reg_30_inst : DFF_X1 port map( D => N39, CK => clk, Q => e_a_30_port, QN
                           => n191);
   e_a_reg_1_inst : DFF_X1 port map( D => N10, CK => clk, Q => e_a_1_port, QN 
                           => net108696);
   e_a_reg_3_inst : DFF_X1 port map( D => N12, CK => clk, Q => e_a_3_port, QN 
                           => net108695);
   e_a_reg_5_inst : DFF_X1 port map( D => N14, CK => clk, Q => e_a_5_port, QN 
                           => net108694);
   e_a_reg_7_inst : DFF_X1 port map( D => N16, CK => clk, Q => e_a_7_port, QN 
                           => net108693);
   e_a_reg_9_inst : DFF_X1 port map( D => N18, CK => clk, Q => e_a_9_port, QN 
                           => net108692);
   e_a_reg_11_inst : DFF_X1 port map( D => N20, CK => clk, Q => e_a_11_port, QN
                           => net108691);
   e_a_reg_13_inst : DFF_X1 port map( D => N22, CK => clk, Q => e_a_13_port, QN
                           => n79_port);
   e_a_reg_15_inst : DFF_X1 port map( D => N24, CK => clk, Q => e_a_15_port, QN
                           => n80_port);
   e_a_reg_17_inst : DFF_X1 port map( D => N26, CK => clk, Q => e_a_17_port, QN
                           => n81_port);
   e_a_reg_19_inst : DFF_X1 port map( D => N28, CK => clk, Q => e_a_19_port, QN
                           => n82_port);
   e_a_reg_21_inst : DFF_X1 port map( D => N30, CK => clk, Q => e_a_21_port, QN
                           => n83_port);
   e_a_reg_23_inst : DFF_X1 port map( D => N32, CK => clk, Q => e_a_23_port, QN
                           => n84_port);
   e_a_reg_25_inst : DFF_X1 port map( D => N34, CK => clk, Q => e_a_25_port, QN
                           => n85_port);
   e_a_reg_27_inst : DFF_X1 port map( D => N36, CK => clk, Q => e_a_27_port, QN
                           => n86_port);
   e_a_reg_29_inst : DFF_X1 port map( D => N38, CK => clk, Q => e_a_29_port, QN
                           => n87_port);
   e_a_reg_31_inst : DFF_X1 port map( D => N40, CK => clk, Q => e_a_31_port, QN
                           => n190);
   adj_final_mod_0_port <= '0';
   adj_final_mod_1_port <= '0';
   adj_final_mod_2_port <= '0';
   adj_final_mod_3_port <= '0';
   adj_final_mod_4_port <= '0';
   adj_final_mod_5_port <= '0';
   adj_final_mod_6_port <= '0';
   adj_final_mod_7_port <= '0';
   adj_final_mod_8_port <= '0';
   adj_final_mod_9_port <= '0';
   adj_final_mod_10_port <= '0';
   adj_final_mod_11_port <= '0';
   adj_final_mod_12_port <= '0';
   adj_final_mod_13_port <= '0';
   adj_final_mod_14_port <= '0';
   ADJUST0 : Adder_DATA_SIZE16 port map( cin => X_Logic0_port, a(15) => a(15), 
                           a(14) => a(14), a(13) => a(13), a(12) => a(12), 
                           a(11) => a(11), a(10) => a(10), a(9) => a(9), a(8) 
                           => a(8), a(7) => a(7), a(6) => a(6), a(5) => a(5), 
                           a(4) => a(4), a(3) => a(3), a(2) => a(2), a(1) => 
                           a(1), a(0) => a(0), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           s(15) => adj_sum_15_port, s(14) => adj_sum_14_port, 
                           s(13) => adj_sum_13_port, s(12) => adj_sum_12_port, 
                           s(11) => adj_sum_11_port, s(10) => adj_sum_10_port, 
                           s(9) => adj_sum_9_port, s(8) => adj_sum_8_port, s(7)
                           => adj_sum_7_port, s(6) => adj_sum_6_port, s(5) => 
                           adj_sum_5_port, s(4) => adj_sum_4_port, s(3) => 
                           adj_sum_3_port, s(2) => adj_sum_2_port, s(1) => 
                           adj_sum_1_port, s(0) => adj_sum_0_port, cout => 
                           adj_cout);
   BEC0 : BoothEncoder port map( din(2) => e_b_2_port, din(1) => e_b_1_port, 
                           din(0) => e_b_0_port, sel(2) => sel_2_port, sel(1) 
                           => sel_1_port, sel(0) => sel_0_port);
   MUX0 : Mux_DATA_SIZE32_1 port map( sel => sel_0_port, din0(31) => 
                           e_a_31_port, din0(30) => e_a_30_port, din0(29) => 
                           e_a_29_port, din0(28) => e_a_28_port, din0(27) => 
                           e_a_27_port, din0(26) => e_a_26_port, din0(25) => 
                           e_a_25_port, din0(24) => e_a_24_port, din0(23) => 
                           e_a_23_port, din0(22) => e_a_22_port, din0(21) => 
                           e_a_21_port, din0(20) => e_a_20_port, din0(19) => 
                           e_a_19_port, din0(18) => e_a_18_port, din0(17) => 
                           e_a_17_port, din0(16) => e_a_16_port, din0(15) => 
                           e_a_15_port, din0(14) => e_a_14_port, din0(13) => 
                           e_a_13_port, din0(12) => e_a_12_port, din0(11) => 
                           e_a_11_port, din0(10) => e_a_10_port, din0(9) => 
                           e_a_9_port, din0(8) => e_a_8_port, din0(7) => 
                           e_a_7_port, din0(6) => e_a_6_port, din0(5) => 
                           e_a_5_port, din0(4) => e_a_4_port, din0(3) => 
                           e_a_3_port, din0(2) => e_a_2_port, din0(1) => 
                           e_a_1_port, din0(0) => e_a_0_port, din1(31) => 
                           e_a_30_port, din1(30) => e_a_29_port, din1(29) => 
                           e_a_28_port, din1(28) => e_a_27_port, din1(27) => 
                           e_a_26_port, din1(26) => e_a_25_port, din1(25) => 
                           e_a_24_port, din1(24) => e_a_23_port, din1(23) => 
                           e_a_22_port, din1(22) => e_a_21_port, din1(21) => 
                           e_a_20_port, din1(20) => e_a_19_port, din1(19) => 
                           e_a_18_port, din1(18) => e_a_17_port, din1(17) => 
                           e_a_16_port, din1(16) => e_a_15_port, din1(15) => 
                           e_a_14_port, din1(14) => e_a_13_port, din1(13) => 
                           e_a_12_port, din1(12) => e_a_11_port, din1(11) => 
                           e_a_10_port, din1(10) => e_a_9_port, din1(9) => 
                           e_a_8_port, din1(8) => e_a_7_port, din1(7) => 
                           e_a_6_port, din1(6) => e_a_5_port, din1(5) => 
                           e_a_4_port, din1(4) => e_a_3_port, din1(3) => 
                           e_a_2_port, din1(2) => e_a_1_port, din1(1) => 
                           e_a_0_port, din1(0) => X_Logic0_port, dout(31) => 
                           mux_out_31_port, dout(30) => mux_out_30_port, 
                           dout(29) => mux_out_29_port, dout(28) => 
                           mux_out_28_port, dout(27) => mux_out_27_port, 
                           dout(26) => mux_out_26_port, dout(25) => 
                           mux_out_25_port, dout(24) => mux_out_24_port, 
                           dout(23) => mux_out_23_port, dout(22) => 
                           mux_out_22_port, dout(21) => mux_out_21_port, 
                           dout(20) => mux_out_20_port, dout(19) => 
                           mux_out_19_port, dout(18) => mux_out_18_port, 
                           dout(17) => mux_out_17_port, dout(16) => 
                           mux_out_16_port, dout(15) => mux_out_15_port, 
                           dout(14) => mux_out_14_port, dout(13) => 
                           mux_out_13_port, dout(12) => mux_out_12_port, 
                           dout(11) => mux_out_11_port, dout(10) => 
                           mux_out_10_port, dout(9) => mux_out_9_port, dout(8) 
                           => mux_out_8_port, dout(7) => mux_out_7_port, 
                           dout(6) => mux_out_6_port, dout(5) => mux_out_5_port
                           , dout(4) => mux_out_4_port, dout(3) => 
                           mux_out_3_port, dout(2) => mux_out_2_port, dout(1) 
                           => mux_out_1_port, dout(0) => mux_out_0_port);
   ADDSUBn : AddSub_DATA_SIZE32_1 port map( as => sel_1_port, a(31) => 
                           add_out_reg_31_port, a(30) => add_out_reg_30_port, 
                           a(29) => add_out_reg_29_port, a(28) => 
                           add_out_reg_28_port, a(27) => add_out_reg_27_port, 
                           a(26) => add_out_reg_26_port, a(25) => 
                           add_out_reg_25_port, a(24) => add_out_reg_24_port, 
                           a(23) => add_out_reg_23_port, a(22) => 
                           add_out_reg_22_port, a(21) => add_out_reg_21_port, 
                           a(20) => add_out_reg_20_port, a(19) => 
                           add_out_reg_19_port, a(18) => add_out_reg_18_port, 
                           a(17) => add_out_reg_17_port, a(16) => 
                           add_out_reg_16_port, a(15) => add_out_reg_15_port, 
                           a(14) => add_out_reg_14_port, a(13) => 
                           add_out_reg_13_port, a(12) => add_out_reg_12_port, 
                           a(11) => add_out_reg_11_port, a(10) => 
                           add_out_reg_10_port, a(9) => add_out_reg_9_port, 
                           a(8) => add_out_reg_8_port, a(7) => 
                           add_out_reg_7_port, a(6) => add_out_reg_6_port, a(5)
                           => add_out_reg_5_port, a(4) => add_out_reg_4_port, 
                           a(3) => add_out_reg_3_port, a(2) => 
                           add_out_reg_2_port, a(1) => add_out_reg_1_port, a(0)
                           => add_out_reg_0_port, b(31) => zero_out_31_port, 
                           b(30) => zero_out_30_port, b(29) => zero_out_29_port
                           , b(28) => zero_out_28_port, b(27) => 
                           zero_out_27_port, b(26) => zero_out_26_port, b(25) 
                           => zero_out_25_port, b(24) => zero_out_24_port, 
                           b(23) => zero_out_23_port, b(22) => zero_out_22_port
                           , b(21) => zero_out_21_port, b(20) => 
                           zero_out_20_port, b(19) => zero_out_19_port, b(18) 
                           => zero_out_18_port, b(17) => zero_out_17_port, 
                           b(16) => zero_out_16_port, b(15) => zero_out_15_port
                           , b(14) => zero_out_14_port, b(13) => 
                           zero_out_13_port, b(12) => zero_out_12_port, b(11) 
                           => zero_out_11_port, b(10) => zero_out_10_port, b(9)
                           => zero_out_9_port, b(8) => zero_out_8_port, b(7) =>
                           zero_out_7_port, b(6) => zero_out_6_port, b(5) => 
                           zero_out_5_port, b(4) => zero_out_4_port, b(3) => 
                           zero_out_3_port, b(2) => zero_out_2_port, b(1) => 
                           zero_out_1_port, b(0) => zero_out_0_port, re(31) => 
                           add_out_31_port, re(30) => add_out_30_port, re(29) 
                           => add_out_29_port, re(28) => add_out_28_port, 
                           re(27) => add_out_27_port, re(26) => add_out_26_port
                           , re(25) => add_out_25_port, re(24) => 
                           add_out_24_port, re(23) => add_out_23_port, re(22) 
                           => add_out_22_port, re(21) => add_out_21_port, 
                           re(20) => add_out_20_port, re(19) => add_out_19_port
                           , re(18) => add_out_18_port, re(17) => 
                           add_out_17_port, re(16) => add_out_16_port, re(15) 
                           => add_out_15_port, re(14) => add_out_14_port, 
                           re(13) => add_out_13_port, re(12) => add_out_12_port
                           , re(11) => add_out_11_port, re(10) => 
                           add_out_10_port, re(9) => add_out_9_port, re(8) => 
                           add_out_8_port, re(7) => add_out_7_port, re(6) => 
                           add_out_6_port, re(5) => add_out_5_port, re(4) => 
                           add_out_4_port, re(3) => add_out_3_port, re(2) => 
                           add_out_2_port, re(1) => add_out_1_port, re(0) => 
                           add_out_0_port, cout => net4348);
   REG0 : Reg_DATA_SIZE32_1 port map( rst => reg_rst, en => en_o, clk => clk, 
                           din(31) => add_out_31_port, din(30) => 
                           add_out_30_port, din(29) => add_out_29_port, din(28)
                           => add_out_28_port, din(27) => add_out_27_port, 
                           din(26) => add_out_26_port, din(25) => 
                           add_out_25_port, din(24) => add_out_24_port, din(23)
                           => add_out_23_port, din(22) => add_out_22_port, 
                           din(21) => add_out_21_port, din(20) => 
                           add_out_20_port, din(19) => add_out_19_port, din(18)
                           => add_out_18_port, din(17) => add_out_17_port, 
                           din(16) => add_out_16_port, din(15) => 
                           add_out_15_port, din(14) => add_out_14_port, din(13)
                           => add_out_13_port, din(12) => add_out_12_port, 
                           din(11) => add_out_11_port, din(10) => 
                           add_out_10_port, din(9) => add_out_9_port, din(8) =>
                           add_out_8_port, din(7) => add_out_7_port, din(6) => 
                           add_out_6_port, din(5) => add_out_5_port, din(4) => 
                           add_out_4_port, din(3) => add_out_3_port, din(2) => 
                           add_out_2_port, din(1) => add_out_1_port, din(0) => 
                           add_out_0_port, dout(31) => add_out_reg_31_port, 
                           dout(30) => add_out_reg_30_port, dout(29) => 
                           add_out_reg_29_port, dout(28) => add_out_reg_28_port
                           , dout(27) => add_out_reg_27_port, dout(26) => 
                           add_out_reg_26_port, dout(25) => add_out_reg_25_port
                           , dout(24) => add_out_reg_24_port, dout(23) => 
                           add_out_reg_23_port, dout(22) => add_out_reg_22_port
                           , dout(21) => add_out_reg_21_port, dout(20) => 
                           add_out_reg_20_port, dout(19) => add_out_reg_19_port
                           , dout(18) => add_out_reg_18_port, dout(17) => 
                           add_out_reg_17_port, dout(16) => add_out_reg_16_port
                           , dout(15) => add_out_reg_15_port, dout(14) => 
                           add_out_reg_14_port, dout(13) => add_out_reg_13_port
                           , dout(12) => add_out_reg_12_port, dout(11) => 
                           add_out_reg_11_port, dout(10) => add_out_reg_10_port
                           , dout(9) => add_out_reg_9_port, dout(8) => 
                           add_out_reg_8_port, dout(7) => add_out_reg_7_port, 
                           dout(6) => add_out_reg_6_port, dout(5) => 
                           add_out_reg_5_port, dout(4) => add_out_reg_4_port, 
                           dout(3) => add_out_reg_3_port, dout(2) => 
                           add_out_reg_2_port, dout(1) => add_out_reg_1_port, 
                           dout(0) => add_out_reg_0_port);
   ADJUST1 : Adder_DATA_SIZE32_5 port map( cin => X_Logic0_port, a(31) => 
                           add_out_reg_31_port, a(30) => add_out_reg_30_port, 
                           a(29) => add_out_reg_29_port, a(28) => 
                           add_out_reg_28_port, a(27) => add_out_reg_27_port, 
                           a(26) => add_out_reg_26_port, a(25) => 
                           add_out_reg_25_port, a(24) => add_out_reg_24_port, 
                           a(23) => add_out_reg_23_port, a(22) => 
                           add_out_reg_22_port, a(21) => add_out_reg_21_port, 
                           a(20) => add_out_reg_20_port, a(19) => 
                           add_out_reg_19_port, a(18) => add_out_reg_18_port, 
                           a(17) => add_out_reg_17_port, a(16) => 
                           add_out_reg_16_port, a(15) => add_out_reg_15_port, 
                           a(14) => add_out_reg_14_port, a(13) => 
                           add_out_reg_13_port, a(12) => add_out_reg_12_port, 
                           a(11) => add_out_reg_11_port, a(10) => 
                           add_out_reg_10_port, a(9) => add_out_reg_9_port, 
                           a(8) => add_out_reg_8_port, a(7) => 
                           add_out_reg_7_port, a(6) => add_out_reg_6_port, a(5)
                           => add_out_reg_5_port, a(4) => add_out_reg_4_port, 
                           a(3) => add_out_reg_3_port, a(2) => 
                           add_out_reg_2_port, a(1) => add_out_reg_1_port, a(0)
                           => add_out_reg_0_port, b(31) => 
                           adj_final_mod_31_port, b(30) => 
                           adj_final_mod_30_port, b(29) => 
                           adj_final_mod_29_port, b(28) => 
                           adj_final_mod_28_port, b(27) => 
                           adj_final_mod_27_port, b(26) => 
                           adj_final_mod_26_port, b(25) => 
                           adj_final_mod_25_port, b(24) => 
                           adj_final_mod_24_port, b(23) => 
                           adj_final_mod_23_port, b(22) => 
                           adj_final_mod_22_port, b(21) => 
                           adj_final_mod_21_port, b(20) => 
                           adj_final_mod_20_port, b(19) => 
                           adj_final_mod_19_port, b(18) => 
                           adj_final_mod_18_port, b(17) => 
                           adj_final_mod_17_port, b(16) => 
                           adj_final_mod_16_port, b(15) => 
                           adj_final_mod_15_port, b(14) => 
                           adj_final_mod_14_port, b(13) => 
                           adj_final_mod_13_port, b(12) => 
                           adj_final_mod_12_port, b(11) => 
                           adj_final_mod_11_port, b(10) => 
                           adj_final_mod_10_port, b(9) => adj_final_mod_9_port,
                           b(8) => adj_final_mod_8_port, b(7) => 
                           adj_final_mod_7_port, b(6) => adj_final_mod_6_port, 
                           b(5) => adj_final_mod_5_port, b(4) => 
                           adj_final_mod_4_port, b(3) => adj_final_mod_3_port, 
                           b(2) => adj_final_mod_2_port, b(1) => 
                           adj_final_mod_1_port, b(0) => adj_final_mod_0_port, 
                           s(31) => o(31), s(30) => o(30), s(29) => o(29), 
                           s(28) => o(28), s(27) => o(27), s(26) => o(26), 
                           s(25) => o(25), s(24) => o(24), s(23) => o(23), 
                           s(22) => o(22), s(21) => o(21), s(20) => o(20), 
                           s(19) => o(19), s(18) => o(18), s(17) => o(17), 
                           s(16) => o(16), s(15) => o(15), s(14) => o(14), 
                           s(13) => o(13), s(12) => o(12), s(11) => o(11), 
                           s(10) => o(10), s(9) => o(9), s(8) => o(8), s(7) => 
                           o(7), s(6) => o(6), s(5) => o(5), s(4) => o(4), s(3)
                           => o(3), s(2) => o(2), s(1) => o(1), s(0) => o(0), 
                           cout => net4347);
   add_189 : BoothMul_DATA_SIZE16_STAGE10_DW01_inc_0 port map( A(31) => 
                           c_state_31_port, A(30) => c_state_30_port, A(29) => 
                           c_state_29_port, A(28) => c_state_28_port, A(27) => 
                           c_state_27_port, A(26) => c_state_26_port, A(25) => 
                           c_state_25_port, A(24) => c_state_24_port, A(23) => 
                           c_state_23_port, A(22) => c_state_22_port, A(21) => 
                           c_state_21_port, A(20) => c_state_20_port, A(19) => 
                           c_state_19_port, A(18) => c_state_18_port, A(17) => 
                           c_state_17_port, A(16) => c_state_16_port, A(15) => 
                           c_state_15_port, A(14) => c_state_14_port, A(13) => 
                           c_state_13_port, A(12) => c_state_12_port, A(11) => 
                           c_state_11_port, A(10) => c_state_10_port, A(9) => 
                           c_state_9_port, A(8) => c_state_8_port, A(7) => 
                           c_state_7_port, A(6) => c_state_6_port, A(5) => 
                           c_state_5_port, A(4) => c_state_4_port, A(3) => 
                           c_state_3_port, A(2) => c_state_2_port, A(1) => 
                           c_state_1_port, A(0) => c_state_0_port, SUM(31) => 
                           N101, SUM(30) => N100, SUM(29) => N99, SUM(28) => 
                           N98, SUM(27) => N97, SUM(26) => N96, SUM(25) => N95,
                           SUM(24) => N94, SUM(23) => N93, SUM(22) => N92, 
                           SUM(21) => N91, SUM(20) => N90, SUM(19) => N89, 
                           SUM(18) => N88, SUM(17) => N87, SUM(16) => N86, 
                           SUM(15) => N85, SUM(14) => N84, SUM(13) => N83, 
                           SUM(12) => N82, SUM(11) => N81, SUM(10) => N80, 
                           SUM(9) => N79, SUM(8) => N78, SUM(7) => N77, SUM(6) 
                           => N76, SUM(5) => N75, SUM(4) => N74, SUM(3) => N73,
                           SUM(2) => N72, SUM(1) => N71, SUM(0) => N70);
   U3 : AND2_X2 port map( A1 => rst, A2 => en_o, ZN => reg_rst);
   U4 : INV_X2 port map( A => n38_port, ZN => en_o);
   U5 : AOI21_X4 port map( B1 => en, B2 => lock, A => n6, ZN => n1);
   U6 : NOR2_X2 port map( A1 => n16_port, A2 => sign, ZN => n14_port);
   U7 : NAND2_X2 port map( A1 => en, A2 => n38_port, ZN => n16_port);
   U8 : AND2_X1 port map( A1 => sel_2_port, A2 => mux_out_9_port, ZN => 
                           zero_out_9_port);
   U9 : AND2_X1 port map( A1 => mux_out_8_port, A2 => sel_2_port, ZN => 
                           zero_out_8_port);
   U10 : AND2_X1 port map( A1 => mux_out_7_port, A2 => sel_2_port, ZN => 
                           zero_out_7_port);
   U11 : AND2_X1 port map( A1 => mux_out_6_port, A2 => sel_2_port, ZN => 
                           zero_out_6_port);
   U12 : AND2_X1 port map( A1 => mux_out_5_port, A2 => sel_2_port, ZN => 
                           zero_out_5_port);
   U13 : AND2_X1 port map( A1 => mux_out_4_port, A2 => sel_2_port, ZN => 
                           zero_out_4_port);
   U14 : AND2_X1 port map( A1 => mux_out_3_port, A2 => sel_2_port, ZN => 
                           zero_out_3_port);
   U15 : AND2_X1 port map( A1 => mux_out_31_port, A2 => sel_2_port, ZN => 
                           zero_out_31_port);
   U16 : AND2_X1 port map( A1 => mux_out_30_port, A2 => sel_2_port, ZN => 
                           zero_out_30_port);
   U17 : AND2_X1 port map( A1 => mux_out_2_port, A2 => sel_2_port, ZN => 
                           zero_out_2_port);
   U18 : AND2_X1 port map( A1 => mux_out_29_port, A2 => sel_2_port, ZN => 
                           zero_out_29_port);
   U19 : AND2_X1 port map( A1 => mux_out_28_port, A2 => sel_2_port, ZN => 
                           zero_out_28_port);
   U20 : AND2_X1 port map( A1 => mux_out_27_port, A2 => sel_2_port, ZN => 
                           zero_out_27_port);
   U21 : AND2_X1 port map( A1 => mux_out_26_port, A2 => sel_2_port, ZN => 
                           zero_out_26_port);
   U22 : AND2_X1 port map( A1 => mux_out_25_port, A2 => sel_2_port, ZN => 
                           zero_out_25_port);
   U23 : AND2_X1 port map( A1 => mux_out_24_port, A2 => sel_2_port, ZN => 
                           zero_out_24_port);
   U24 : AND2_X1 port map( A1 => mux_out_23_port, A2 => sel_2_port, ZN => 
                           zero_out_23_port);
   U25 : AND2_X1 port map( A1 => mux_out_22_port, A2 => sel_2_port, ZN => 
                           zero_out_22_port);
   U26 : AND2_X1 port map( A1 => mux_out_21_port, A2 => sel_2_port, ZN => 
                           zero_out_21_port);
   U27 : AND2_X1 port map( A1 => mux_out_20_port, A2 => sel_2_port, ZN => 
                           zero_out_20_port);
   U28 : AND2_X1 port map( A1 => mux_out_1_port, A2 => sel_2_port, ZN => 
                           zero_out_1_port);
   U29 : AND2_X1 port map( A1 => mux_out_19_port, A2 => sel_2_port, ZN => 
                           zero_out_19_port);
   U30 : AND2_X1 port map( A1 => mux_out_18_port, A2 => sel_2_port, ZN => 
                           zero_out_18_port);
   U31 : AND2_X1 port map( A1 => mux_out_17_port, A2 => sel_2_port, ZN => 
                           zero_out_17_port);
   U32 : AND2_X1 port map( A1 => mux_out_16_port, A2 => sel_2_port, ZN => 
                           zero_out_16_port);
   U33 : AND2_X1 port map( A1 => mux_out_15_port, A2 => sel_2_port, ZN => 
                           zero_out_15_port);
   U34 : AND2_X1 port map( A1 => mux_out_14_port, A2 => sel_2_port, ZN => 
                           zero_out_14_port);
   U35 : AND2_X1 port map( A1 => mux_out_13_port, A2 => sel_2_port, ZN => 
                           zero_out_13_port);
   U36 : AND2_X1 port map( A1 => mux_out_12_port, A2 => sel_2_port, ZN => 
                           zero_out_12_port);
   U37 : AND2_X1 port map( A1 => mux_out_11_port, A2 => sel_2_port, ZN => 
                           zero_out_11_port);
   U38 : AND2_X1 port map( A1 => mux_out_10_port, A2 => sel_2_port, ZN => 
                           zero_out_10_port);
   U39 : AND2_X1 port map( A1 => mux_out_0_port, A2 => sel_2_port, ZN => 
                           zero_out_0_port);
   U40 : AND2_X1 port map( A1 => N79, A2 => n1, ZN => n_state_9_port);
   U41 : AND2_X1 port map( A1 => N78, A2 => n1, ZN => n_state_8_port);
   U42 : AND2_X1 port map( A1 => N77, A2 => n1, ZN => n_state_7_port);
   U43 : AND2_X1 port map( A1 => N76, A2 => n1, ZN => n_state_6_port);
   U44 : AND2_X1 port map( A1 => N75, A2 => n1, ZN => n_state_5_port);
   U45 : AND2_X1 port map( A1 => N74, A2 => n1, ZN => n_state_4_port);
   U46 : AND2_X1 port map( A1 => N73, A2 => n1, ZN => n_state_3_port);
   U47 : AND2_X1 port map( A1 => N101, A2 => n1, ZN => n_state_31_port);
   U48 : AND2_X1 port map( A1 => N100, A2 => n1, ZN => n_state_30_port);
   U49 : AND2_X1 port map( A1 => N72, A2 => n1, ZN => n_state_2_port);
   U50 : AND2_X1 port map( A1 => N99, A2 => n1, ZN => n_state_29_port);
   U51 : AND2_X1 port map( A1 => N98, A2 => n1, ZN => n_state_28_port);
   U52 : AND2_X1 port map( A1 => N97, A2 => n1, ZN => n_state_27_port);
   U53 : AND2_X1 port map( A1 => N96, A2 => n1, ZN => n_state_26_port);
   U54 : AND2_X1 port map( A1 => N95, A2 => n1, ZN => n_state_25_port);
   U55 : AND2_X1 port map( A1 => N94, A2 => n1, ZN => n_state_24_port);
   U56 : AND2_X1 port map( A1 => N93, A2 => n1, ZN => n_state_23_port);
   U57 : AND2_X1 port map( A1 => N92, A2 => n1, ZN => n_state_22_port);
   U58 : AND2_X1 port map( A1 => N91, A2 => n1, ZN => n_state_21_port);
   U59 : AND2_X1 port map( A1 => N90, A2 => n1, ZN => n_state_20_port);
   U60 : AND2_X1 port map( A1 => N71, A2 => n1, ZN => n_state_1_port);
   U61 : AND2_X1 port map( A1 => N89, A2 => n1, ZN => n_state_19_port);
   U62 : AND2_X1 port map( A1 => N88, A2 => n1, ZN => n_state_18_port);
   U63 : AND2_X1 port map( A1 => N87, A2 => n1, ZN => n_state_17_port);
   U64 : AND2_X1 port map( A1 => N86, A2 => n1, ZN => n_state_16_port);
   U65 : AND2_X1 port map( A1 => N85, A2 => n1, ZN => n_state_15_port);
   U66 : AND2_X1 port map( A1 => N84, A2 => n1, ZN => n_state_14_port);
   U67 : AND2_X1 port map( A1 => N83, A2 => n1, ZN => n_state_13_port);
   U68 : AND2_X1 port map( A1 => N82, A2 => n1, ZN => n_state_12_port);
   U69 : AND2_X1 port map( A1 => N81, A2 => n1, ZN => n_state_11_port);
   U70 : AND2_X1 port map( A1 => N80, A2 => n1, ZN => n_state_10_port);
   U71 : INV_X1 port map( A => n2, ZN => n_state_0_port);
   U72 : AOI21_X1 port map( B1 => n1, B2 => N70, A => n3, ZN => n2);
   U73 : AND4_X1 port map( A1 => en, A2 => n53_port, A3 => n4, A4 => n211, ZN 
                           => n3);
   U74 : NOR2_X1 port map( A1 => lock, A2 => n5, ZN => n4);
   U75 : AOI21_X1 port map( B1 => n7, B2 => n8, A => c_state_31_port, ZN => n6)
                           ;
   U76 : MUX2_X1 port map( A => n5, B => n54_port, S => c_state_0_port, Z => n8
                           );
   U77 : OAI22_X1 port map( A1 => n189, A2 => n9_port, B1 => n10_port, B2 => 
                           n11_port, ZN => n210);
   U78 : XOR2_X1 port map( A => adj_sum_15_port, B => adj_cout, Z => n11_port);
   U79 : OAI22_X1 port map( A1 => n188, A2 => n9_port, B1 => adj_sum_15_port, 
                           B2 => n10_port, ZN => n209);
   U80 : INV_X1 port map( A => n14_port, ZN => n10_port);
   U81 : INV_X1 port map( A => n15_port, ZN => n208);
   U82 : AOI22_X1 port map( A1 => adj_sum_14_port, A2 => n14_port, B1 => 
                           n16_port, B2 => adj_final_mod_29_port, ZN => 
                           n15_port);
   U83 : INV_X1 port map( A => n17_port, ZN => n207);
   U84 : AOI22_X1 port map( A1 => adj_sum_13_port, A2 => n14_port, B1 => 
                           n16_port, B2 => adj_final_mod_28_port, ZN => 
                           n17_port);
   U85 : INV_X1 port map( A => n18_port, ZN => n206);
   U86 : AOI22_X1 port map( A1 => adj_sum_12_port, A2 => n14_port, B1 => 
                           n16_port, B2 => adj_final_mod_27_port, ZN => 
                           n18_port);
   U87 : INV_X1 port map( A => n19_port, ZN => n205);
   U88 : AOI22_X1 port map( A1 => adj_sum_11_port, A2 => n14_port, B1 => 
                           n16_port, B2 => adj_final_mod_26_port, ZN => 
                           n19_port);
   U89 : INV_X1 port map( A => n20_port, ZN => n204);
   U90 : AOI22_X1 port map( A1 => adj_sum_10_port, A2 => n14_port, B1 => 
                           n16_port, B2 => adj_final_mod_25_port, ZN => 
                           n20_port);
   U91 : INV_X1 port map( A => n21_port, ZN => n203);
   U92 : AOI22_X1 port map( A1 => adj_sum_9_port, A2 => n14_port, B1 => 
                           n16_port, B2 => adj_final_mod_24_port, ZN => 
                           n21_port);
   U93 : INV_X1 port map( A => n25_port, ZN => n202);
   U94 : AOI22_X1 port map( A1 => adj_sum_8_port, A2 => n14_port, B1 => 
                           n16_port, B2 => adj_final_mod_23_port, ZN => 
                           n25_port);
   U95 : INV_X1 port map( A => n26_port, ZN => n201);
   U96 : AOI22_X1 port map( A1 => adj_sum_7_port, A2 => n14_port, B1 => 
                           n16_port, B2 => adj_final_mod_22_port, ZN => 
                           n26_port);
   U97 : INV_X1 port map( A => n27_port, ZN => n200);
   U98 : AOI22_X1 port map( A1 => adj_sum_6_port, A2 => n14_port, B1 => 
                           n16_port, B2 => adj_final_mod_21_port, ZN => 
                           n27_port);
   U99 : INV_X1 port map( A => n32_port, ZN => n199);
   U100 : AOI22_X1 port map( A1 => adj_sum_5_port, A2 => n14_port, B1 => 
                           n16_port, B2 => adj_final_mod_20_port, ZN => 
                           n32_port);
   U101 : INV_X1 port map( A => n33_port, ZN => n198);
   U102 : AOI22_X1 port map( A1 => adj_sum_4_port, A2 => n14_port, B1 => 
                           n16_port, B2 => adj_final_mod_19_port, ZN => 
                           n33_port);
   U103 : INV_X1 port map( A => n34_port, ZN => n197);
   U104 : AOI22_X1 port map( A1 => adj_sum_3_port, A2 => n14_port, B1 => 
                           n16_port, B2 => adj_final_mod_18_port, ZN => 
                           n34_port);
   U105 : INV_X1 port map( A => n35_port, ZN => n196);
   U106 : AOI22_X1 port map( A1 => adj_sum_2_port, A2 => n14_port, B1 => 
                           n16_port, B2 => adj_final_mod_17_port, ZN => 
                           n35_port);
   U107 : INV_X1 port map( A => n36_port, ZN => n195);
   U108 : AOI22_X1 port map( A1 => adj_sum_1_port, A2 => n14_port, B1 => 
                           n16_port, B2 => adj_final_mod_16_port, ZN => 
                           n36_port);
   U109 : INV_X1 port map( A => n37_port, ZN => n194);
   U110 : AOI22_X1 port map( A1 => adj_sum_0_port, A2 => n14_port, B1 => 
                           n16_port, B2 => adj_final_mod_15_port, ZN => 
                           n37_port);
   U111 : AND2_X1 port map( A1 => a(0), A2 => n9_port, ZN => N9);
   U112 : AND3_X1 port map( A1 => b(15), A2 => n9_port, A3 => sign, ZN => N57);
   U113 : AND2_X1 port map( A1 => b(14), A2 => n9_port, ZN => N56);
   U114 : MUX2_X1 port map( A => b(13), B => e_b_16_port, S => n16_port, Z => 
                           N55);
   U115 : MUX2_X1 port map( A => b(12), B => e_b_15_port, S => n16_port, Z => 
                           N54);
   U116 : MUX2_X1 port map( A => b(11), B => e_b_14_port, S => n16_port, Z => 
                           N53);
   U117 : MUX2_X1 port map( A => b(10), B => e_b_13_port, S => n16_port, Z => 
                           N52);
   U118 : MUX2_X1 port map( A => b(9), B => e_b_12_port, S => n16_port, Z => 
                           N51);
   U119 : MUX2_X1 port map( A => b(8), B => e_b_11_port, S => n16_port, Z => 
                           N50);
   U120 : MUX2_X1 port map( A => b(7), B => e_b_10_port, S => n16_port, Z => 
                           N49);
   U121 : MUX2_X1 port map( A => b(6), B => e_b_9_port, S => n16_port, Z => N48
                           );
   U122 : MUX2_X1 port map( A => b(5), B => e_b_8_port, S => n16_port, Z => N47
                           );
   U123 : MUX2_X1 port map( A => b(4), B => e_b_7_port, S => n16_port, Z => N46
                           );
   U124 : MUX2_X1 port map( A => b(3), B => e_b_6_port, S => n16_port, Z => N45
                           );
   U125 : MUX2_X1 port map( A => b(2), B => e_b_5_port, S => n16_port, Z => N44
                           );
   U126 : MUX2_X1 port map( A => b(1), B => e_b_4_port, S => n16_port, Z => N43
                           );
   U127 : MUX2_X1 port map( A => b(0), B => e_b_3_port, S => n16_port, Z => N42
                           );
   U128 : NOR2_X1 port map( A1 => n58, A2 => n9_port, ZN => N41);
   U129 : OAI21_X1 port map( B1 => n87_port, B2 => n9_port, A => n39_port, ZN 
                           => N40);
   U130 : OAI21_X1 port map( B1 => n72_port, B2 => n9_port, A => n39_port, ZN 
                           => N39);
   U131 : OAI21_X1 port map( B1 => n86_port, B2 => n9_port, A => n39_port, ZN 
                           => N38);
   U132 : OAI21_X1 port map( B1 => n71_port, B2 => n9_port, A => n39_port, ZN 
                           => N37);
   U133 : OAI21_X1 port map( B1 => n85_port, B2 => n9_port, A => n39_port, ZN 
                           => N36);
   U134 : OAI21_X1 port map( B1 => n70_port, B2 => n9_port, A => n39_port, ZN 
                           => N35);
   U135 : OAI21_X1 port map( B1 => n84_port, B2 => n9_port, A => n39_port, ZN 
                           => N34);
   U136 : OAI21_X1 port map( B1 => n69, B2 => n9_port, A => n39_port, ZN => N33
                           );
   U137 : OAI21_X1 port map( B1 => n83_port, B2 => n9_port, A => n39_port, ZN 
                           => N32);
   U138 : OAI21_X1 port map( B1 => n68, B2 => n9_port, A => n39_port, ZN => N31
                           );
   U139 : OAI21_X1 port map( B1 => n82_port, B2 => n9_port, A => n39_port, ZN 
                           => N30);
   U140 : OAI21_X1 port map( B1 => n67, B2 => n9_port, A => n39_port, ZN => N29
                           );
   U141 : OAI21_X1 port map( B1 => n81_port, B2 => n9_port, A => n39_port, ZN 
                           => N28);
   U142 : OAI21_X1 port map( B1 => n66, B2 => n9_port, A => n39_port, ZN => N27
                           );
   U143 : OAI21_X1 port map( B1 => n80_port, B2 => n9_port, A => n39_port, ZN 
                           => N26);
   U144 : OAI21_X1 port map( B1 => n65, B2 => n9_port, A => n39_port, ZN => N25
                           );
   U145 : OAI21_X1 port map( B1 => n79_port, B2 => n9_port, A => n39_port, ZN 
                           => N24);
   U146 : NAND3_X1 port map( A1 => sign, A2 => n9_port, A3 => a(15), ZN => 
                           n39_port);
   U147 : MUX2_X1 port map( A => a(14), B => e_a_12_port, S => n16_port, Z => 
                           N23);
   U148 : MUX2_X1 port map( A => a(13), B => e_a_11_port, S => n16_port, Z => 
                           N22);
   U149 : MUX2_X1 port map( A => a(12), B => e_a_10_port, S => n16_port, Z => 
                           N21);
   U150 : MUX2_X1 port map( A => a(11), B => e_a_9_port, S => n16_port, Z => 
                           N20);
   U151 : MUX2_X1 port map( A => a(10), B => e_a_8_port, S => n16_port, Z => 
                           N19);
   U152 : MUX2_X1 port map( A => a(9), B => e_a_7_port, S => n16_port, Z => N18
                           );
   U153 : MUX2_X1 port map( A => a(8), B => e_a_6_port, S => n16_port, Z => N17
                           );
   U154 : MUX2_X1 port map( A => a(7), B => e_a_5_port, S => n16_port, Z => N16
                           );
   U155 : MUX2_X1 port map( A => a(6), B => e_a_4_port, S => n16_port, Z => N15
                           );
   U156 : MUX2_X1 port map( A => a(5), B => e_a_3_port, S => n16_port, Z => N14
                           );
   U157 : MUX2_X1 port map( A => a(4), B => e_a_2_port, S => n16_port, Z => N13
                           );
   U158 : MUX2_X1 port map( A => a(3), B => e_a_1_port, S => n16_port, Z => N12
                           );
   U159 : MUX2_X1 port map( A => a(2), B => e_a_0_port, S => n16_port, Z => N11
                           );
   U160 : AND2_X1 port map( A1 => a(1), A2 => n9_port, ZN => N10);
   U161 : INV_X1 port map( A => n16_port, ZN => n9_port);
   U162 : OAI211_X1 port map( C1 => n5, C2 => c_state_0_port, A => n7, B => 
                           n53_port, ZN => n38_port);
   U163 : AND3_X1 port map( A1 => n40_port, A2 => n41_port, A3 => n42_port, ZN 
                           => n7);
   U164 : INV_X1 port map( A => n43_port, ZN => n41_port);
   U165 : AOI21_X1 port map( B1 => n13_port, B2 => n55_port, A => n54_port, ZN 
                           => n43_port);
   U166 : NAND4_X1 port map( A1 => n42_port, A2 => n40_port, A3 => n13_port, A4
                           => n44_port, ZN => n5);
   U167 : AND2_X1 port map( A1 => n55_port, A2 => n54_port, ZN => n44_port);
   U168 : AND2_X1 port map( A1 => n45_port, A2 => n46_port, ZN => n40_port);
   U169 : NOR4_X1 port map( A1 => n47_port, A2 => c_state_16_port, A3 => 
                           c_state_14_port, A4 => c_state_15_port, ZN => 
                           n46_port);
   U170 : NAND4_X1 port map( A1 => n24_port, A2 => n23_port, A3 => n22_port, A4
                           => n12_port, ZN => n47_port);
   U171 : NOR4_X1 port map( A1 => n48_port, A2 => c_state_23_port, A3 => 
                           c_state_21_port, A4 => c_state_22_port, ZN => 
                           n45_port);
   U172 : NAND4_X1 port map( A1 => n31_port, A2 => n30_port, A3 => n29_port, A4
                           => n28_port, ZN => n48_port);
   U173 : AND2_X1 port map( A1 => n49_port, A2 => n50_port, ZN => n42_port);
   U174 : NOR4_X1 port map( A1 => n51_port, A2 => c_state_30_port, A3 => 
                           c_state_27_port, A4 => c_state_26_port, ZN => 
                           n50_port);
   U175 : NAND4_X1 port map( A1 => n60, A2 => n61, A3 => n62, A4 => n63, ZN => 
                           n51_port);
   U176 : NOR4_X1 port map( A1 => n52_port, A2 => c_state_6_port, A3 => 
                           c_state_8_port, A4 => c_state_7_port, ZN => n49_port
                           );
   U177 : NAND3_X1 port map( A1 => n57_port, A2 => n59, A3 => n56_port, ZN => 
                           n52_port);

end SYN_booth_mul_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Shifter_DATA_SIZE32 is

   port( l_r, l_a, s_r : in std_logic;  a, b : in std_logic_vector (31 downto 
         0);  o : out std_logic_vector (31 downto 0));

end Shifter_DATA_SIZE32;

architecture SYN_shifter_arch of Shifter_DATA_SIZE32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component Shifter_DATA_SIZE32_DW_rbsh_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component Shifter_DATA_SIZE32_DW_lbsh_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component Shifter_DATA_SIZE32_DW_sra_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component Shifter_DATA_SIZE32_DW_rash_0
      port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH
            : in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out
            std_logic_vector (31 downto 0));
   end component;
   
   component Shifter_DATA_SIZE32_DW_sla_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component Shifter_DATA_SIZE32_DW01_ash_0
      port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH
            : in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out
            std_logic_vector (31 downto 0));
   end component;
   
   signal N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, 
      N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37
      , N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, 
      N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66
      , N67, N68, N69, N70, N71, N72, N108, N109, N110, N111, N112, N113, N114,
      N115, N116, N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, 
      N127, N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, 
      N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, 
      N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, 
      N163, N164, N165, N166, N167, N168, N169, N170, N171, N205, N206, N207, 
      N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, 
      N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231, 
      N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, 
      N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, 
      N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267, 
      N268, n14_port, n15_port, n16_port, n17_port, n18_port, n19_port, n1, n2,
      n3, n4, n5, n6, n7, n8, n9_port, n10_port, n11_port, n12_port, n13_port, 
      n20_port, n21_port, n22_port, n23_port, n24_port, n25_port, n26_port, 
      n27_port, n28_port, n29_port, n30_port, n31_port, n32_port, n33_port, 
      n34_port, n35_port, n36_port, n37_port, n38_port, n39_port, n40_port, 
      n41_port, n42_port, n43_port, n44_port, n45_port, n46_port, n47_port, 
      n48_port, n49_port, n50_port, n51_port, n52_port, n53_port, n54_port, 
      n55_port, n56_port, n57_port, n58_port, n59_port, n60_port, n61_port, 
      n62_port, n63_port, n64_port, n65_port, n66_port, n67_port, n68_port, 
      n69_port, n70_port, n71_port, n72_port, n73, n74, n75, n76, n77, n78, n79
      , n80, n81, n82, n83, n84 : std_logic;

begin
   
   n14_port <= '0';
   n15_port <= '0';
   n16_port <= '0';
   n17_port <= '0';
   n18_port <= '0';
   n19_port <= '0';
   C93 : Shifter_DATA_SIZE32_DW01_ash_0 port map( A(31) => a(31), A(30) => 
                           a(30), A(29) => a(29), A(28) => a(28), A(27) => 
                           a(27), A(26) => a(26), A(25) => a(25), A(24) => 
                           a(24), A(23) => a(23), A(22) => a(22), A(21) => 
                           a(21), A(20) => a(20), A(19) => a(19), A(18) => 
                           a(18), A(17) => a(17), A(16) => a(16), A(15) => 
                           a(15), A(14) => a(14), A(13) => a(13), A(12) => 
                           a(12), A(11) => a(11), A(10) => a(10), A(9) => a(9),
                           A(8) => a(8), A(7) => a(7), A(6) => a(6), A(5) => 
                           a(5), A(4) => a(4), A(3) => a(3), A(2) => a(2), A(1)
                           => a(1), A(0) => a(0), DATA_TC => n14_port, SH(4) =>
                           n8, SH(3) => b(3), SH(2) => b(2), SH(1) => b(1), 
                           SH(0) => b(0), SH_TC => n14_port, B(31) => N268, 
                           B(30) => N267, B(29) => N266, B(28) => N265, B(27) 
                           => N264, B(26) => N263, B(25) => N262, B(24) => N261
                           , B(23) => N260, B(22) => N259, B(21) => N258, B(20)
                           => N257, B(19) => N256, B(18) => N255, B(17) => N254
                           , B(16) => N253, B(15) => N252, B(14) => N251, B(13)
                           => N250, B(12) => N249, B(11) => N248, B(10) => N247
                           , B(9) => N246, B(8) => N245, B(7) => N244, B(6) => 
                           N243, B(5) => N242, B(4) => N241, B(3) => N240, B(2)
                           => N239, B(1) => N238, B(0) => N237);
   C91 : Shifter_DATA_SIZE32_DW_sla_0 port map( A(31) => a(31), A(30) => a(30),
                           A(29) => a(29), A(28) => a(28), A(27) => a(27), 
                           A(26) => a(26), A(25) => a(25), A(24) => a(24), 
                           A(23) => a(23), A(22) => a(22), A(21) => a(21), 
                           A(20) => a(20), A(19) => a(19), A(18) => a(18), 
                           A(17) => a(17), A(16) => a(16), A(15) => a(15), 
                           A(14) => a(14), A(13) => a(13), A(12) => a(12), 
                           A(11) => a(11), A(10) => a(10), A(9) => a(9), A(8) 
                           => a(8), A(7) => a(7), A(6) => a(6), A(5) => a(5), 
                           A(4) => a(4), A(3) => a(3), A(2) => a(2), A(1) => 
                           a(1), A(0) => a(0), SH(4) => n8, SH(3) => b(3), 
                           SH(2) => b(2), SH(1) => b(1), SH(0) => b(0), SH_TC 
                           => n15_port, B(31) => N236, B(30) => N235, B(29) => 
                           N234, B(28) => N233, B(27) => N232, B(26) => N231, 
                           B(25) => N230, B(24) => N229, B(23) => N228, B(22) 
                           => N227, B(21) => N226, B(20) => N225, B(19) => N224
                           , B(18) => N223, B(17) => N222, B(16) => N221, B(15)
                           => N220, B(14) => N219, B(13) => N218, B(12) => N217
                           , B(11) => N216, B(10) => N215, B(9) => N214, B(8) 
                           => N213, B(7) => N212, B(6) => N211, B(5) => N210, 
                           B(4) => N209, B(3) => N208, B(2) => N207, B(1) => 
                           N206, B(0) => N205);
   C54 : Shifter_DATA_SIZE32_DW_rash_0 port map( A(31) => a(31), A(30) => a(30)
                           , A(29) => a(29), A(28) => a(28), A(27) => a(27), 
                           A(26) => a(26), A(25) => a(25), A(24) => a(24), 
                           A(23) => a(23), A(22) => a(22), A(21) => a(21), 
                           A(20) => a(20), A(19) => a(19), A(18) => a(18), 
                           A(17) => a(17), A(16) => a(16), A(15) => a(15), 
                           A(14) => a(14), A(13) => a(13), A(12) => a(12), 
                           A(11) => a(11), A(10) => a(10), A(9) => a(9), A(8) 
                           => a(8), A(7) => a(7), A(6) => a(6), A(5) => a(5), 
                           A(4) => a(4), A(3) => a(3), A(2) => a(2), A(1) => 
                           a(1), A(0) => a(0), DATA_TC => n16_port, SH(4) => n8
                           , SH(3) => b(3), SH(2) => b(2), SH(1) => b(1), SH(0)
                           => b(0), SH_TC => n16_port, B(31) => N171, B(30) => 
                           N170, B(29) => N169, B(28) => N168, B(27) => N167, 
                           B(26) => N166, B(25) => N165, B(24) => N164, B(23) 
                           => N163, B(22) => N162, B(21) => N161, B(20) => N160
                           , B(19) => N159, B(18) => N158, B(17) => N157, B(16)
                           => N156, B(15) => N155, B(14) => N154, B(13) => N153
                           , B(12) => N152, B(11) => N151, B(10) => N150, B(9) 
                           => N149, B(8) => N148, B(7) => N147, B(6) => N146, 
                           B(5) => N145, B(4) => N144, B(3) => N143, B(2) => 
                           N142, B(1) => N141, B(0) => N140);
   C52 : Shifter_DATA_SIZE32_DW_sra_0 port map( A(31) => a(31), A(30) => a(30),
                           A(29) => a(29), A(28) => a(28), A(27) => a(27), 
                           A(26) => a(26), A(25) => a(25), A(24) => a(24), 
                           A(23) => a(23), A(22) => a(22), A(21) => a(21), 
                           A(20) => a(20), A(19) => a(19), A(18) => a(18), 
                           A(17) => a(17), A(16) => a(16), A(15) => a(15), 
                           A(14) => a(14), A(13) => a(13), A(12) => a(12), 
                           A(11) => a(11), A(10) => a(10), A(9) => a(9), A(8) 
                           => a(8), A(7) => a(7), A(6) => a(6), A(5) => a(5), 
                           A(4) => a(4), A(3) => a(3), A(2) => a(2), A(1) => 
                           a(1), A(0) => a(0), SH(4) => n8, SH(3) => b(3), 
                           SH(2) => b(2), SH(1) => b(1), SH(0) => b(0), SH_TC 
                           => n17_port, B(31) => N139, B(30) => N138, B(29) => 
                           N137, B(28) => N136, B(27) => N135, B(26) => N134, 
                           B(25) => N133, B(24) => N132, B(23) => N131, B(22) 
                           => N130, B(21) => N129, B(20) => N128, B(19) => N127
                           , B(18) => N126, B(17) => N125, B(16) => N124, B(15)
                           => N123, B(14) => N122, B(13) => N121, B(12) => N120
                           , B(11) => N119, B(10) => N118, B(9) => N117, B(8) 
                           => N116, B(7) => N115, B(6) => N114, B(5) => N113, 
                           B(4) => N112, B(3) => N111, B(2) => N110, B(1) => 
                           N109, B(0) => N108);
   C12 : Shifter_DATA_SIZE32_DW_lbsh_0 port map( A(31) => a(31), A(30) => a(30)
                           , A(29) => a(29), A(28) => a(28), A(27) => a(27), 
                           A(26) => a(26), A(25) => a(25), A(24) => a(24), 
                           A(23) => a(23), A(22) => a(22), A(21) => a(21), 
                           A(20) => a(20), A(19) => a(19), A(18) => a(18), 
                           A(17) => a(17), A(16) => a(16), A(15) => a(15), 
                           A(14) => a(14), A(13) => a(13), A(12) => a(12), 
                           A(11) => a(11), A(10) => a(10), A(9) => a(9), A(8) 
                           => a(8), A(7) => a(7), A(6) => a(6), A(5) => a(5), 
                           A(4) => a(4), A(3) => a(3), A(2) => a(2), A(1) => 
                           a(1), A(0) => a(0), SH(4) => n8, SH(3) => b(3), 
                           SH(2) => b(2), SH(1) => b(1), SH(0) => b(0), SH_TC 
                           => n18_port, B(31) => N72, B(30) => N71, B(29) => 
                           N70, B(28) => N69, B(27) => N68, B(26) => N67, B(25)
                           => N66, B(24) => N65, B(23) => N64, B(22) => N63, 
                           B(21) => N62, B(20) => N61, B(19) => N60, B(18) => 
                           N59, B(17) => N58, B(16) => N57, B(15) => N56, B(14)
                           => N55, B(13) => N54, B(12) => N53, B(11) => N52, 
                           B(10) => N51, B(9) => N50, B(8) => N49, B(7) => N48,
                           B(6) => N47, B(5) => N46, B(4) => N45, B(3) => N44, 
                           B(2) => N43, B(1) => N42, B(0) => N41);
   C10 : Shifter_DATA_SIZE32_DW_rbsh_0 port map( A(31) => a(31), A(30) => a(30)
                           , A(29) => a(29), A(28) => a(28), A(27) => a(27), 
                           A(26) => a(26), A(25) => a(25), A(24) => a(24), 
                           A(23) => a(23), A(22) => a(22), A(21) => a(21), 
                           A(20) => a(20), A(19) => a(19), A(18) => a(18), 
                           A(17) => a(17), A(16) => a(16), A(15) => a(15), 
                           A(14) => a(14), A(13) => a(13), A(12) => a(12), 
                           A(11) => a(11), A(10) => a(10), A(9) => a(9), A(8) 
                           => a(8), A(7) => a(7), A(6) => a(6), A(5) => a(5), 
                           A(4) => a(4), A(3) => a(3), A(2) => a(2), A(1) => 
                           a(1), A(0) => a(0), SH(4) => n8, SH(3) => b(3), 
                           SH(2) => b(2), SH(1) => b(1), SH(0) => b(0), SH_TC 
                           => n19_port, B(31) => N40, B(30) => N39, B(29) => 
                           N38, B(28) => N37, B(27) => N36, B(26) => N35, B(25)
                           => N34, B(24) => N33, B(23) => N32, B(22) => N31, 
                           B(21) => N30, B(20) => N29, B(19) => N28, B(18) => 
                           N27, B(17) => N26, B(16) => N25, B(15) => N24, B(14)
                           => N23, B(13) => N22, B(12) => N21, B(11) => N20, 
                           B(10) => N19, B(9) => N18, B(8) => N17, B(7) => N16,
                           B(6) => N15, B(5) => N14, B(4) => N13, B(3) => N12, 
                           B(2) => N11, B(1) => N10, B(0) => N9);
   U5 : NOR2_X4 port map( A1 => n84, A2 => n82, ZN => n11_port);
   U6 : CLKBUF_X1 port map( A => n13_port, Z => n1);
   U7 : NOR2_X4 port map( A1 => n84, A2 => l_r, ZN => n12_port);
   U8 : OR3_X1 port map( A1 => l_r, A2 => s_r, A3 => l_a, ZN => n2);
   U9 : INV_X2 port map( A => n2, ZN => n3);
   U10 : OR3_X1 port map( A1 => l_a, A2 => s_r, A3 => n82, ZN => n4);
   U13 : INV_X2 port map( A => n4, ZN => n5);
   U14 : OR3_X1 port map( A1 => l_r, A2 => s_r, A3 => n83, ZN => n6);
   U15 : INV_X2 port map( A => n6, ZN => n7);
   U16 : CLKBUF_X3 port map( A => b(4), Z => n8);
   U17 : NAND2_X1 port map( A1 => n9_port, A2 => n10_port, ZN => o(9));
   U18 : AOI222_X1 port map( A1 => N214, A2 => n7, B1 => N149, B2 => n5, C1 => 
                           N246, C2 => n3, ZN => n10_port);
   U19 : AOI222_X1 port map( A1 => N18, A2 => n11_port, B1 => N50, B2 => 
                           n12_port, C1 => N117, C2 => n1, ZN => n9_port);
   U20 : NAND2_X1 port map( A1 => n20_port, A2 => n21_port, ZN => o(8));
   U21 : AOI222_X1 port map( A1 => N213, A2 => n7, B1 => N148, B2 => n5, C1 => 
                           N245, C2 => n3, ZN => n21_port);
   U22 : AOI222_X1 port map( A1 => N17, A2 => n11_port, B1 => N49, B2 => 
                           n12_port, C1 => N116, C2 => n1, ZN => n20_port);
   U23 : NAND2_X1 port map( A1 => n22_port, A2 => n23_port, ZN => o(7));
   U24 : AOI222_X1 port map( A1 => N212, A2 => n7, B1 => N147, B2 => n5, C1 => 
                           N244, C2 => n3, ZN => n23_port);
   U25 : AOI222_X1 port map( A1 => N16, A2 => n11_port, B1 => N48, B2 => 
                           n12_port, C1 => N115, C2 => n1, ZN => n22_port);
   U26 : NAND2_X1 port map( A1 => n24_port, A2 => n25_port, ZN => o(6));
   U27 : AOI222_X1 port map( A1 => N211, A2 => n7, B1 => N146, B2 => n5, C1 => 
                           N243, C2 => n3, ZN => n25_port);
   U28 : AOI222_X1 port map( A1 => N15, A2 => n11_port, B1 => N47, B2 => 
                           n12_port, C1 => N114, C2 => n1, ZN => n24_port);
   U29 : NAND2_X1 port map( A1 => n26_port, A2 => n27_port, ZN => o(5));
   U30 : AOI222_X1 port map( A1 => N210, A2 => n7, B1 => N145, B2 => n5, C1 => 
                           N242, C2 => n3, ZN => n27_port);
   U31 : AOI222_X1 port map( A1 => N14, A2 => n11_port, B1 => N46, B2 => 
                           n12_port, C1 => N113, C2 => n1, ZN => n26_port);
   U32 : NAND2_X1 port map( A1 => n28_port, A2 => n29_port, ZN => o(4));
   U33 : AOI222_X1 port map( A1 => N209, A2 => n7, B1 => N144, B2 => n5, C1 => 
                           N241, C2 => n3, ZN => n29_port);
   U34 : AOI222_X1 port map( A1 => N13, A2 => n11_port, B1 => N45, B2 => 
                           n12_port, C1 => N112, C2 => n1, ZN => n28_port);
   U35 : NAND2_X1 port map( A1 => n30_port, A2 => n31_port, ZN => o(3));
   U36 : AOI222_X1 port map( A1 => N208, A2 => n7, B1 => N143, B2 => n5, C1 => 
                           N240, C2 => n3, ZN => n31_port);
   U37 : AOI222_X1 port map( A1 => N12, A2 => n11_port, B1 => N44, B2 => 
                           n12_port, C1 => N111, C2 => n1, ZN => n30_port);
   U38 : NAND2_X1 port map( A1 => n32_port, A2 => n33_port, ZN => o(31));
   U39 : AOI222_X1 port map( A1 => N236, A2 => n7, B1 => N171, B2 => n5, C1 => 
                           N268, C2 => n3, ZN => n33_port);
   U40 : AOI222_X1 port map( A1 => N40, A2 => n11_port, B1 => N72, B2 => 
                           n12_port, C1 => N139, C2 => n1, ZN => n32_port);
   U41 : NAND2_X1 port map( A1 => n34_port, A2 => n35_port, ZN => o(30));
   U42 : AOI222_X1 port map( A1 => N235, A2 => n7, B1 => N170, B2 => n5, C1 => 
                           N267, C2 => n3, ZN => n35_port);
   U43 : AOI222_X1 port map( A1 => N39, A2 => n11_port, B1 => N71, B2 => 
                           n12_port, C1 => N138, C2 => n1, ZN => n34_port);
   U44 : NAND2_X1 port map( A1 => n36_port, A2 => n37_port, ZN => o(2));
   U45 : AOI222_X1 port map( A1 => N207, A2 => n7, B1 => N142, B2 => n5, C1 => 
                           N239, C2 => n3, ZN => n37_port);
   U46 : AOI222_X1 port map( A1 => N11, A2 => n11_port, B1 => N43, B2 => 
                           n12_port, C1 => N110, C2 => n1, ZN => n36_port);
   U47 : NAND2_X1 port map( A1 => n38_port, A2 => n39_port, ZN => o(29));
   U48 : AOI222_X1 port map( A1 => N234, A2 => n7, B1 => N169, B2 => n5, C1 => 
                           N266, C2 => n3, ZN => n39_port);
   U49 : AOI222_X1 port map( A1 => N38, A2 => n11_port, B1 => N70, B2 => 
                           n12_port, C1 => N137, C2 => n1, ZN => n38_port);
   U50 : NAND2_X1 port map( A1 => n40_port, A2 => n41_port, ZN => o(28));
   U51 : AOI222_X1 port map( A1 => N233, A2 => n7, B1 => N168, B2 => n5, C1 => 
                           N265, C2 => n3, ZN => n41_port);
   U52 : AOI222_X1 port map( A1 => N37, A2 => n11_port, B1 => N69, B2 => 
                           n12_port, C1 => N136, C2 => n1, ZN => n40_port);
   U53 : NAND2_X1 port map( A1 => n42_port, A2 => n43_port, ZN => o(27));
   U54 : AOI222_X1 port map( A1 => N232, A2 => n7, B1 => N167, B2 => n5, C1 => 
                           N264, C2 => n3, ZN => n43_port);
   U55 : AOI222_X1 port map( A1 => N36, A2 => n11_port, B1 => N68, B2 => 
                           n12_port, C1 => N135, C2 => n1, ZN => n42_port);
   U56 : NAND2_X1 port map( A1 => n44_port, A2 => n45_port, ZN => o(26));
   U57 : AOI222_X1 port map( A1 => N231, A2 => n7, B1 => N166, B2 => n5, C1 => 
                           N263, C2 => n3, ZN => n45_port);
   U58 : AOI222_X1 port map( A1 => N35, A2 => n11_port, B1 => N67, B2 => 
                           n12_port, C1 => N134, C2 => n1, ZN => n44_port);
   U59 : NAND2_X1 port map( A1 => n46_port, A2 => n47_port, ZN => o(25));
   U60 : AOI222_X1 port map( A1 => N230, A2 => n7, B1 => N165, B2 => n5, C1 => 
                           N262, C2 => n3, ZN => n47_port);
   U61 : AOI222_X1 port map( A1 => N34, A2 => n11_port, B1 => N66, B2 => 
                           n12_port, C1 => N133, C2 => n1, ZN => n46_port);
   U62 : NAND2_X1 port map( A1 => n48_port, A2 => n49_port, ZN => o(24));
   U63 : AOI222_X1 port map( A1 => N229, A2 => n7, B1 => N164, B2 => n5, C1 => 
                           N261, C2 => n3, ZN => n49_port);
   U64 : AOI222_X1 port map( A1 => N33, A2 => n11_port, B1 => N65, B2 => 
                           n12_port, C1 => N132, C2 => n1, ZN => n48_port);
   U65 : NAND2_X1 port map( A1 => n50_port, A2 => n51_port, ZN => o(23));
   U66 : AOI222_X1 port map( A1 => N228, A2 => n7, B1 => N163, B2 => n5, C1 => 
                           N260, C2 => n3, ZN => n51_port);
   U67 : AOI222_X1 port map( A1 => N32, A2 => n11_port, B1 => N64, B2 => 
                           n12_port, C1 => N131, C2 => n1, ZN => n50_port);
   U68 : NAND2_X1 port map( A1 => n52_port, A2 => n53_port, ZN => o(22));
   U69 : AOI222_X1 port map( A1 => N227, A2 => n7, B1 => N162, B2 => n5, C1 => 
                           N259, C2 => n3, ZN => n53_port);
   U70 : AOI222_X1 port map( A1 => N31, A2 => n11_port, B1 => N63, B2 => 
                           n12_port, C1 => N130, C2 => n1, ZN => n52_port);
   U71 : NAND2_X1 port map( A1 => n54_port, A2 => n55_port, ZN => o(21));
   U72 : AOI222_X1 port map( A1 => N226, A2 => n7, B1 => N161, B2 => n5, C1 => 
                           N258, C2 => n3, ZN => n55_port);
   U73 : AOI222_X1 port map( A1 => N30, A2 => n11_port, B1 => N62, B2 => 
                           n12_port, C1 => N129, C2 => n1, ZN => n54_port);
   U74 : NAND2_X1 port map( A1 => n56_port, A2 => n57_port, ZN => o(20));
   U75 : AOI222_X1 port map( A1 => N225, A2 => n7, B1 => N160, B2 => n5, C1 => 
                           N257, C2 => n3, ZN => n57_port);
   U76 : AOI222_X1 port map( A1 => N29, A2 => n11_port, B1 => N61, B2 => 
                           n12_port, C1 => N128, C2 => n1, ZN => n56_port);
   U77 : NAND2_X1 port map( A1 => n58_port, A2 => n59_port, ZN => o(1));
   U78 : AOI222_X1 port map( A1 => N206, A2 => n7, B1 => N141, B2 => n5, C1 => 
                           N238, C2 => n3, ZN => n59_port);
   U79 : AOI222_X1 port map( A1 => N10, A2 => n11_port, B1 => N42, B2 => 
                           n12_port, C1 => N109, C2 => n1, ZN => n58_port);
   U80 : NAND2_X1 port map( A1 => n60_port, A2 => n61_port, ZN => o(19));
   U81 : AOI222_X1 port map( A1 => N224, A2 => n7, B1 => N159, B2 => n5, C1 => 
                           N256, C2 => n3, ZN => n61_port);
   U82 : AOI222_X1 port map( A1 => N28, A2 => n11_port, B1 => N60, B2 => 
                           n12_port, C1 => N127, C2 => n1, ZN => n60_port);
   U83 : NAND2_X1 port map( A1 => n62_port, A2 => n63_port, ZN => o(18));
   U84 : AOI222_X1 port map( A1 => N223, A2 => n7, B1 => N158, B2 => n5, C1 => 
                           N255, C2 => n3, ZN => n63_port);
   U85 : AOI222_X1 port map( A1 => N27, A2 => n11_port, B1 => N59, B2 => 
                           n12_port, C1 => N126, C2 => n1, ZN => n62_port);
   U86 : NAND2_X1 port map( A1 => n64_port, A2 => n65_port, ZN => o(17));
   U87 : AOI222_X1 port map( A1 => N222, A2 => n7, B1 => N157, B2 => n5, C1 => 
                           N254, C2 => n3, ZN => n65_port);
   U88 : AOI222_X1 port map( A1 => N26, A2 => n11_port, B1 => N58, B2 => 
                           n12_port, C1 => N125, C2 => n1, ZN => n64_port);
   U89 : NAND2_X1 port map( A1 => n66_port, A2 => n67_port, ZN => o(16));
   U90 : AOI222_X1 port map( A1 => N221, A2 => n7, B1 => N156, B2 => n5, C1 => 
                           N253, C2 => n3, ZN => n67_port);
   U91 : AOI222_X1 port map( A1 => N25, A2 => n11_port, B1 => N57, B2 => 
                           n12_port, C1 => N124, C2 => n13_port, ZN => n66_port
                           );
   U92 : NAND2_X1 port map( A1 => n68_port, A2 => n69_port, ZN => o(15));
   U93 : AOI222_X1 port map( A1 => N220, A2 => n7, B1 => N155, B2 => n5, C1 => 
                           N252, C2 => n3, ZN => n69_port);
   U94 : AOI222_X1 port map( A1 => N24, A2 => n11_port, B1 => N56, B2 => 
                           n12_port, C1 => N123, C2 => n13_port, ZN => n68_port
                           );
   U95 : NAND2_X1 port map( A1 => n70_port, A2 => n71_port, ZN => o(14));
   U96 : AOI222_X1 port map( A1 => N219, A2 => n7, B1 => N154, B2 => n5, C1 => 
                           N251, C2 => n3, ZN => n71_port);
   U97 : AOI222_X1 port map( A1 => N23, A2 => n11_port, B1 => N55, B2 => 
                           n12_port, C1 => N122, C2 => n13_port, ZN => n70_port
                           );
   U98 : NAND2_X1 port map( A1 => n72_port, A2 => n73, ZN => o(13));
   U99 : AOI222_X1 port map( A1 => N218, A2 => n7, B1 => N153, B2 => n5, C1 => 
                           N250, C2 => n3, ZN => n73);
   U100 : AOI222_X1 port map( A1 => N22, A2 => n11_port, B1 => N54, B2 => 
                           n12_port, C1 => N121, C2 => n13_port, ZN => n72_port
                           );
   U101 : NAND2_X1 port map( A1 => n74, A2 => n75, ZN => o(12));
   U102 : AOI222_X1 port map( A1 => N217, A2 => n7, B1 => N152, B2 => n5, C1 =>
                           N249, C2 => n3, ZN => n75);
   U103 : AOI222_X1 port map( A1 => N21, A2 => n11_port, B1 => N53, B2 => 
                           n12_port, C1 => N120, C2 => n13_port, ZN => n74);
   U104 : NAND2_X1 port map( A1 => n76, A2 => n77, ZN => o(11));
   U105 : AOI222_X1 port map( A1 => N216, A2 => n7, B1 => N151, B2 => n5, C1 =>
                           N248, C2 => n3, ZN => n77);
   U106 : AOI222_X1 port map( A1 => N20, A2 => n11_port, B1 => N52, B2 => 
                           n12_port, C1 => N119, C2 => n13_port, ZN => n76);
   U107 : NAND2_X1 port map( A1 => n78, A2 => n79, ZN => o(10));
   U108 : AOI222_X1 port map( A1 => N215, A2 => n7, B1 => N150, B2 => n5, C1 =>
                           N247, C2 => n3, ZN => n79);
   U109 : AOI222_X1 port map( A1 => N19, A2 => n11_port, B1 => N51, B2 => 
                           n12_port, C1 => N118, C2 => n13_port, ZN => n78);
   U110 : NAND2_X1 port map( A1 => n80, A2 => n81, ZN => o(0));
   U111 : AOI222_X1 port map( A1 => N205, A2 => n7, B1 => N140, B2 => n5, C1 =>
                           N237, C2 => n3, ZN => n81);
   U112 : AOI222_X1 port map( A1 => N9, A2 => n11_port, B1 => N41, B2 => 
                           n12_port, C1 => N108, C2 => n1, ZN => n80);
   U113 : NOR3_X1 port map( A1 => n82, A2 => s_r, A3 => n83, ZN => n13_port);
   U114 : INV_X1 port map( A => l_a, ZN => n83);
   U115 : INV_X1 port map( A => l_r, ZN => n82);
   U116 : INV_X1 port map( A => s_r, ZN => n84);

end SYN_shifter_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity P4Adder_DATA_SIZE32_SPARSITY4_0 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end P4Adder_DATA_SIZE32_SPARSITY4_0;

architecture SYN_p4_adder_arch of P4Adder_DATA_SIZE32_SPARSITY4_0 is

   component AdderSumGenerator_DATA_SIZE32_SPARSITY4_0
      port( a, b : in std_logic_vector (31 downto 0);  cin : in 
            std_logic_vector (7 downto 0);  sum : out std_logic_vector (31 
            downto 0));
   end component;
   
   component P4CarryGenerator_DATA_SIZE32_SPARSITY4_0
      port( a, b : in std_logic_vector (31 downto 0);  cin : in std_logic;  
            cout : out std_logic_vector (7 downto 0));
   end component;
   
   signal carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port,
      carry_2_port, carry_1_port : std_logic;

begin
   
   CG0 : P4CarryGenerator_DATA_SIZE32_SPARSITY4_0 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), cin => cin, 
                           cout(7) => cout, cout(6) => carry_7_port, cout(5) =>
                           carry_6_port, cout(4) => carry_5_port, cout(3) => 
                           carry_4_port, cout(2) => carry_3_port, cout(1) => 
                           carry_2_port, cout(0) => carry_1_port);
   SG0 : AdderSumGenerator_DATA_SIZE32_SPARSITY4_0 port map( a(31) => a(31), 
                           a(30) => a(30), a(29) => a(29), a(28) => a(28), 
                           a(27) => a(27), a(26) => a(26), a(25) => a(25), 
                           a(24) => a(24), a(23) => a(23), a(22) => a(22), 
                           a(21) => a(21), a(20) => a(20), a(19) => a(19), 
                           a(18) => a(18), a(17) => a(17), a(16) => a(16), 
                           a(15) => a(15), a(14) => a(14), a(13) => a(13), 
                           a(12) => a(12), a(11) => a(11), a(10) => a(10), a(9)
                           => a(9), a(8) => a(8), a(7) => a(7), a(6) => a(6), 
                           a(5) => a(5), a(4) => a(4), a(3) => a(3), a(2) => 
                           a(2), a(1) => a(1), a(0) => a(0), b(31) => b(31), 
                           b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), cin(7) => 
                           carry_7_port, cin(6) => carry_6_port, cin(5) => 
                           carry_5_port, cin(4) => carry_4_port, cin(3) => 
                           carry_3_port, cin(2) => carry_2_port, cin(1) => 
                           carry_1_port, cin(0) => cin, sum(31) => s(31), 
                           sum(30) => s(30), sum(29) => s(29), sum(28) => s(28)
                           , sum(27) => s(27), sum(26) => s(26), sum(25) => 
                           s(25), sum(24) => s(24), sum(23) => s(23), sum(22) 
                           => s(22), sum(21) => s(21), sum(20) => s(20), 
                           sum(19) => s(19), sum(18) => s(18), sum(17) => s(17)
                           , sum(16) => s(16), sum(15) => s(15), sum(14) => 
                           s(14), sum(13) => s(13), sum(12) => s(12), sum(11) 
                           => s(11), sum(10) => s(10), sum(9) => s(9), sum(8) 
                           => s(8), sum(7) => s(7), sum(6) => s(6), sum(5) => 
                           s(5), sum(4) => s(4), sum(3) => s(3), sum(2) => s(2)
                           , sum(1) => s(1), sum(0) => s(0));

end SYN_p4_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux4_DATA_SIZE32 is

   port( sel : in std_logic_vector (1 downto 0);  din0, din1, din2, din3 : in 
         std_logic_vector (31 downto 0);  dout : out std_logic_vector (31 
         downto 0));

end Mux4_DATA_SIZE32;

architecture SYN_mux4_arch of Mux4_DATA_SIZE32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70 : std_logic;

begin
   
   U3 : NOR2_X4 port map( A1 => n69, A2 => sel(0), ZN => n4);
   U4 : NOR2_X4 port map( A1 => sel(0), A2 => sel(1), ZN => n6);
   U5 : NOR2_X4 port map( A1 => n69, A2 => n70, ZN => n5);
   U6 : NOR2_X4 port map( A1 => n70, A2 => sel(1), ZN => n3);
   U7 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => dout(31));
   U8 : AOI22_X1 port map( A1 => din1(31), A2 => n3, B1 => din2(31), B2 => n4, 
                           ZN => n2);
   U9 : AOI22_X1 port map( A1 => din3(31), A2 => n5, B1 => din0(31), B2 => n6, 
                           ZN => n1);
   U10 : NAND2_X1 port map( A1 => n7, A2 => n8, ZN => dout(24));
   U11 : AOI22_X1 port map( A1 => din1(24), A2 => n3, B1 => din2(24), B2 => n4,
                           ZN => n8);
   U12 : AOI22_X1 port map( A1 => din3(24), A2 => n5, B1 => din0(24), B2 => n6,
                           ZN => n7);
   U13 : NAND2_X1 port map( A1 => n9, A2 => n10, ZN => dout(23));
   U14 : AOI22_X1 port map( A1 => din1(23), A2 => n3, B1 => din2(23), B2 => n4,
                           ZN => n10);
   U15 : AOI22_X1 port map( A1 => din3(23), A2 => n5, B1 => din0(23), B2 => n6,
                           ZN => n9);
   U16 : NAND2_X1 port map( A1 => n11, A2 => n12, ZN => dout(22));
   U17 : AOI22_X1 port map( A1 => din1(22), A2 => n3, B1 => din2(22), B2 => n4,
                           ZN => n12);
   U18 : AOI22_X1 port map( A1 => din3(22), A2 => n5, B1 => din0(22), B2 => n6,
                           ZN => n11);
   U19 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => dout(21));
   U20 : AOI22_X1 port map( A1 => din1(21), A2 => n3, B1 => din2(21), B2 => n4,
                           ZN => n14);
   U21 : AOI22_X1 port map( A1 => din3(21), A2 => n5, B1 => din0(21), B2 => n6,
                           ZN => n13);
   U22 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => dout(20));
   U23 : AOI22_X1 port map( A1 => din1(20), A2 => n3, B1 => din2(20), B2 => n4,
                           ZN => n16);
   U24 : AOI22_X1 port map( A1 => din3(20), A2 => n5, B1 => din0(20), B2 => n6,
                           ZN => n15);
   U25 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => dout(19));
   U26 : AOI22_X1 port map( A1 => din1(19), A2 => n3, B1 => din2(19), B2 => n4,
                           ZN => n18);
   U27 : AOI22_X1 port map( A1 => din3(19), A2 => n5, B1 => din0(19), B2 => n6,
                           ZN => n17);
   U28 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => dout(18));
   U29 : AOI22_X1 port map( A1 => din1(18), A2 => n3, B1 => din2(18), B2 => n4,
                           ZN => n20);
   U30 : AOI22_X1 port map( A1 => din3(18), A2 => n5, B1 => din0(18), B2 => n6,
                           ZN => n19);
   U31 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => dout(17));
   U32 : AOI22_X1 port map( A1 => din1(17), A2 => n3, B1 => din2(17), B2 => n4,
                           ZN => n22);
   U33 : AOI22_X1 port map( A1 => din3(17), A2 => n5, B1 => din0(17), B2 => n6,
                           ZN => n21);
   U34 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => dout(16));
   U35 : AOI22_X1 port map( A1 => din1(16), A2 => n3, B1 => din2(16), B2 => n4,
                           ZN => n24);
   U36 : AOI22_X1 port map( A1 => din3(16), A2 => n5, B1 => din0(16), B2 => n6,
                           ZN => n23);
   U37 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => dout(15));
   U38 : AOI22_X1 port map( A1 => din1(15), A2 => n3, B1 => din2(15), B2 => n4,
                           ZN => n26);
   U39 : AOI22_X1 port map( A1 => din3(15), A2 => n5, B1 => din0(15), B2 => n6,
                           ZN => n25);
   U40 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => dout(14));
   U41 : AOI22_X1 port map( A1 => din1(14), A2 => n3, B1 => din2(14), B2 => n4,
                           ZN => n28);
   U42 : AOI22_X1 port map( A1 => din3(14), A2 => n5, B1 => din0(14), B2 => n6,
                           ZN => n27);
   U43 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => dout(13));
   U44 : AOI22_X1 port map( A1 => din1(13), A2 => n3, B1 => din2(13), B2 => n4,
                           ZN => n30);
   U45 : AOI22_X1 port map( A1 => din3(13), A2 => n5, B1 => din0(13), B2 => n6,
                           ZN => n29);
   U46 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => dout(12));
   U47 : AOI22_X1 port map( A1 => din1(12), A2 => n3, B1 => din2(12), B2 => n4,
                           ZN => n32);
   U48 : AOI22_X1 port map( A1 => din3(12), A2 => n5, B1 => din0(12), B2 => n6,
                           ZN => n31);
   U49 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => dout(11));
   U50 : AOI22_X1 port map( A1 => din1(11), A2 => n3, B1 => din2(11), B2 => n4,
                           ZN => n34);
   U51 : AOI22_X1 port map( A1 => din3(11), A2 => n5, B1 => din0(11), B2 => n6,
                           ZN => n33);
   U52 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => dout(10));
   U53 : AOI22_X1 port map( A1 => din1(10), A2 => n3, B1 => din2(10), B2 => n4,
                           ZN => n36);
   U54 : AOI22_X1 port map( A1 => din3(10), A2 => n5, B1 => din0(10), B2 => n6,
                           ZN => n35);
   U55 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => dout(9));
   U56 : AOI22_X1 port map( A1 => din1(9), A2 => n3, B1 => din2(9), B2 => n4, 
                           ZN => n38);
   U57 : AOI22_X1 port map( A1 => din3(9), A2 => n5, B1 => din0(9), B2 => n6, 
                           ZN => n37);
   U58 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => dout(8));
   U59 : AOI22_X1 port map( A1 => din1(8), A2 => n3, B1 => din2(8), B2 => n4, 
                           ZN => n40);
   U60 : AOI22_X1 port map( A1 => din3(8), A2 => n5, B1 => din0(8), B2 => n6, 
                           ZN => n39);
   U61 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => dout(7));
   U62 : AOI22_X1 port map( A1 => din1(7), A2 => n3, B1 => din2(7), B2 => n4, 
                           ZN => n42);
   U63 : AOI22_X1 port map( A1 => din3(7), A2 => n5, B1 => din0(7), B2 => n6, 
                           ZN => n41);
   U64 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => dout(6));
   U65 : AOI22_X1 port map( A1 => din1(6), A2 => n3, B1 => din2(6), B2 => n4, 
                           ZN => n44);
   U66 : AOI22_X1 port map( A1 => din3(6), A2 => n5, B1 => din0(6), B2 => n6, 
                           ZN => n43);
   U67 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => dout(5));
   U68 : AOI22_X1 port map( A1 => din1(5), A2 => n3, B1 => din2(5), B2 => n4, 
                           ZN => n46);
   U69 : AOI22_X1 port map( A1 => din3(5), A2 => n5, B1 => din0(5), B2 => n6, 
                           ZN => n45);
   U70 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => dout(4));
   U71 : AOI22_X1 port map( A1 => din1(4), A2 => n3, B1 => din2(4), B2 => n4, 
                           ZN => n48);
   U72 : AOI22_X1 port map( A1 => din3(4), A2 => n5, B1 => din0(4), B2 => n6, 
                           ZN => n47);
   U73 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => dout(3));
   U74 : AOI22_X1 port map( A1 => din1(3), A2 => n3, B1 => din2(3), B2 => n4, 
                           ZN => n50);
   U75 : AOI22_X1 port map( A1 => din3(3), A2 => n5, B1 => din0(3), B2 => n6, 
                           ZN => n49);
   U76 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => dout(2));
   U77 : AOI22_X1 port map( A1 => din1(2), A2 => n3, B1 => din2(2), B2 => n4, 
                           ZN => n52);
   U78 : AOI22_X1 port map( A1 => din3(2), A2 => n5, B1 => din0(2), B2 => n6, 
                           ZN => n51);
   U79 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => dout(1));
   U80 : AOI22_X1 port map( A1 => din1(1), A2 => n3, B1 => din2(1), B2 => n4, 
                           ZN => n54);
   U81 : AOI22_X1 port map( A1 => din3(1), A2 => n5, B1 => din0(1), B2 => n6, 
                           ZN => n53);
   U82 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => dout(0));
   U83 : AOI22_X1 port map( A1 => din1(0), A2 => n3, B1 => din2(0), B2 => n4, 
                           ZN => n56);
   U84 : AOI22_X1 port map( A1 => din3(0), A2 => n5, B1 => din0(0), B2 => n6, 
                           ZN => n55);
   U85 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => dout(30));
   U86 : AOI22_X1 port map( A1 => din1(30), A2 => n3, B1 => din2(30), B2 => n4,
                           ZN => n58);
   U87 : AOI22_X1 port map( A1 => din3(30), A2 => n5, B1 => din0(30), B2 => n6,
                           ZN => n57);
   U88 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => dout(29));
   U89 : AOI22_X1 port map( A1 => din1(29), A2 => n3, B1 => din2(29), B2 => n4,
                           ZN => n60);
   U90 : AOI22_X1 port map( A1 => din3(29), A2 => n5, B1 => din0(29), B2 => n6,
                           ZN => n59);
   U91 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => dout(28));
   U92 : AOI22_X1 port map( A1 => din1(28), A2 => n3, B1 => din2(28), B2 => n4,
                           ZN => n62);
   U93 : AOI22_X1 port map( A1 => din3(28), A2 => n5, B1 => din0(28), B2 => n6,
                           ZN => n61);
   U94 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => dout(27));
   U95 : AOI22_X1 port map( A1 => din1(27), A2 => n3, B1 => din2(27), B2 => n4,
                           ZN => n64);
   U96 : AOI22_X1 port map( A1 => din3(27), A2 => n5, B1 => din0(27), B2 => n6,
                           ZN => n63);
   U97 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => dout(26));
   U98 : AOI22_X1 port map( A1 => din1(26), A2 => n3, B1 => din2(26), B2 => n4,
                           ZN => n66);
   U99 : AOI22_X1 port map( A1 => din3(26), A2 => n5, B1 => din0(26), B2 => n6,
                           ZN => n65);
   U100 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => dout(25));
   U101 : AOI22_X1 port map( A1 => din1(25), A2 => n3, B1 => din2(25), B2 => n4
                           , ZN => n68);
   U102 : AOI22_X1 port map( A1 => din3(25), A2 => n5, B1 => din0(25), B2 => n6
                           , ZN => n67);
   U103 : INV_X1 port map( A => sel(0), ZN => n70);
   U104 : INV_X1 port map( A => sel(1), ZN => n69);

end SYN_mux4_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Div_DATA_SIZE32_DIV_STAGE34_SQRT_STAGE18 is

   port( rst, clk, en, lock, sign, func : in std_logic;  a, b : in 
         std_logic_vector (31 downto 0);  o : out std_logic_vector (31 downto 
         0));

end Div_DATA_SIZE32_DIV_STAGE34_SQRT_STAGE18;

architecture SYN_div_arch of Div_DATA_SIZE32_DIV_STAGE34_SQRT_STAGE18 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X8
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X4
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X2
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component Div_DATA_SIZE32_DIV_STAGE34_SQRT_STAGE18_DW01_inc_0
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component AddSub_DATA_SIZE32_2
      port( as : in std_logic;  a, b : in std_logic_vector (31 downto 0);  re :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;
   
   component Sipo_DATA_SIZE32
      port( rst, en, clk, din : in std_logic;  dout : out std_logic_vector (31 
            downto 0));
   end component;
   
   component Reg_DATA_SIZE64
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (63 downto 
            0);  dout : out std_logic_vector (63 downto 0));
   end component;
   
   component AddSub_DATA_SIZE64
      port( as : in std_logic;  a, b : in std_logic_vector (63 downto 0);  re :
            out std_logic_vector (63 downto 0);  cout : out std_logic);
   end component;
   
   component Mux_DATA_SIZE64
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (63 downto 0)
            ;  dout : out std_logic_vector (63 downto 0));
   end component;
   
   component AddSub_DATA_SIZE32_3
      port( as : in std_logic;  a, b : in std_logic_vector (31 downto 0);  re :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;
   
   component AddSub_DATA_SIZE32_0
      port( as : in std_logic;  a, b : in std_logic_vector (31 downto 0);  re :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic0_port, a_mod_63_port, a_mod_62_port, a_mod_61_port, 
      a_mod_60_port, a_mod_59_port, a_mod_58_port, a_mod_57_port, a_mod_56_port
      , a_mod_55_port, a_mod_54_port, a_mod_53_port, a_mod_52_port, 
      a_mod_51_port, a_mod_50_port, a_mod_49_port, a_mod_48_port, a_mod_47_port
      , a_mod_46_port, a_mod_45_port, a_mod_44_port, a_mod_43_port, 
      a_mod_42_port, a_mod_41_port, a_mod_40_port, a_mod_39_port, a_mod_38_port
      , a_mod_37_port, a_mod_36_port, a_mod_35_port, a_mod_34_port, 
      a_mod_33_port, a_mod_32_port, a_mod_31_port, a_mod_30_port, a_mod_29_port
      , a_mod_28_port, a_mod_27_port, a_mod_26_port, a_mod_25_port, 
      a_mod_24_port, a_mod_23_port, a_mod_22_port, a_mod_21_port, a_mod_20_port
      , a_mod_19_port, a_mod_18_port, a_mod_17_port, a_mod_16_port, 
      a_mod_15_port, a_mod_14_port, a_mod_13_port, a_mod_12_port, a_mod_11_port
      , a_mod_10_port, a_mod_9_port, a_mod_8_port, a_mod_7_port, a_mod_6_port, 
      a_mod_5_port, a_mod_4_port, a_mod_3_port, a_mod_2_port, a_mod_1_port, 
      a_mod_0_port, inv_q_flag_mod, inv_a_flag, inv_b_flag, a_adj_31_port, 
      a_adj_30_port, a_adj_29_port, a_adj_28_port, a_adj_27_port, a_adj_26_port
      , a_adj_25_port, a_adj_24_port, a_adj_23_port, a_adj_22_port, 
      a_adj_21_port, a_adj_20_port, a_adj_19_port, a_adj_18_port, a_adj_17_port
      , a_adj_16_port, a_adj_15_port, a_adj_14_port, a_adj_13_port, 
      a_adj_12_port, a_adj_11_port, a_adj_10_port, a_adj_9_port, a_adj_8_port, 
      a_adj_7_port, a_adj_6_port, a_adj_5_port, a_adj_4_port, a_adj_3_port, 
      a_adj_2_port, a_adj_1_port, a_adj_0_port, b_adj_31_port, b_adj_30_port, 
      b_adj_29_port, b_adj_28_port, b_adj_27_port, b_adj_26_port, b_adj_25_port
      , b_adj_24_port, b_adj_23_port, b_adj_22_port, b_adj_21_port, 
      b_adj_20_port, b_adj_19_port, b_adj_18_port, b_adj_17_port, b_adj_16_port
      , b_adj_15_port, b_adj_14_port, b_adj_13_port, b_adj_12_port, 
      b_adj_11_port, b_adj_10_port, b_adj_9_port, b_adj_8_port, b_adj_7_port, 
      b_adj_6_port, b_adj_5_port, b_adj_4_port, b_adj_3_port, b_adj_2_port, 
      b_adj_1_port, b_adj_0_port, r_63_port, r_62_port, r_61_port, r_60_port, 
      r_59_port, r_58_port, r_57_port, r_56_port, r_55_port, r_54_port, 
      r_53_port, r_52_port, r_51_port, r_50_port, r_49_port, r_48_port, 
      r_47_port, r_46_port, r_45_port, r_44_port, r_43_port, r_42_port, 
      r_41_port, r_40_port, r_39_port, r_38_port, r_37_port, r_36_port, 
      r_35_port, r_34_port, r_33_port, r_32_port, r_31_port, r_30_port, 
      r_29_port, r_28_port, r_27_port, r_26_port, r_25_port, r_24_port, 
      r_23_port, r_22_port, r_21_port, r_20_port, r_19_port, r_18_port, 
      r_17_port, r_16_port, r_15_port, r_14_port, r_13_port, r_12_port, 
      r_11_port, r_10_port, r_9_port, r_8_port, r_7_port, r_6_port, r_5_port, 
      r_4_port, r_3_port, r_2_port, r_1_port, r_0_port, a_mux_63_port, 
      a_mux_62_port, a_mux_61_port, a_mux_60_port, a_mux_59_port, a_mux_58_port
      , a_mux_57_port, a_mux_56_port, a_mux_55_port, a_mux_54_port, 
      a_mux_53_port, a_mux_52_port, a_mux_51_port, a_mux_50_port, a_mux_49_port
      , a_mux_48_port, a_mux_47_port, a_mux_46_port, a_mux_45_port, 
      a_mux_44_port, a_mux_43_port, a_mux_42_port, a_mux_41_port, a_mux_40_port
      , a_mux_39_port, a_mux_38_port, a_mux_37_port, a_mux_36_port, 
      a_mux_35_port, a_mux_34_port, a_mux_33_port, a_mux_32_port, a_mux_31_port
      , a_mux_30_port, a_mux_29_port, a_mux_28_port, a_mux_27_port, 
      a_mux_26_port, a_mux_25_port, a_mux_24_port, a_mux_23_port, a_mux_22_port
      , a_mux_21_port, a_mux_20_port, a_mux_19_port, a_mux_18_port, 
      a_mux_17_port, a_mux_16_port, a_mux_15_port, a_mux_14_port, a_mux_13_port
      , a_mux_12_port, a_mux_11_port, a_mux_10_port, a_mux_9_port, a_mux_8_port
      , a_mux_7_port, a_mux_6_port, a_mux_5_port, a_mux_4_port, a_mux_3_port, 
      a_mux_2_port, a_mux_1_port, a_mux_0_port, not_r_sign, a_shf_63_port, 
      a_shf_62_port, a_shf_61_port, a_shf_60_port, a_shf_59_port, a_shf_58_port
      , a_shf_57_port, a_shf_56_port, a_shf_55_port, a_shf_54_port, 
      a_shf_53_port, a_shf_52_port, a_shf_51_port, a_shf_50_port, a_shf_49_port
      , a_shf_48_port, a_shf_47_port, a_shf_46_port, a_shf_45_port, 
      a_shf_44_port, a_shf_43_port, a_shf_42_port, a_shf_41_port, a_shf_40_port
      , a_shf_39_port, a_shf_38_port, a_shf_37_port, a_shf_36_port, 
      a_shf_35_port, a_shf_34_port, a_shf_33_port, a_shf_32_port, a_shf_31_port
      , a_shf_30_port, a_shf_29_port, a_shf_28_port, a_shf_27_port, 
      a_shf_26_port, a_shf_25_port, a_shf_24_port, a_shf_23_port, a_shf_22_port
      , a_shf_21_port, a_shf_20_port, a_shf_19_port, a_shf_18_port, 
      a_shf_17_port, a_shf_16_port, a_shf_15_port, a_shf_14_port, a_shf_13_port
      , a_shf_12_port, a_shf_11_port, a_shf_10_port, a_shf_9_port, a_shf_8_port
      , a_shf_7_port, a_shf_6_port, a_shf_5_port, a_shf_4_port, a_shf_3_port, 
      a_shf_2_port, a_shf_1_port, q_31_port, q_30_port, b_shf_sqrt_63_port, 
      b_shf_sqrt_62_port, b_shf_sqrt_61_port, b_shf_sqrt_60_port, 
      b_shf_sqrt_59_port, b_shf_sqrt_58_port, b_shf_sqrt_57_port, 
      b_shf_sqrt_56_port, b_shf_sqrt_55_port, b_shf_sqrt_54_port, 
      b_shf_sqrt_53_port, b_shf_sqrt_52_port, b_shf_sqrt_51_port, 
      b_shf_sqrt_50_port, b_shf_sqrt_49_port, b_shf_sqrt_48_port, 
      b_shf_sqrt_47_port, b_shf_sqrt_46_port, b_shf_sqrt_45_port, 
      b_shf_sqrt_44_port, b_shf_sqrt_43_port, b_shf_sqrt_42_port, 
      b_shf_sqrt_41_port, b_shf_sqrt_40_port, b_shf_sqrt_39_port, 
      b_shf_sqrt_38_port, b_shf_sqrt_37_port, b_shf_sqrt_36_port, 
      b_shf_sqrt_35_port, b_shf_sqrt_34_port, b_shf_63_port, b_shf_62_port, 
      b_shf_61_port, b_shf_60_port, b_shf_59_port, b_shf_58_port, b_shf_57_port
      , b_shf_56_port, b_shf_55_port, b_shf_54_port, b_shf_53_port, 
      b_shf_52_port, b_shf_51_port, b_shf_50_port, b_shf_49_port, b_shf_48_port
      , b_shf_47_port, b_shf_46_port, b_shf_45_port, b_shf_44_port, 
      b_shf_43_port, b_shf_42_port, b_shf_41_port, b_shf_40_port, b_shf_39_port
      , b_shf_38_port, b_shf_37_port, b_shf_36_port, b_shf_35_port, 
      b_shf_34_port, b_shf_33_port, b_shf_32_port, b_shf_31_port, b_shf_30_port
      , b_shf_29_port, b_shf_28_port, b_shf_27_port, b_shf_26_port, 
      b_shf_25_port, b_shf_24_port, b_shf_23_port, b_shf_22_port, b_shf_21_port
      , b_shf_20_port, b_shf_19_port, b_shf_18_port, b_shf_17_port, 
      b_shf_16_port, b_shf_15_port, b_shf_14_port, b_shf_13_port, b_shf_12_port
      , b_shf_11_port, b_shf_10_port, b_shf_9_port, b_shf_8_port, b_shf_7_port,
      b_shf_6_port, b_shf_5_port, b_shf_4_port, b_shf_3_port, b_shf_2_port, 
      b_shf_1_port, b_shf_0_port, r_es_63_port, r_es_62_port, r_es_61_port, 
      r_es_60_port, r_es_59_port, r_es_58_port, r_es_57_port, r_es_56_port, 
      r_es_55_port, r_es_54_port, r_es_53_port, r_es_52_port, r_es_51_port, 
      r_es_50_port, r_es_49_port, r_es_48_port, r_es_47_port, r_es_46_port, 
      r_es_45_port, r_es_44_port, r_es_43_port, r_es_42_port, r_es_41_port, 
      r_es_40_port, r_es_39_port, r_es_38_port, r_es_37_port, r_es_36_port, 
      r_es_35_port, r_es_34_port, r_es_33_port, r_es_32_port, r_es_31_port, 
      r_es_30_port, r_es_29_port, r_es_28_port, r_es_27_port, r_es_26_port, 
      r_es_25_port, r_es_24_port, r_es_23_port, r_es_22_port, r_es_21_port, 
      r_es_20_port, r_es_19_port, r_es_18_port, r_es_17_port, r_es_16_port, 
      r_es_15_port, r_es_14_port, r_es_13_port, r_es_12_port, r_es_11_port, 
      r_es_10_port, r_es_9_port, r_es_8_port, r_es_7_port, r_es_6_port, 
      r_es_5_port, r_es_4_port, r_es_3_port, r_es_2_port, r_es_1_port, 
      r_es_0_port, en_r, not_r_es_sign, n_state_31_port, n_state_30_port, 
      n_state_29_port, n_state_28_port, n_state_27_port, n_state_26_port, 
      n_state_25_port, n_state_24_port, n_state_23_port, n_state_22_port, 
      n_state_21_port, n_state_20_port, n_state_19_port, n_state_18_port, 
      n_state_17_port, n_state_16_port, n_state_15_port, n_state_14_port, 
      n_state_13_port, n_state_12_port, n_state_11_port, n_state_10_port, 
      n_state_9_port, n_state_8_port, n_state_7_port, n_state_6_port, 
      n_state_5_port, n_state_4_port, n_state_3_port, n_state_2_port, 
      n_state_1_port, n_state_0_port, c_state_31_port, c_state_30_port, 
      c_state_29_port, c_state_28_port, c_state_27_port, c_state_26_port, 
      c_state_25_port, c_state_24_port, c_state_23_port, c_state_22_port, 
      c_state_21_port, c_state_20_port, c_state_19_port, c_state_18_port, 
      c_state_17_port, c_state_16_port, c_state_15_port, c_state_14_port, 
      c_state_13_port, c_state_12_port, c_state_11_port, c_state_10_port, 
      c_state_9_port, c_state_8_port, c_state_7_port, c_state_6_port, 
      c_state_5_port, c_state_4_port, c_state_3_port, c_state_2_port, 
      c_state_1_port, c_state_0_port, N17, N18, N19, N20, N21, N22, N23, N24, 
      N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39
      , N40, N41, N42, N43, N44, N45, N46, N47, N48, net3927, net3928, net3929,
      net3930, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307
      , n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
      n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, 
      n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, 
      n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, 
      n356, n357, n358, n359, n360, n361, n362, n371, n372, n373, n374, n1, n2,
      n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17_port, 
      n18_port, n19_port, n20_port, n21_port, n22_port, n23_port, n24_port, 
      n25_port, n26_port, n27_port, n28_port, n29_port, n30_port, n31_port, 
      n32_port, n33_port, n34_port, n35_port, n36_port, n37_port, n38_port, 
      n39_port, n40_port, n41_port, n42_port, n43_port, n44_port, n45_port, 
      n46_port, n47_port, n48_port, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
      n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86
      , net108616, net108617, net108618, net108619, net108620, net108621, 
      net108622, net108623, net108624, net108625, net108626, net108627, 
      net108628, net108629, net108630, net108631, net108632, net108633, 
      net108634, net108635, net108636, net108637, net108638, net108639, 
      net108640, net108641, net108642, net108643, net108644, net108645, 
      net108646, net108647, net108648, net108649, net108650, net108651, 
      net108652, net108653, net108654, net108655, net108656, net108657, 
      net108658, net108659, net108660, net108661, net108662, net108663, 
      net108664, net108665, net108666, net108667, net108668, net108669, 
      net108670, net108671, net108672, net108673, net108674, net108675, 
      net108676, net108677, net108678, net108679, net108680, net108681, 
      net108682, net108683, net108684, net108685, net108686, net108687, 
      net108688, net108689, net108690 : std_logic;

begin
   
   X_Logic0_port <= '0';
   c_state_reg_0_inst : DFFR_X1 port map( D => n_state_0_port, CK => clk, RN =>
                           rst, Q => c_state_0_port, QN => n362);
   c_state_reg_10_inst : DFFR_X1 port map( D => n_state_10_port, CK => clk, RN 
                           => rst, Q => c_state_10_port, QN => net108690);
   c_state_reg_1_inst : DFFR_X1 port map( D => n_state_1_port, CK => clk, RN =>
                           rst, Q => c_state_1_port, QN => n373);
   c_state_reg_2_inst : DFFR_X1 port map( D => n_state_2_port, CK => clk, RN =>
                           rst, Q => c_state_2_port, QN => n77);
   c_state_reg_3_inst : DFFR_X1 port map( D => n_state_3_port, CK => clk, RN =>
                           rst, Q => c_state_3_port, QN => n78);
   c_state_reg_4_inst : DFFR_X1 port map( D => n_state_4_port, CK => clk, RN =>
                           rst, Q => c_state_4_port, QN => n76);
   c_state_reg_5_inst : DFFR_X1 port map( D => n_state_5_port, CK => clk, RN =>
                           rst, Q => c_state_5_port, QN => n82);
   c_state_reg_6_inst : DFFR_X1 port map( D => n_state_6_port, CK => clk, RN =>
                           rst, Q => c_state_6_port, QN => n79);
   c_state_reg_7_inst : DFFR_X1 port map( D => n_state_7_port, CK => clk, RN =>
                           rst, Q => c_state_7_port, QN => n80);
   c_state_reg_8_inst : DFFR_X1 port map( D => n_state_8_port, CK => clk, RN =>
                           rst, Q => c_state_8_port, QN => n81);
   c_state_reg_9_inst : DFFR_X1 port map( D => n_state_9_port, CK => clk, RN =>
                           rst, Q => c_state_9_port, QN => net108689);
   c_state_reg_11_inst : DFFR_X1 port map( D => n_state_11_port, CK => clk, RN 
                           => rst, Q => c_state_11_port, QN => net108688);
   c_state_reg_12_inst : DFFR_X1 port map( D => n_state_12_port, CK => clk, RN 
                           => rst, Q => c_state_12_port, QN => net108687);
   c_state_reg_13_inst : DFFR_X1 port map( D => n_state_13_port, CK => clk, RN 
                           => rst, Q => c_state_13_port, QN => n74);
   c_state_reg_14_inst : DFFR_X1 port map( D => n_state_14_port, CK => clk, RN 
                           => rst, Q => c_state_14_port, QN => n75);
   c_state_reg_15_inst : DFFR_X1 port map( D => n_state_15_port, CK => clk, RN 
                           => rst, Q => c_state_15_port, QN => n73);
   c_state_reg_16_inst : DFFR_X1 port map( D => n_state_16_port, CK => clk, RN 
                           => rst, Q => c_state_16_port, QN => net108686);
   c_state_reg_17_inst : DFFR_X1 port map( D => n_state_17_port, CK => clk, RN 
                           => rst, Q => c_state_17_port, QN => net108685);
   c_state_reg_18_inst : DFFR_X1 port map( D => n_state_18_port, CK => clk, RN 
                           => rst, Q => c_state_18_port, QN => n371);
   c_state_reg_19_inst : DFFR_X1 port map( D => n_state_19_port, CK => clk, RN 
                           => rst, Q => c_state_19_port, QN => n372);
   c_state_reg_20_inst : DFFR_X1 port map( D => n_state_20_port, CK => clk, RN 
                           => rst, Q => c_state_20_port, QN => n374);
   c_state_reg_21_inst : DFFR_X1 port map( D => n_state_21_port, CK => clk, RN 
                           => rst, Q => c_state_21_port, QN => net108684);
   c_state_reg_22_inst : DFFR_X1 port map( D => n_state_22_port, CK => clk, RN 
                           => rst, Q => c_state_22_port, QN => n86);
   c_state_reg_23_inst : DFFR_X1 port map( D => n_state_23_port, CK => clk, RN 
                           => rst, Q => c_state_23_port, QN => net108683);
   c_state_reg_24_inst : DFFR_X1 port map( D => n_state_24_port, CK => clk, RN 
                           => rst, Q => c_state_24_port, QN => net108682);
   c_state_reg_25_inst : DFFR_X1 port map( D => n_state_25_port, CK => clk, RN 
                           => rst, Q => c_state_25_port, QN => n83);
   c_state_reg_26_inst : DFFR_X1 port map( D => n_state_26_port, CK => clk, RN 
                           => rst, Q => c_state_26_port, QN => n84);
   c_state_reg_27_inst : DFFR_X1 port map( D => n_state_27_port, CK => clk, RN 
                           => rst, Q => c_state_27_port, QN => n85);
   c_state_reg_28_inst : DFFR_X1 port map( D => n_state_28_port, CK => clk, RN 
                           => rst, Q => c_state_28_port, QN => net108681);
   c_state_reg_29_inst : DFFR_X1 port map( D => n_state_29_port, CK => clk, RN 
                           => rst, Q => c_state_29_port, QN => net108680);
   c_state_reg_30_inst : DFFR_X1 port map( D => n_state_30_port, CK => clk, RN 
                           => rst, Q => c_state_30_port, QN => net108679);
   c_state_reg_31_inst : DFFR_X1 port map( D => n_state_31_port, CK => clk, RN 
                           => rst, Q => c_state_31_port, QN => n72);
   a_mod_reg_0_inst : DFF_X1 port map( D => n361, CK => clk, Q => a_mod_0_port,
                           QN => net108678);
   a_mod_reg_1_inst : DFF_X1 port map( D => n360, CK => clk, Q => a_mod_1_port,
                           QN => net108677);
   a_mod_reg_2_inst : DFF_X1 port map( D => n359, CK => clk, Q => a_mod_2_port,
                           QN => net108676);
   a_mod_reg_3_inst : DFF_X1 port map( D => n358, CK => clk, Q => a_mod_3_port,
                           QN => net108675);
   a_mod_reg_4_inst : DFF_X1 port map( D => n357, CK => clk, Q => a_mod_4_port,
                           QN => net108674);
   a_mod_reg_5_inst : DFF_X1 port map( D => n356, CK => clk, Q => a_mod_5_port,
                           QN => net108673);
   a_mod_reg_6_inst : DFF_X1 port map( D => n355, CK => clk, Q => a_mod_6_port,
                           QN => net108672);
   a_mod_reg_7_inst : DFF_X1 port map( D => n354, CK => clk, Q => a_mod_7_port,
                           QN => net108671);
   a_mod_reg_8_inst : DFF_X1 port map( D => n353, CK => clk, Q => a_mod_8_port,
                           QN => net108670);
   a_mod_reg_9_inst : DFF_X1 port map( D => n352, CK => clk, Q => a_mod_9_port,
                           QN => net108669);
   a_mod_reg_10_inst : DFF_X1 port map( D => n351, CK => clk, Q => 
                           a_mod_10_port, QN => net108668);
   a_mod_reg_11_inst : DFF_X1 port map( D => n350, CK => clk, Q => 
                           a_mod_11_port, QN => net108667);
   a_mod_reg_12_inst : DFF_X1 port map( D => n349, CK => clk, Q => 
                           a_mod_12_port, QN => net108666);
   a_mod_reg_13_inst : DFF_X1 port map( D => n348, CK => clk, Q => 
                           a_mod_13_port, QN => net108665);
   a_mod_reg_14_inst : DFF_X1 port map( D => n347, CK => clk, Q => 
                           a_mod_14_port, QN => net108664);
   a_mod_reg_15_inst : DFF_X1 port map( D => n346, CK => clk, Q => 
                           a_mod_15_port, QN => net108663);
   a_mod_reg_16_inst : DFF_X1 port map( D => n345, CK => clk, Q => 
                           a_mod_16_port, QN => net108662);
   a_mod_reg_17_inst : DFF_X1 port map( D => n344, CK => clk, Q => 
                           a_mod_17_port, QN => net108661);
   a_mod_reg_18_inst : DFF_X1 port map( D => n343, CK => clk, Q => 
                           a_mod_18_port, QN => net108660);
   a_mod_reg_19_inst : DFF_X1 port map( D => n342, CK => clk, Q => 
                           a_mod_19_port, QN => net108659);
   a_mod_reg_20_inst : DFF_X1 port map( D => n341, CK => clk, Q => 
                           a_mod_20_port, QN => net108658);
   a_mod_reg_21_inst : DFF_X1 port map( D => n340, CK => clk, Q => 
                           a_mod_21_port, QN => net108657);
   a_mod_reg_22_inst : DFF_X1 port map( D => n339, CK => clk, Q => 
                           a_mod_22_port, QN => net108656);
   a_mod_reg_23_inst : DFF_X1 port map( D => n338, CK => clk, Q => 
                           a_mod_23_port, QN => net108655);
   a_mod_reg_24_inst : DFF_X1 port map( D => n337, CK => clk, Q => 
                           a_mod_24_port, QN => net108654);
   a_mod_reg_25_inst : DFF_X1 port map( D => n336, CK => clk, Q => 
                           a_mod_25_port, QN => net108653);
   a_mod_reg_26_inst : DFF_X1 port map( D => n335, CK => clk, Q => 
                           a_mod_26_port, QN => net108652);
   a_mod_reg_27_inst : DFF_X1 port map( D => n334, CK => clk, Q => 
                           a_mod_27_port, QN => net108651);
   a_mod_reg_28_inst : DFF_X1 port map( D => n333, CK => clk, Q => 
                           a_mod_28_port, QN => net108650);
   a_mod_reg_29_inst : DFF_X1 port map( D => n332, CK => clk, Q => 
                           a_mod_29_port, QN => net108649);
   a_mod_reg_30_inst : DFF_X1 port map( D => n331, CK => clk, Q => 
                           a_mod_30_port, QN => net108648);
   a_mod_reg_31_inst : DFF_X1 port map( D => n330, CK => clk, Q => 
                           a_mod_31_port, QN => net108647);
   b_mod_reg_32_inst : DFF_X1 port map( D => n329, CK => clk, Q => n31_port, QN
                           => n71);
   b_mod_reg_33_inst : DFF_X1 port map( D => n328, CK => clk, Q => n70, QN => 
                           net108646);
   b_mod_reg_34_inst : DFF_X1 port map( D => n327, CK => clk, Q => n30_port, QN
                           => net108645);
   b_mod_reg_35_inst : DFF_X1 port map( D => n326, CK => clk, Q => n29_port, QN
                           => net108644);
   b_mod_reg_36_inst : DFF_X1 port map( D => n325, CK => clk, Q => n28_port, QN
                           => net108643);
   b_mod_reg_37_inst : DFF_X1 port map( D => n324, CK => clk, Q => n27_port, QN
                           => net108642);
   b_mod_reg_38_inst : DFF_X1 port map( D => n323, CK => clk, Q => n26_port, QN
                           => net108641);
   b_mod_reg_39_inst : DFF_X1 port map( D => n322, CK => clk, Q => n25_port, QN
                           => net108640);
   b_mod_reg_40_inst : DFF_X1 port map( D => n321, CK => clk, Q => n24_port, QN
                           => net108639);
   b_mod_reg_41_inst : DFF_X1 port map( D => n320, CK => clk, Q => n23_port, QN
                           => net108638);
   b_mod_reg_42_inst : DFF_X1 port map( D => n319, CK => clk, Q => n22_port, QN
                           => net108637);
   b_mod_reg_43_inst : DFF_X1 port map( D => n318, CK => clk, Q => n21_port, QN
                           => net108636);
   b_mod_reg_44_inst : DFF_X1 port map( D => n317, CK => clk, Q => n20_port, QN
                           => net108635);
   b_mod_reg_45_inst : DFF_X1 port map( D => n316, CK => clk, Q => n19_port, QN
                           => net108634);
   b_mod_reg_46_inst : DFF_X1 port map( D => n315, CK => clk, Q => n18_port, QN
                           => net108633);
   b_mod_reg_47_inst : DFF_X1 port map( D => n314, CK => clk, Q => n17_port, QN
                           => net108632);
   b_mod_reg_48_inst : DFF_X1 port map( D => n313, CK => clk, Q => n16, QN => 
                           net108631);
   b_mod_reg_49_inst : DFF_X1 port map( D => n312, CK => clk, Q => n15, QN => 
                           net108630);
   b_mod_reg_50_inst : DFF_X1 port map( D => n311, CK => clk, Q => n14, QN => 
                           net108629);
   b_mod_reg_51_inst : DFF_X1 port map( D => n310, CK => clk, Q => n13, QN => 
                           net108628);
   b_mod_reg_52_inst : DFF_X1 port map( D => n309, CK => clk, Q => n12, QN => 
                           net108627);
   b_mod_reg_53_inst : DFF_X1 port map( D => n308, CK => clk, Q => n11, QN => 
                           net108626);
   b_mod_reg_54_inst : DFF_X1 port map( D => n307, CK => clk, Q => n10, QN => 
                           net108625);
   b_mod_reg_55_inst : DFF_X1 port map( D => n306, CK => clk, Q => n9, QN => 
                           net108624);
   b_mod_reg_56_inst : DFF_X1 port map( D => n305, CK => clk, Q => n8, QN => 
                           net108623);
   b_mod_reg_57_inst : DFF_X1 port map( D => n304, CK => clk, Q => n7, QN => 
                           net108622);
   b_mod_reg_58_inst : DFF_X1 port map( D => n303, CK => clk, Q => n6, QN => 
                           net108621);
   b_mod_reg_59_inst : DFF_X1 port map( D => n302, CK => clk, Q => n5, QN => 
                           net108620);
   b_mod_reg_60_inst : DFF_X1 port map( D => n301, CK => clk, Q => n4, QN => 
                           net108619);
   b_mod_reg_61_inst : DFF_X1 port map( D => n300, CK => clk, Q => n3, QN => 
                           net108618);
   b_mod_reg_62_inst : DFF_X1 port map( D => n299, CK => clk, Q => n2, QN => 
                           net108617);
   b_mod_reg_63_inst : DFF_X1 port map( D => n298, CK => clk, Q => n1, QN => 
                           net108616);
   b_shf_31_port <= '0';
   b_shf_30_port <= '0';
   b_shf_29_port <= '0';
   b_shf_28_port <= '0';
   b_shf_27_port <= '0';
   b_shf_26_port <= '0';
   b_shf_25_port <= '0';
   b_shf_24_port <= '0';
   b_shf_23_port <= '0';
   b_shf_22_port <= '0';
   b_shf_21_port <= '0';
   b_shf_20_port <= '0';
   b_shf_19_port <= '0';
   b_shf_18_port <= '0';
   b_shf_17_port <= '0';
   b_shf_16_port <= '0';
   b_shf_15_port <= '0';
   b_shf_14_port <= '0';
   b_shf_13_port <= '0';
   b_shf_12_port <= '0';
   b_shf_11_port <= '0';
   b_shf_10_port <= '0';
   b_shf_9_port <= '0';
   b_shf_8_port <= '0';
   b_shf_7_port <= '0';
   b_shf_6_port <= '0';
   b_shf_5_port <= '0';
   b_shf_4_port <= '0';
   b_shf_3_port <= '0';
   b_shf_2_port <= '0';
   b_shf_1_port <= '0';
   b_shf_0_port <= '0';
   a_mod_63_port <= '0';
   a_mod_62_port <= '0';
   a_mod_61_port <= '0';
   a_mod_60_port <= '0';
   a_mod_59_port <= '0';
   a_mod_58_port <= '0';
   a_mod_57_port <= '0';
   a_mod_56_port <= '0';
   a_mod_55_port <= '0';
   a_mod_54_port <= '0';
   a_mod_53_port <= '0';
   a_mod_52_port <= '0';
   a_mod_51_port <= '0';
   a_mod_50_port <= '0';
   a_mod_49_port <= '0';
   a_mod_48_port <= '0';
   a_mod_47_port <= '0';
   a_mod_46_port <= '0';
   a_mod_45_port <= '0';
   a_mod_44_port <= '0';
   a_mod_43_port <= '0';
   a_mod_42_port <= '0';
   a_mod_41_port <= '0';
   a_mod_40_port <= '0';
   a_mod_39_port <= '0';
   a_mod_38_port <= '0';
   a_mod_37_port <= '0';
   a_mod_36_port <= '0';
   a_mod_35_port <= '0';
   a_mod_34_port <= '0';
   a_mod_33_port <= '0';
   a_mod_32_port <= '0';
   ADJUST0a : AddSub_DATA_SIZE32_0 port map( as => inv_a_flag, a(31) => 
                           X_Logic0_port, a(30) => X_Logic0_port, a(29) => 
                           X_Logic0_port, a(28) => X_Logic0_port, a(27) => 
                           X_Logic0_port, a(26) => X_Logic0_port, a(25) => 
                           X_Logic0_port, a(24) => X_Logic0_port, a(23) => 
                           X_Logic0_port, a(22) => X_Logic0_port, a(21) => 
                           X_Logic0_port, a(20) => X_Logic0_port, a(19) => 
                           X_Logic0_port, a(18) => X_Logic0_port, a(17) => 
                           X_Logic0_port, a(16) => X_Logic0_port, a(15) => 
                           X_Logic0_port, a(14) => X_Logic0_port, a(13) => 
                           X_Logic0_port, a(12) => X_Logic0_port, a(11) => 
                           X_Logic0_port, a(10) => X_Logic0_port, a(9) => 
                           X_Logic0_port, a(8) => X_Logic0_port, a(7) => 
                           X_Logic0_port, a(6) => X_Logic0_port, a(5) => 
                           X_Logic0_port, a(4) => X_Logic0_port, a(3) => 
                           X_Logic0_port, a(2) => X_Logic0_port, a(1) => 
                           X_Logic0_port, a(0) => X_Logic0_port, b(31) => a(31)
                           , b(30) => a(30), b(29) => a(29), b(28) => a(28), 
                           b(27) => a(27), b(26) => a(26), b(25) => a(25), 
                           b(24) => a(24), b(23) => a(23), b(22) => a(22), 
                           b(21) => a(21), b(20) => a(20), b(19) => a(19), 
                           b(18) => a(18), b(17) => a(17), b(16) => a(16), 
                           b(15) => a(15), b(14) => a(14), b(13) => a(13), 
                           b(12) => a(12), b(11) => a(11), b(10) => a(10), b(9)
                           => a(9), b(8) => a(8), b(7) => a(7), b(6) => a(6), 
                           b(5) => a(5), b(4) => a(4), b(3) => a(3), b(2) => 
                           a(2), b(1) => a(1), b(0) => a(0), re(31) => 
                           a_adj_31_port, re(30) => a_adj_30_port, re(29) => 
                           a_adj_29_port, re(28) => a_adj_28_port, re(27) => 
                           a_adj_27_port, re(26) => a_adj_26_port, re(25) => 
                           a_adj_25_port, re(24) => a_adj_24_port, re(23) => 
                           a_adj_23_port, re(22) => a_adj_22_port, re(21) => 
                           a_adj_21_port, re(20) => a_adj_20_port, re(19) => 
                           a_adj_19_port, re(18) => a_adj_18_port, re(17) => 
                           a_adj_17_port, re(16) => a_adj_16_port, re(15) => 
                           a_adj_15_port, re(14) => a_adj_14_port, re(13) => 
                           a_adj_13_port, re(12) => a_adj_12_port, re(11) => 
                           a_adj_11_port, re(10) => a_adj_10_port, re(9) => 
                           a_adj_9_port, re(8) => a_adj_8_port, re(7) => 
                           a_adj_7_port, re(6) => a_adj_6_port, re(5) => 
                           a_adj_5_port, re(4) => a_adj_4_port, re(3) => 
                           a_adj_3_port, re(2) => a_adj_2_port, re(1) => 
                           a_adj_1_port, re(0) => a_adj_0_port, cout => net3930
                           );
   ADJUST0b : AddSub_DATA_SIZE32_3 port map( as => inv_b_flag, a(31) => 
                           X_Logic0_port, a(30) => X_Logic0_port, a(29) => 
                           X_Logic0_port, a(28) => X_Logic0_port, a(27) => 
                           X_Logic0_port, a(26) => X_Logic0_port, a(25) => 
                           X_Logic0_port, a(24) => X_Logic0_port, a(23) => 
                           X_Logic0_port, a(22) => X_Logic0_port, a(21) => 
                           X_Logic0_port, a(20) => X_Logic0_port, a(19) => 
                           X_Logic0_port, a(18) => X_Logic0_port, a(17) => 
                           X_Logic0_port, a(16) => X_Logic0_port, a(15) => 
                           X_Logic0_port, a(14) => X_Logic0_port, a(13) => 
                           X_Logic0_port, a(12) => X_Logic0_port, a(11) => 
                           X_Logic0_port, a(10) => X_Logic0_port, a(9) => 
                           X_Logic0_port, a(8) => X_Logic0_port, a(7) => 
                           X_Logic0_port, a(6) => X_Logic0_port, a(5) => 
                           X_Logic0_port, a(4) => X_Logic0_port, a(3) => 
                           X_Logic0_port, a(2) => X_Logic0_port, a(1) => 
                           X_Logic0_port, a(0) => X_Logic0_port, b(31) => b(31)
                           , b(30) => b(30), b(29) => b(29), b(28) => b(28), 
                           b(27) => b(27), b(26) => b(26), b(25) => b(25), 
                           b(24) => b(24), b(23) => b(23), b(22) => b(22), 
                           b(21) => b(21), b(20) => b(20), b(19) => b(19), 
                           b(18) => b(18), b(17) => b(17), b(16) => b(16), 
                           b(15) => b(15), b(14) => b(14), b(13) => b(13), 
                           b(12) => b(12), b(11) => b(11), b(10) => b(10), b(9)
                           => b(9), b(8) => b(8), b(7) => b(7), b(6) => b(6), 
                           b(5) => b(5), b(4) => b(4), b(3) => b(3), b(2) => 
                           b(2), b(1) => b(1), b(0) => b(0), re(31) => 
                           b_adj_31_port, re(30) => b_adj_30_port, re(29) => 
                           b_adj_29_port, re(28) => b_adj_28_port, re(27) => 
                           b_adj_27_port, re(26) => b_adj_26_port, re(25) => 
                           b_adj_25_port, re(24) => b_adj_24_port, re(23) => 
                           b_adj_23_port, re(22) => b_adj_22_port, re(21) => 
                           b_adj_21_port, re(20) => b_adj_20_port, re(19) => 
                           b_adj_19_port, re(18) => b_adj_18_port, re(17) => 
                           b_adj_17_port, re(16) => b_adj_16_port, re(15) => 
                           b_adj_15_port, re(14) => b_adj_14_port, re(13) => 
                           b_adj_13_port, re(12) => b_adj_12_port, re(11) => 
                           b_adj_11_port, re(10) => b_adj_10_port, re(9) => 
                           b_adj_9_port, re(8) => b_adj_8_port, re(7) => 
                           b_adj_7_port, re(6) => b_adj_6_port, re(5) => 
                           b_adj_5_port, re(4) => b_adj_4_port, re(3) => 
                           b_adj_3_port, re(2) => b_adj_2_port, re(1) => 
                           b_adj_1_port, re(0) => b_adj_0_port, cout => net3929
                           );
   MUXa : Mux_DATA_SIZE64 port map( sel => n37_port, din0(63) => a_mod_63_port,
                           din0(62) => a_mod_62_port, din0(61) => a_mod_61_port
                           , din0(60) => a_mod_60_port, din0(59) => 
                           a_mod_59_port, din0(58) => a_mod_58_port, din0(57) 
                           => a_mod_57_port, din0(56) => a_mod_56_port, 
                           din0(55) => a_mod_55_port, din0(54) => a_mod_54_port
                           , din0(53) => a_mod_53_port, din0(52) => 
                           a_mod_52_port, din0(51) => a_mod_51_port, din0(50) 
                           => a_mod_50_port, din0(49) => a_mod_49_port, 
                           din0(48) => a_mod_48_port, din0(47) => a_mod_47_port
                           , din0(46) => a_mod_46_port, din0(45) => 
                           a_mod_45_port, din0(44) => a_mod_44_port, din0(43) 
                           => a_mod_43_port, din0(42) => a_mod_42_port, 
                           din0(41) => a_mod_41_port, din0(40) => a_mod_40_port
                           , din0(39) => a_mod_39_port, din0(38) => 
                           a_mod_38_port, din0(37) => a_mod_37_port, din0(36) 
                           => a_mod_36_port, din0(35) => a_mod_35_port, 
                           din0(34) => a_mod_34_port, din0(33) => a_mod_33_port
                           , din0(32) => a_mod_32_port, din0(31) => 
                           a_mod_31_port, din0(30) => a_mod_30_port, din0(29) 
                           => a_mod_29_port, din0(28) => a_mod_28_port, 
                           din0(27) => a_mod_27_port, din0(26) => a_mod_26_port
                           , din0(25) => a_mod_25_port, din0(24) => 
                           a_mod_24_port, din0(23) => a_mod_23_port, din0(22) 
                           => a_mod_22_port, din0(21) => a_mod_21_port, 
                           din0(20) => a_mod_20_port, din0(19) => a_mod_19_port
                           , din0(18) => a_mod_18_port, din0(17) => 
                           a_mod_17_port, din0(16) => a_mod_16_port, din0(15) 
                           => a_mod_15_port, din0(14) => a_mod_14_port, 
                           din0(13) => a_mod_13_port, din0(12) => a_mod_12_port
                           , din0(11) => a_mod_11_port, din0(10) => 
                           a_mod_10_port, din0(9) => a_mod_9_port, din0(8) => 
                           a_mod_8_port, din0(7) => a_mod_7_port, din0(6) => 
                           a_mod_6_port, din0(5) => a_mod_5_port, din0(4) => 
                           a_mod_4_port, din0(3) => a_mod_3_port, din0(2) => 
                           a_mod_2_port, din0(1) => a_mod_1_port, din0(0) => 
                           a_mod_0_port, din1(63) => r_63_port, din1(62) => 
                           r_62_port, din1(61) => r_61_port, din1(60) => 
                           r_60_port, din1(59) => r_59_port, din1(58) => 
                           r_58_port, din1(57) => r_57_port, din1(56) => 
                           r_56_port, din1(55) => r_55_port, din1(54) => 
                           r_54_port, din1(53) => r_53_port, din1(52) => 
                           r_52_port, din1(51) => r_51_port, din1(50) => 
                           r_50_port, din1(49) => r_49_port, din1(48) => 
                           r_48_port, din1(47) => r_47_port, din1(46) => 
                           r_46_port, din1(45) => r_45_port, din1(44) => 
                           r_44_port, din1(43) => r_43_port, din1(42) => 
                           r_42_port, din1(41) => r_41_port, din1(40) => 
                           r_40_port, din1(39) => r_39_port, din1(38) => 
                           r_38_port, din1(37) => r_37_port, din1(36) => 
                           r_36_port, din1(35) => r_35_port, din1(34) => 
                           r_34_port, din1(33) => r_33_port, din1(32) => 
                           r_32_port, din1(31) => r_31_port, din1(30) => 
                           r_30_port, din1(29) => r_29_port, din1(28) => 
                           r_28_port, din1(27) => r_27_port, din1(26) => 
                           r_26_port, din1(25) => r_25_port, din1(24) => 
                           r_24_port, din1(23) => r_23_port, din1(22) => 
                           r_22_port, din1(21) => r_21_port, din1(20) => 
                           r_20_port, din1(19) => r_19_port, din1(18) => 
                           r_18_port, din1(17) => r_17_port, din1(16) => 
                           r_16_port, din1(15) => r_15_port, din1(14) => 
                           r_14_port, din1(13) => r_13_port, din1(12) => 
                           r_12_port, din1(11) => r_11_port, din1(10) => 
                           r_10_port, din1(9) => r_9_port, din1(8) => r_8_port,
                           din1(7) => r_7_port, din1(6) => r_6_port, din1(5) =>
                           r_5_port, din1(4) => r_4_port, din1(3) => r_3_port, 
                           din1(2) => r_2_port, din1(1) => r_1_port, din1(0) =>
                           r_0_port, dout(63) => a_mux_63_port, dout(62) => 
                           a_mux_62_port, dout(61) => a_mux_61_port, dout(60) 
                           => a_mux_60_port, dout(59) => a_mux_59_port, 
                           dout(58) => a_mux_58_port, dout(57) => a_mux_57_port
                           , dout(56) => a_mux_56_port, dout(55) => 
                           a_mux_55_port, dout(54) => a_mux_54_port, dout(53) 
                           => a_mux_53_port, dout(52) => a_mux_52_port, 
                           dout(51) => a_mux_51_port, dout(50) => a_mux_50_port
                           , dout(49) => a_mux_49_port, dout(48) => 
                           a_mux_48_port, dout(47) => a_mux_47_port, dout(46) 
                           => a_mux_46_port, dout(45) => a_mux_45_port, 
                           dout(44) => a_mux_44_port, dout(43) => a_mux_43_port
                           , dout(42) => a_mux_42_port, dout(41) => 
                           a_mux_41_port, dout(40) => a_mux_40_port, dout(39) 
                           => a_mux_39_port, dout(38) => a_mux_38_port, 
                           dout(37) => a_mux_37_port, dout(36) => a_mux_36_port
                           , dout(35) => a_mux_35_port, dout(34) => 
                           a_mux_34_port, dout(33) => a_mux_33_port, dout(32) 
                           => a_mux_32_port, dout(31) => a_mux_31_port, 
                           dout(30) => a_mux_30_port, dout(29) => a_mux_29_port
                           , dout(28) => a_mux_28_port, dout(27) => 
                           a_mux_27_port, dout(26) => a_mux_26_port, dout(25) 
                           => a_mux_25_port, dout(24) => a_mux_24_port, 
                           dout(23) => a_mux_23_port, dout(22) => a_mux_22_port
                           , dout(21) => a_mux_21_port, dout(20) => 
                           a_mux_20_port, dout(19) => a_mux_19_port, dout(18) 
                           => a_mux_18_port, dout(17) => a_mux_17_port, 
                           dout(16) => a_mux_16_port, dout(15) => a_mux_15_port
                           , dout(14) => a_mux_14_port, dout(13) => 
                           a_mux_13_port, dout(12) => a_mux_12_port, dout(11) 
                           => a_mux_11_port, dout(10) => a_mux_10_port, dout(9)
                           => a_mux_9_port, dout(8) => a_mux_8_port, dout(7) =>
                           a_mux_7_port, dout(6) => a_mux_6_port, dout(5) => 
                           a_mux_5_port, dout(4) => a_mux_4_port, dout(3) => 
                           a_mux_3_port, dout(2) => a_mux_2_port, dout(1) => 
                           a_mux_1_port, dout(0) => a_mux_0_port);
   ADD0 : AddSub_DATA_SIZE64 port map( as => not_r_sign, a(63) => a_shf_63_port
                           , a(62) => a_shf_62_port, a(61) => a_shf_61_port, 
                           a(60) => a_shf_60_port, a(59) => a_shf_59_port, 
                           a(58) => a_shf_58_port, a(57) => a_shf_57_port, 
                           a(56) => a_shf_56_port, a(55) => a_shf_55_port, 
                           a(54) => a_shf_54_port, a(53) => a_shf_53_port, 
                           a(52) => a_shf_52_port, a(51) => a_shf_51_port, 
                           a(50) => a_shf_50_port, a(49) => a_shf_49_port, 
                           a(48) => a_shf_48_port, a(47) => a_shf_47_port, 
                           a(46) => a_shf_46_port, a(45) => a_shf_45_port, 
                           a(44) => a_shf_44_port, a(43) => a_shf_43_port, 
                           a(42) => a_shf_42_port, a(41) => a_shf_41_port, 
                           a(40) => a_shf_40_port, a(39) => a_shf_39_port, 
                           a(38) => a_shf_38_port, a(37) => a_shf_37_port, 
                           a(36) => a_shf_36_port, a(35) => a_shf_35_port, 
                           a(34) => a_shf_34_port, a(33) => a_shf_33_port, 
                           a(32) => a_shf_32_port, a(31) => a_shf_31_port, 
                           a(30) => a_shf_30_port, a(29) => a_shf_29_port, 
                           a(28) => a_shf_28_port, a(27) => a_shf_27_port, 
                           a(26) => a_shf_26_port, a(25) => a_shf_25_port, 
                           a(24) => a_shf_24_port, a(23) => a_shf_23_port, 
                           a(22) => a_shf_22_port, a(21) => a_shf_21_port, 
                           a(20) => a_shf_20_port, a(19) => a_shf_19_port, 
                           a(18) => a_shf_18_port, a(17) => a_shf_17_port, 
                           a(16) => a_shf_16_port, a(15) => a_shf_15_port, 
                           a(14) => a_shf_14_port, a(13) => a_shf_13_port, 
                           a(12) => a_shf_12_port, a(11) => a_shf_11_port, 
                           a(10) => a_shf_10_port, a(9) => a_shf_9_port, a(8) 
                           => a_shf_8_port, a(7) => a_shf_7_port, a(6) => 
                           a_shf_6_port, a(5) => a_shf_5_port, a(4) => 
                           a_shf_4_port, a(3) => a_shf_3_port, a(2) => 
                           a_shf_2_port, a(1) => a_shf_1_port, a(0) => 
                           X_Logic0_port, b(63) => b_shf_63_port, b(62) => 
                           b_shf_62_port, b(61) => b_shf_61_port, b(60) => 
                           b_shf_60_port, b(59) => b_shf_59_port, b(58) => 
                           b_shf_58_port, b(57) => b_shf_57_port, b(56) => 
                           b_shf_56_port, b(55) => b_shf_55_port, b(54) => 
                           b_shf_54_port, b(53) => b_shf_53_port, b(52) => 
                           b_shf_52_port, b(51) => b_shf_51_port, b(50) => 
                           b_shf_50_port, b(49) => b_shf_49_port, b(48) => 
                           b_shf_48_port, b(47) => b_shf_47_port, b(46) => 
                           b_shf_46_port, b(45) => b_shf_45_port, b(44) => 
                           b_shf_44_port, b(43) => b_shf_43_port, b(42) => 
                           b_shf_42_port, b(41) => b_shf_41_port, b(40) => 
                           b_shf_40_port, b(39) => b_shf_39_port, b(38) => 
                           b_shf_38_port, b(37) => b_shf_37_port, b(36) => 
                           b_shf_36_port, b(35) => b_shf_35_port, b(34) => 
                           b_shf_34_port, b(33) => b_shf_33_port, b(32) => 
                           b_shf_32_port, b(31) => b_shf_31_port, b(30) => 
                           b_shf_30_port, b(29) => b_shf_29_port, b(28) => 
                           b_shf_28_port, b(27) => b_shf_27_port, b(26) => 
                           b_shf_26_port, b(25) => b_shf_25_port, b(24) => 
                           b_shf_24_port, b(23) => b_shf_23_port, b(22) => 
                           b_shf_22_port, b(21) => b_shf_21_port, b(20) => 
                           b_shf_20_port, b(19) => b_shf_19_port, b(18) => 
                           b_shf_18_port, b(17) => b_shf_17_port, b(16) => 
                           b_shf_16_port, b(15) => b_shf_15_port, b(14) => 
                           b_shf_14_port, b(13) => b_shf_13_port, b(12) => 
                           b_shf_12_port, b(11) => b_shf_11_port, b(10) => 
                           b_shf_10_port, b(9) => b_shf_9_port, b(8) => 
                           b_shf_8_port, b(7) => b_shf_7_port, b(6) => 
                           b_shf_6_port, b(5) => b_shf_5_port, b(4) => 
                           b_shf_4_port, b(3) => b_shf_3_port, b(2) => 
                           b_shf_2_port, b(1) => b_shf_1_port, b(0) => 
                           b_shf_0_port, re(63) => r_es_63_port, re(62) => 
                           r_es_62_port, re(61) => r_es_61_port, re(60) => 
                           r_es_60_port, re(59) => r_es_59_port, re(58) => 
                           r_es_58_port, re(57) => r_es_57_port, re(56) => 
                           r_es_56_port, re(55) => r_es_55_port, re(54) => 
                           r_es_54_port, re(53) => r_es_53_port, re(52) => 
                           r_es_52_port, re(51) => r_es_51_port, re(50) => 
                           r_es_50_port, re(49) => r_es_49_port, re(48) => 
                           r_es_48_port, re(47) => r_es_47_port, re(46) => 
                           r_es_46_port, re(45) => r_es_45_port, re(44) => 
                           r_es_44_port, re(43) => r_es_43_port, re(42) => 
                           r_es_42_port, re(41) => r_es_41_port, re(40) => 
                           r_es_40_port, re(39) => r_es_39_port, re(38) => 
                           r_es_38_port, re(37) => r_es_37_port, re(36) => 
                           r_es_36_port, re(35) => r_es_35_port, re(34) => 
                           r_es_34_port, re(33) => r_es_33_port, re(32) => 
                           r_es_32_port, re(31) => r_es_31_port, re(30) => 
                           r_es_30_port, re(29) => r_es_29_port, re(28) => 
                           r_es_28_port, re(27) => r_es_27_port, re(26) => 
                           r_es_26_port, re(25) => r_es_25_port, re(24) => 
                           r_es_24_port, re(23) => r_es_23_port, re(22) => 
                           r_es_22_port, re(21) => r_es_21_port, re(20) => 
                           r_es_20_port, re(19) => r_es_19_port, re(18) => 
                           r_es_18_port, re(17) => r_es_17_port, re(16) => 
                           r_es_16_port, re(15) => r_es_15_port, re(14) => 
                           r_es_14_port, re(13) => r_es_13_port, re(12) => 
                           r_es_12_port, re(11) => r_es_11_port, re(10) => 
                           r_es_10_port, re(9) => r_es_9_port, re(8) => 
                           r_es_8_port, re(7) => r_es_7_port, re(6) => 
                           r_es_6_port, re(5) => r_es_5_port, re(4) => 
                           r_es_4_port, re(3) => r_es_3_port, re(2) => 
                           r_es_2_port, re(1) => r_es_1_port, re(0) => 
                           r_es_0_port, cout => net3928);
   REG_R : Reg_DATA_SIZE64 port map( rst => n33_port, en => n38_port, clk => 
                           clk, din(63) => r_es_63_port, din(62) => 
                           r_es_62_port, din(61) => r_es_61_port, din(60) => 
                           r_es_60_port, din(59) => r_es_59_port, din(58) => 
                           r_es_58_port, din(57) => r_es_57_port, din(56) => 
                           r_es_56_port, din(55) => r_es_55_port, din(54) => 
                           r_es_54_port, din(53) => r_es_53_port, din(52) => 
                           r_es_52_port, din(51) => r_es_51_port, din(50) => 
                           r_es_50_port, din(49) => r_es_49_port, din(48) => 
                           r_es_48_port, din(47) => r_es_47_port, din(46) => 
                           r_es_46_port, din(45) => r_es_45_port, din(44) => 
                           r_es_44_port, din(43) => r_es_43_port, din(42) => 
                           r_es_42_port, din(41) => r_es_41_port, din(40) => 
                           r_es_40_port, din(39) => r_es_39_port, din(38) => 
                           r_es_38_port, din(37) => r_es_37_port, din(36) => 
                           r_es_36_port, din(35) => r_es_35_port, din(34) => 
                           r_es_34_port, din(33) => r_es_33_port, din(32) => 
                           r_es_32_port, din(31) => r_es_31_port, din(30) => 
                           r_es_30_port, din(29) => r_es_29_port, din(28) => 
                           r_es_28_port, din(27) => r_es_27_port, din(26) => 
                           r_es_26_port, din(25) => r_es_25_port, din(24) => 
                           r_es_24_port, din(23) => r_es_23_port, din(22) => 
                           r_es_22_port, din(21) => r_es_21_port, din(20) => 
                           r_es_20_port, din(19) => r_es_19_port, din(18) => 
                           r_es_18_port, din(17) => r_es_17_port, din(16) => 
                           r_es_16_port, din(15) => r_es_15_port, din(14) => 
                           r_es_14_port, din(13) => r_es_13_port, din(12) => 
                           r_es_12_port, din(11) => r_es_11_port, din(10) => 
                           r_es_10_port, din(9) => r_es_9_port, din(8) => 
                           r_es_8_port, din(7) => r_es_7_port, din(6) => 
                           r_es_6_port, din(5) => r_es_5_port, din(4) => 
                           r_es_4_port, din(3) => r_es_3_port, din(2) => 
                           r_es_2_port, din(1) => r_es_1_port, din(0) => 
                           r_es_0_port, dout(63) => r_63_port, dout(62) => 
                           r_62_port, dout(61) => r_61_port, dout(60) => 
                           r_60_port, dout(59) => r_59_port, dout(58) => 
                           r_58_port, dout(57) => r_57_port, dout(56) => 
                           r_56_port, dout(55) => r_55_port, dout(54) => 
                           r_54_port, dout(53) => r_53_port, dout(52) => 
                           r_52_port, dout(51) => r_51_port, dout(50) => 
                           r_50_port, dout(49) => r_49_port, dout(48) => 
                           r_48_port, dout(47) => r_47_port, dout(46) => 
                           r_46_port, dout(45) => r_45_port, dout(44) => 
                           r_44_port, dout(43) => r_43_port, dout(42) => 
                           r_42_port, dout(41) => r_41_port, dout(40) => 
                           r_40_port, dout(39) => r_39_port, dout(38) => 
                           r_38_port, dout(37) => r_37_port, dout(36) => 
                           r_36_port, dout(35) => r_35_port, dout(34) => 
                           r_34_port, dout(33) => r_33_port, dout(32) => 
                           r_32_port, dout(31) => r_31_port, dout(30) => 
                           r_30_port, dout(29) => r_29_port, dout(28) => 
                           r_28_port, dout(27) => r_27_port, dout(26) => 
                           r_26_port, dout(25) => r_25_port, dout(24) => 
                           r_24_port, dout(23) => r_23_port, dout(22) => 
                           r_22_port, dout(21) => r_21_port, dout(20) => 
                           r_20_port, dout(19) => r_19_port, dout(18) => 
                           r_18_port, dout(17) => r_17_port, dout(16) => 
                           r_16_port, dout(15) => r_15_port, dout(14) => 
                           r_14_port, dout(13) => r_13_port, dout(12) => 
                           r_12_port, dout(11) => r_11_port, dout(10) => 
                           r_10_port, dout(9) => r_9_port, dout(8) => r_8_port,
                           dout(7) => r_7_port, dout(6) => r_6_port, dout(5) =>
                           r_5_port, dout(4) => r_4_port, dout(3) => r_3_port, 
                           dout(2) => r_2_port, dout(1) => r_1_port, dout(0) =>
                           r_0_port);
   REG_Q : Sipo_DATA_SIZE32 port map( rst => n34_port, en => n38_port, clk => 
                           clk, din => not_r_es_sign, dout(31) => q_31_port, 
                           dout(30) => q_30_port, dout(29) => 
                           b_shf_sqrt_63_port, dout(28) => b_shf_sqrt_62_port, 
                           dout(27) => b_shf_sqrt_61_port, dout(26) => 
                           b_shf_sqrt_60_port, dout(25) => b_shf_sqrt_59_port, 
                           dout(24) => b_shf_sqrt_58_port, dout(23) => 
                           b_shf_sqrt_57_port, dout(22) => b_shf_sqrt_56_port, 
                           dout(21) => b_shf_sqrt_55_port, dout(20) => 
                           b_shf_sqrt_54_port, dout(19) => b_shf_sqrt_53_port, 
                           dout(18) => b_shf_sqrt_52_port, dout(17) => 
                           b_shf_sqrt_51_port, dout(16) => b_shf_sqrt_50_port, 
                           dout(15) => b_shf_sqrt_49_port, dout(14) => 
                           b_shf_sqrt_48_port, dout(13) => b_shf_sqrt_47_port, 
                           dout(12) => b_shf_sqrt_46_port, dout(11) => 
                           b_shf_sqrt_45_port, dout(10) => b_shf_sqrt_44_port, 
                           dout(9) => b_shf_sqrt_43_port, dout(8) => 
                           b_shf_sqrt_42_port, dout(7) => b_shf_sqrt_41_port, 
                           dout(6) => b_shf_sqrt_40_port, dout(5) => 
                           b_shf_sqrt_39_port, dout(4) => b_shf_sqrt_38_port, 
                           dout(3) => b_shf_sqrt_37_port, dout(2) => 
                           b_shf_sqrt_36_port, dout(1) => b_shf_sqrt_35_port, 
                           dout(0) => b_shf_sqrt_34_port);
   ADJUST : AddSub_DATA_SIZE32_2 port map( as => inv_q_flag_mod, a(31) => 
                           X_Logic0_port, a(30) => X_Logic0_port, a(29) => 
                           X_Logic0_port, a(28) => X_Logic0_port, a(27) => 
                           X_Logic0_port, a(26) => X_Logic0_port, a(25) => 
                           X_Logic0_port, a(24) => X_Logic0_port, a(23) => 
                           X_Logic0_port, a(22) => X_Logic0_port, a(21) => 
                           X_Logic0_port, a(20) => X_Logic0_port, a(19) => 
                           X_Logic0_port, a(18) => X_Logic0_port, a(17) => 
                           X_Logic0_port, a(16) => X_Logic0_port, a(15) => 
                           X_Logic0_port, a(14) => X_Logic0_port, a(13) => 
                           X_Logic0_port, a(12) => X_Logic0_port, a(11) => 
                           X_Logic0_port, a(10) => X_Logic0_port, a(9) => 
                           X_Logic0_port, a(8) => X_Logic0_port, a(7) => 
                           X_Logic0_port, a(6) => X_Logic0_port, a(5) => 
                           X_Logic0_port, a(4) => X_Logic0_port, a(3) => 
                           X_Logic0_port, a(2) => X_Logic0_port, a(1) => 
                           X_Logic0_port, a(0) => X_Logic0_port, b(31) => 
                           q_31_port, b(30) => q_30_port, b(29) => 
                           b_shf_sqrt_63_port, b(28) => b_shf_sqrt_62_port, 
                           b(27) => b_shf_sqrt_61_port, b(26) => 
                           b_shf_sqrt_60_port, b(25) => b_shf_sqrt_59_port, 
                           b(24) => b_shf_sqrt_58_port, b(23) => 
                           b_shf_sqrt_57_port, b(22) => b_shf_sqrt_56_port, 
                           b(21) => b_shf_sqrt_55_port, b(20) => 
                           b_shf_sqrt_54_port, b(19) => b_shf_sqrt_53_port, 
                           b(18) => b_shf_sqrt_52_port, b(17) => 
                           b_shf_sqrt_51_port, b(16) => b_shf_sqrt_50_port, 
                           b(15) => b_shf_sqrt_49_port, b(14) => 
                           b_shf_sqrt_48_port, b(13) => b_shf_sqrt_47_port, 
                           b(12) => b_shf_sqrt_46_port, b(11) => 
                           b_shf_sqrt_45_port, b(10) => b_shf_sqrt_44_port, 
                           b(9) => b_shf_sqrt_43_port, b(8) => 
                           b_shf_sqrt_42_port, b(7) => b_shf_sqrt_41_port, b(6)
                           => b_shf_sqrt_40_port, b(5) => b_shf_sqrt_39_port, 
                           b(4) => b_shf_sqrt_38_port, b(3) => 
                           b_shf_sqrt_37_port, b(2) => b_shf_sqrt_36_port, b(1)
                           => b_shf_sqrt_35_port, b(0) => b_shf_sqrt_34_port, 
                           re(31) => o(31), re(30) => o(30), re(29) => o(29), 
                           re(28) => o(28), re(27) => o(27), re(26) => o(26), 
                           re(25) => o(25), re(24) => o(24), re(23) => o(23), 
                           re(22) => o(22), re(21) => o(21), re(20) => o(20), 
                           re(19) => o(19), re(18) => o(18), re(17) => o(17), 
                           re(16) => o(16), re(15) => o(15), re(14) => o(14), 
                           re(13) => o(13), re(12) => o(12), re(11) => o(11), 
                           re(10) => o(10), re(9) => o(9), re(8) => o(8), re(7)
                           => o(7), re(6) => o(6), re(5) => o(5), re(4) => o(4)
                           , re(3) => o(3), re(2) => o(2), re(1) => o(1), re(0)
                           => o(0), cout => net3927);
   add_197 : Div_DATA_SIZE32_DIV_STAGE34_SQRT_STAGE18_DW01_inc_0 port map( 
                           A(31) => c_state_31_port, A(30) => c_state_30_port, 
                           A(29) => c_state_29_port, A(28) => c_state_28_port, 
                           A(27) => c_state_27_port, A(26) => c_state_26_port, 
                           A(25) => c_state_25_port, A(24) => c_state_24_port, 
                           A(23) => c_state_23_port, A(22) => c_state_22_port, 
                           A(21) => c_state_21_port, A(20) => c_state_20_port, 
                           A(19) => c_state_19_port, A(18) => c_state_18_port, 
                           A(17) => c_state_17_port, A(16) => c_state_16_port, 
                           A(15) => c_state_15_port, A(14) => c_state_14_port, 
                           A(13) => c_state_13_port, A(12) => c_state_12_port, 
                           A(11) => c_state_11_port, A(10) => c_state_10_port, 
                           A(9) => c_state_9_port, A(8) => c_state_8_port, A(7)
                           => c_state_7_port, A(6) => c_state_6_port, A(5) => 
                           c_state_5_port, A(4) => c_state_4_port, A(3) => 
                           c_state_3_port, A(2) => c_state_2_port, A(1) => 
                           c_state_1_port, A(0) => c_state_0_port, SUM(31) => 
                           N48, SUM(30) => N47, SUM(29) => N46, SUM(28) => N45,
                           SUM(27) => N44, SUM(26) => N43, SUM(25) => N42, 
                           SUM(24) => N41, SUM(23) => N40, SUM(22) => N39, 
                           SUM(21) => N38, SUM(20) => N37, SUM(19) => N36, 
                           SUM(18) => N35, SUM(17) => N34, SUM(16) => N33, 
                           SUM(15) => N32, SUM(14) => N31, SUM(13) => N30, 
                           SUM(12) => N29, SUM(11) => N28, SUM(10) => N27, 
                           SUM(9) => N26, SUM(8) => N25, SUM(7) => N24, SUM(6) 
                           => N23, SUM(5) => N22, SUM(4) => N21, SUM(3) => N20,
                           SUM(2) => N19, SUM(1) => N18, SUM(0) => N17);
   inv_q_flag_mod_reg : DFF_X2 port map( D => n297, CK => clk, Q => 
                           inv_q_flag_mod, QN => n35_port);
   U3 : AOI22_X4 port map( A1 => en, A2 => lock, B1 => n46_port, B2 => n72, ZN 
                           => n41_port);
   U4 : INV_X2 port map( A => n52, ZN => inv_a_flag);
   U5 : INV_X2 port map( A => n51, ZN => inv_b_flag);
   U6 : NAND2_X1 port map( A1 => rst, A2 => n40_port, ZN => n32_port);
   U7 : INV_X4 port map( A => n32_port, ZN => n33_port);
   U8 : INV_X2 port map( A => n32_port, ZN => n34_port);
   U9 : INV_X8 port map( A => func, ZN => n53);
   U10 : INV_X4 port map( A => a_mux_63_port, ZN => not_r_sign);
   U11 : OR3_X1 port map( A1 => n47_port, A2 => n45_port, A3 => c_state_31_port
                           , ZN => n36_port);
   U12 : INV_X4 port map( A => n36_port, ZN => n37_port);
   U13 : BUF_X2 port map( A => en_r, Z => n38_port);
   U14 : BUF_X2 port map( A => en_r, Z => n39_port);
   U15 : BUF_X1 port map( A => en_r, Z => n40_port);
   U16 : INV_X1 port map( A => r_es_63_port, ZN => not_r_es_sign);
   U17 : AND2_X1 port map( A1 => N26, A2 => n41_port, ZN => n_state_9_port);
   U18 : AND2_X1 port map( A1 => N25, A2 => n41_port, ZN => n_state_8_port);
   U19 : AND2_X1 port map( A1 => N24, A2 => n41_port, ZN => n_state_7_port);
   U20 : AND2_X1 port map( A1 => N23, A2 => n41_port, ZN => n_state_6_port);
   U21 : AND2_X1 port map( A1 => N22, A2 => n41_port, ZN => n_state_5_port);
   U22 : AND2_X1 port map( A1 => N21, A2 => n41_port, ZN => n_state_4_port);
   U23 : AND2_X1 port map( A1 => N20, A2 => n41_port, ZN => n_state_3_port);
   U24 : AND2_X1 port map( A1 => N48, A2 => n41_port, ZN => n_state_31_port);
   U25 : AND2_X1 port map( A1 => N47, A2 => n41_port, ZN => n_state_30_port);
   U26 : AND2_X1 port map( A1 => N19, A2 => n41_port, ZN => n_state_2_port);
   U27 : AND2_X1 port map( A1 => N46, A2 => n41_port, ZN => n_state_29_port);
   U28 : AND2_X1 port map( A1 => N45, A2 => n41_port, ZN => n_state_28_port);
   U29 : AND2_X1 port map( A1 => N44, A2 => n41_port, ZN => n_state_27_port);
   U30 : AND2_X1 port map( A1 => N43, A2 => n41_port, ZN => n_state_26_port);
   U31 : AND2_X1 port map( A1 => N42, A2 => n41_port, ZN => n_state_25_port);
   U32 : AND2_X1 port map( A1 => N41, A2 => n41_port, ZN => n_state_24_port);
   U33 : AND2_X1 port map( A1 => N40, A2 => n41_port, ZN => n_state_23_port);
   U34 : AND2_X1 port map( A1 => N39, A2 => n41_port, ZN => n_state_22_port);
   U35 : AND2_X1 port map( A1 => N38, A2 => n41_port, ZN => n_state_21_port);
   U36 : AND2_X1 port map( A1 => N37, A2 => n41_port, ZN => n_state_20_port);
   U37 : AND2_X1 port map( A1 => N18, A2 => n41_port, ZN => n_state_1_port);
   U38 : AND2_X1 port map( A1 => N36, A2 => n41_port, ZN => n_state_19_port);
   U39 : AND2_X1 port map( A1 => N35, A2 => n41_port, ZN => n_state_18_port);
   U40 : AND2_X1 port map( A1 => N34, A2 => n41_port, ZN => n_state_17_port);
   U41 : AND2_X1 port map( A1 => N33, A2 => n41_port, ZN => n_state_16_port);
   U42 : AND2_X1 port map( A1 => N32, A2 => n41_port, ZN => n_state_15_port);
   U43 : AND2_X1 port map( A1 => N31, A2 => n41_port, ZN => n_state_14_port);
   U44 : AND2_X1 port map( A1 => N30, A2 => n41_port, ZN => n_state_13_port);
   U45 : AND2_X1 port map( A1 => N29, A2 => n41_port, ZN => n_state_12_port);
   U46 : AND2_X1 port map( A1 => N28, A2 => n41_port, ZN => n_state_11_port);
   U47 : AND2_X1 port map( A1 => N27, A2 => n41_port, ZN => n_state_10_port);
   U48 : INV_X1 port map( A => n42_port, ZN => n_state_0_port);
   U49 : AOI21_X1 port map( B1 => n41_port, B2 => N17, A => n43_port, ZN => 
                           n42_port);
   U50 : AND4_X1 port map( A1 => en, A2 => n362, A3 => n44_port, A4 => n45_port
                           , ZN => n43_port);
   U51 : NOR2_X1 port map( A1 => lock, A2 => c_state_31_port, ZN => n44_port);
   U52 : OR2_X1 port map( A1 => n47_port, A2 => n48_port, ZN => n46_port);
   U53 : MUX2_X1 port map( A => n49, B => n45_port, S => n362, Z => n48_port);
   U54 : MUX2_X1 port map( A => a_adj_0_port, B => a_mod_0_port, S => n40_port,
                           Z => n361);
   U55 : MUX2_X1 port map( A => a_adj_1_port, B => a_mod_1_port, S => n39_port,
                           Z => n360);
   U56 : MUX2_X1 port map( A => a_adj_2_port, B => a_mod_2_port, S => n39_port,
                           Z => n359);
   U57 : MUX2_X1 port map( A => a_adj_3_port, B => a_mod_3_port, S => n39_port,
                           Z => n358);
   U58 : MUX2_X1 port map( A => a_adj_4_port, B => a_mod_4_port, S => n39_port,
                           Z => n357);
   U59 : MUX2_X1 port map( A => a_adj_5_port, B => a_mod_5_port, S => n39_port,
                           Z => n356);
   U60 : MUX2_X1 port map( A => a_adj_6_port, B => a_mod_6_port, S => n39_port,
                           Z => n355);
   U61 : MUX2_X1 port map( A => a_adj_7_port, B => a_mod_7_port, S => n39_port,
                           Z => n354);
   U62 : MUX2_X1 port map( A => a_adj_8_port, B => a_mod_8_port, S => n39_port,
                           Z => n353);
   U63 : MUX2_X1 port map( A => a_adj_9_port, B => a_mod_9_port, S => n39_port,
                           Z => n352);
   U64 : MUX2_X1 port map( A => a_adj_10_port, B => a_mod_10_port, S => 
                           n39_port, Z => n351);
   U65 : MUX2_X1 port map( A => a_adj_11_port, B => a_mod_11_port, S => 
                           n39_port, Z => n350);
   U66 : MUX2_X1 port map( A => a_adj_12_port, B => a_mod_12_port, S => 
                           n39_port, Z => n349);
   U67 : MUX2_X1 port map( A => a_adj_13_port, B => a_mod_13_port, S => 
                           n39_port, Z => n348);
   U68 : MUX2_X1 port map( A => a_adj_14_port, B => a_mod_14_port, S => 
                           n39_port, Z => n347);
   U69 : MUX2_X1 port map( A => a_adj_15_port, B => a_mod_15_port, S => 
                           n39_port, Z => n346);
   U70 : MUX2_X1 port map( A => a_adj_16_port, B => a_mod_16_port, S => 
                           n39_port, Z => n345);
   U71 : MUX2_X1 port map( A => a_adj_17_port, B => a_mod_17_port, S => 
                           n39_port, Z => n344);
   U72 : MUX2_X1 port map( A => a_adj_18_port, B => a_mod_18_port, S => 
                           n39_port, Z => n343);
   U73 : MUX2_X1 port map( A => a_adj_19_port, B => a_mod_19_port, S => 
                           n39_port, Z => n342);
   U74 : MUX2_X1 port map( A => a_adj_20_port, B => a_mod_20_port, S => 
                           n39_port, Z => n341);
   U75 : MUX2_X1 port map( A => a_adj_21_port, B => a_mod_21_port, S => 
                           n39_port, Z => n340);
   U76 : MUX2_X1 port map( A => a_adj_22_port, B => a_mod_22_port, S => 
                           n39_port, Z => n339);
   U77 : MUX2_X1 port map( A => a_adj_23_port, B => a_mod_23_port, S => 
                           n39_port, Z => n338);
   U78 : MUX2_X1 port map( A => a_adj_24_port, B => a_mod_24_port, S => 
                           n39_port, Z => n337);
   U79 : MUX2_X1 port map( A => a_adj_25_port, B => a_mod_25_port, S => 
                           n39_port, Z => n336);
   U80 : MUX2_X1 port map( A => a_adj_26_port, B => a_mod_26_port, S => 
                           n39_port, Z => n335);
   U81 : MUX2_X1 port map( A => a_adj_27_port, B => a_mod_27_port, S => 
                           n39_port, Z => n334);
   U82 : MUX2_X1 port map( A => a_adj_28_port, B => a_mod_28_port, S => 
                           n39_port, Z => n333);
   U83 : MUX2_X1 port map( A => a_adj_29_port, B => a_mod_29_port, S => 
                           n39_port, Z => n332);
   U84 : MUX2_X1 port map( A => a_adj_30_port, B => a_mod_30_port, S => 
                           n39_port, Z => n331);
   U85 : MUX2_X1 port map( A => a_adj_31_port, B => a_mod_31_port, S => 
                           n39_port, Z => n330);
   U86 : MUX2_X1 port map( A => b_adj_0_port, B => n31_port, S => n39_port, Z 
                           => n329);
   U87 : MUX2_X1 port map( A => b_adj_1_port, B => n70, S => n39_port, Z => 
                           n328);
   U88 : MUX2_X1 port map( A => b_adj_2_port, B => n30_port, S => n39_port, Z 
                           => n327);
   U89 : MUX2_X1 port map( A => b_adj_3_port, B => n29_port, S => n38_port, Z 
                           => n326);
   U90 : MUX2_X1 port map( A => b_adj_4_port, B => n28_port, S => n38_port, Z 
                           => n325);
   U91 : MUX2_X1 port map( A => b_adj_5_port, B => n27_port, S => n38_port, Z 
                           => n324);
   U92 : MUX2_X1 port map( A => b_adj_6_port, B => n26_port, S => n38_port, Z 
                           => n323);
   U93 : MUX2_X1 port map( A => b_adj_7_port, B => n25_port, S => n38_port, Z 
                           => n322);
   U94 : MUX2_X1 port map( A => b_adj_8_port, B => n24_port, S => n38_port, Z 
                           => n321);
   U95 : MUX2_X1 port map( A => b_adj_9_port, B => n23_port, S => n38_port, Z 
                           => n320);
   U96 : MUX2_X1 port map( A => b_adj_10_port, B => n22_port, S => n38_port, Z 
                           => n319);
   U97 : MUX2_X1 port map( A => b_adj_11_port, B => n21_port, S => n38_port, Z 
                           => n318);
   U98 : MUX2_X1 port map( A => b_adj_12_port, B => n20_port, S => n38_port, Z 
                           => n317);
   U99 : MUX2_X1 port map( A => b_adj_13_port, B => n19_port, S => n38_port, Z 
                           => n316);
   U100 : MUX2_X1 port map( A => b_adj_14_port, B => n18_port, S => n38_port, Z
                           => n315);
   U101 : MUX2_X1 port map( A => b_adj_15_port, B => n17_port, S => n38_port, Z
                           => n314);
   U102 : MUX2_X1 port map( A => b_adj_16_port, B => n16, S => n38_port, Z => 
                           n313);
   U103 : MUX2_X1 port map( A => b_adj_17_port, B => n15, S => n38_port, Z => 
                           n312);
   U104 : MUX2_X1 port map( A => b_adj_18_port, B => n14, S => n38_port, Z => 
                           n311);
   U105 : MUX2_X1 port map( A => b_adj_19_port, B => n13, S => n38_port, Z => 
                           n310);
   U106 : MUX2_X1 port map( A => b_adj_20_port, B => n12, S => n38_port, Z => 
                           n309);
   U107 : MUX2_X1 port map( A => b_adj_21_port, B => n11, S => n38_port, Z => 
                           n308);
   U108 : MUX2_X1 port map( A => b_adj_22_port, B => n10, S => n38_port, Z => 
                           n307);
   U109 : MUX2_X1 port map( A => b_adj_23_port, B => n9, S => n38_port, Z => 
                           n306);
   U110 : MUX2_X1 port map( A => b_adj_24_port, B => n8, S => n38_port, Z => 
                           n305);
   U111 : MUX2_X1 port map( A => b_adj_25_port, B => n7, S => n38_port, Z => 
                           n304);
   U112 : MUX2_X1 port map( A => b_adj_26_port, B => n6, S => n38_port, Z => 
                           n303);
   U113 : MUX2_X1 port map( A => b_adj_27_port, B => n5, S => n38_port, Z => 
                           n302);
   U114 : MUX2_X1 port map( A => b_adj_28_port, B => n4, S => n38_port, Z => 
                           n301);
   U115 : MUX2_X1 port map( A => b_adj_29_port, B => n3, S => n38_port, Z => 
                           n300);
   U116 : MUX2_X1 port map( A => b_adj_30_port, B => n2, S => n38_port, Z => 
                           n299);
   U117 : MUX2_X1 port map( A => b_adj_31_port, B => n1, S => n38_port, Z => 
                           n298);
   U118 : MUX2_X1 port map( A => n50, B => inv_q_flag_mod, S => n39_port, Z => 
                           n297);
   U119 : OAI22_X1 port map( A1 => a(31), A2 => n51, B1 => b(31), B2 => n52, ZN
                           => n50);
   U120 : NAND3_X1 port map( A1 => sign, A2 => n53, A3 => b(31), ZN => n51);
   U121 : NAND3_X1 port map( A1 => a(31), A2 => n53, A3 => sign, ZN => n52);
   U122 : OR2_X1 port map( A1 => n37_port, A2 => n54, ZN => en_r);
   U123 : NOR3_X1 port map( A1 => c_state_31_port, A2 => n362, A3 => n55, ZN =>
                           n54);
   U124 : INV_X1 port map( A => n55, ZN => n45_port);
   U125 : NAND4_X1 port map( A1 => n77, A2 => n78, A3 => n76, A4 => n56, ZN => 
                           n55);
   U126 : AND3_X1 port map( A1 => n82, A2 => n57, A3 => n373, ZN => n56);
   U127 : OAI211_X1 port map( C1 => n58, C2 => n59, A => n60, B => n57, ZN => 
                           n47_port);
   U128 : AND4_X1 port map( A1 => n61, A2 => n62, A3 => n63, A4 => n64, ZN => 
                           n57);
   U129 : NOR4_X1 port map( A1 => n65, A2 => c_state_28_port, A3 => 
                           c_state_24_port, A4 => c_state_23_port, ZN => n64);
   U130 : NAND4_X1 port map( A1 => n86, A2 => n374, A3 => n372, A4 => n371, ZN 
                           => n65);
   U131 : NOR4_X1 port map( A1 => n66, A2 => c_state_9_port, A3 => 
                           c_state_29_port, A4 => c_state_30_port, ZN => n63);
   U132 : NAND3_X1 port map( A1 => n84, A2 => n85, A3 => n83, ZN => n66);
   U133 : NOR4_X1 port map( A1 => n67, A2 => c_state_12_port, A3 => 
                           c_state_11_port, A4 => c_state_10_port, ZN => n62);
   U134 : NAND3_X1 port map( A1 => n80, A2 => n81, A3 => n79, ZN => n67);
   U135 : NOR4_X1 port map( A1 => n68, A2 => c_state_21_port, A3 => 
                           c_state_17_port, A4 => c_state_16_port, ZN => n61);
   U136 : NAND3_X1 port map( A1 => n74, A2 => n75, A3 => n73, ZN => n68);
   U137 : INV_X1 port map( A => n69, ZN => n60);
   U138 : AOI21_X1 port map( B1 => n53, B2 => n76, A => n82, ZN => n69);
   U139 : INV_X1 port map( A => n49, ZN => n59);
   U140 : OAI21_X1 port map( B1 => n76, B2 => n53, A => n82, ZN => n49);
   U141 : AND3_X1 port map( A1 => n77, A2 => n373, A3 => n78, ZN => n58);
   U142 : MUX2_X1 port map( A => b_shf_sqrt_63_port, B => n1, S => n53, Z => 
                           b_shf_63_port);
   U143 : MUX2_X1 port map( A => b_shf_sqrt_62_port, B => n2, S => n53, Z => 
                           b_shf_62_port);
   U144 : MUX2_X1 port map( A => b_shf_sqrt_61_port, B => n3, S => n53, Z => 
                           b_shf_61_port);
   U145 : MUX2_X1 port map( A => b_shf_sqrt_60_port, B => n4, S => n53, Z => 
                           b_shf_60_port);
   U146 : MUX2_X1 port map( A => b_shf_sqrt_59_port, B => n5, S => n53, Z => 
                           b_shf_59_port);
   U147 : MUX2_X1 port map( A => b_shf_sqrt_58_port, B => n6, S => n53, Z => 
                           b_shf_58_port);
   U148 : MUX2_X1 port map( A => b_shf_sqrt_57_port, B => n7, S => n53, Z => 
                           b_shf_57_port);
   U149 : MUX2_X1 port map( A => b_shf_sqrt_56_port, B => n8, S => n53, Z => 
                           b_shf_56_port);
   U150 : MUX2_X1 port map( A => b_shf_sqrt_55_port, B => n9, S => n53, Z => 
                           b_shf_55_port);
   U151 : MUX2_X1 port map( A => b_shf_sqrt_54_port, B => n10, S => n53, Z => 
                           b_shf_54_port);
   U152 : MUX2_X1 port map( A => b_shf_sqrt_53_port, B => n11, S => n53, Z => 
                           b_shf_53_port);
   U153 : MUX2_X1 port map( A => b_shf_sqrt_52_port, B => n12, S => n53, Z => 
                           b_shf_52_port);
   U154 : MUX2_X1 port map( A => b_shf_sqrt_51_port, B => n13, S => n53, Z => 
                           b_shf_51_port);
   U155 : MUX2_X1 port map( A => b_shf_sqrt_50_port, B => n14, S => n53, Z => 
                           b_shf_50_port);
   U156 : MUX2_X1 port map( A => b_shf_sqrt_49_port, B => n15, S => n53, Z => 
                           b_shf_49_port);
   U157 : MUX2_X1 port map( A => b_shf_sqrt_48_port, B => n16, S => n53, Z => 
                           b_shf_48_port);
   U158 : MUX2_X1 port map( A => b_shf_sqrt_47_port, B => n17_port, S => n53, Z
                           => b_shf_47_port);
   U159 : MUX2_X1 port map( A => b_shf_sqrt_46_port, B => n18_port, S => n53, Z
                           => b_shf_46_port);
   U160 : MUX2_X1 port map( A => b_shf_sqrt_45_port, B => n19_port, S => n53, Z
                           => b_shf_45_port);
   U161 : MUX2_X1 port map( A => b_shf_sqrt_44_port, B => n20_port, S => n53, Z
                           => b_shf_44_port);
   U162 : MUX2_X1 port map( A => b_shf_sqrt_43_port, B => n21_port, S => n53, Z
                           => b_shf_43_port);
   U163 : MUX2_X1 port map( A => b_shf_sqrt_42_port, B => n22_port, S => n53, Z
                           => b_shf_42_port);
   U164 : MUX2_X1 port map( A => b_shf_sqrt_41_port, B => n23_port, S => n53, Z
                           => b_shf_41_port);
   U165 : MUX2_X1 port map( A => b_shf_sqrt_40_port, B => n24_port, S => n53, Z
                           => b_shf_40_port);
   U166 : MUX2_X1 port map( A => b_shf_sqrt_39_port, B => n25_port, S => n53, Z
                           => b_shf_39_port);
   U167 : MUX2_X1 port map( A => b_shf_sqrt_38_port, B => n26_port, S => n53, Z
                           => b_shf_38_port);
   U168 : MUX2_X1 port map( A => b_shf_sqrt_37_port, B => n27_port, S => n53, Z
                           => b_shf_37_port);
   U169 : MUX2_X1 port map( A => b_shf_sqrt_36_port, B => n28_port, S => n53, Z
                           => b_shf_36_port);
   U170 : MUX2_X1 port map( A => b_shf_sqrt_35_port, B => n29_port, S => n53, Z
                           => b_shf_35_port);
   U171 : MUX2_X1 port map( A => b_shf_sqrt_34_port, B => n30_port, S => n53, Z
                           => b_shf_34_port);
   U172 : MUX2_X1 port map( A => a_mux_63_port, B => n70, S => n53, Z => 
                           b_shf_33_port);
   U173 : NAND2_X1 port map( A1 => n71, A2 => n53, ZN => b_shf_32_port);
   U174 : MUX2_X1 port map( A => a_mux_7_port, B => a_mux_8_port, S => n53, Z 
                           => a_shf_9_port);
   U175 : MUX2_X1 port map( A => a_mux_6_port, B => a_mux_7_port, S => n53, Z 
                           => a_shf_8_port);
   U176 : MUX2_X1 port map( A => a_mux_5_port, B => a_mux_6_port, S => n53, Z 
                           => a_shf_7_port);
   U177 : MUX2_X1 port map( A => a_mux_4_port, B => a_mux_5_port, S => n53, Z 
                           => a_shf_6_port);
   U178 : MUX2_X1 port map( A => a_mux_61_port, B => a_mux_62_port, S => n53, Z
                           => a_shf_63_port);
   U179 : MUX2_X1 port map( A => a_mux_60_port, B => a_mux_61_port, S => n53, Z
                           => a_shf_62_port);
   U180 : MUX2_X1 port map( A => a_mux_59_port, B => a_mux_60_port, S => n53, Z
                           => a_shf_61_port);
   U181 : MUX2_X1 port map( A => a_mux_58_port, B => a_mux_59_port, S => n53, Z
                           => a_shf_60_port);
   U182 : MUX2_X1 port map( A => a_mux_3_port, B => a_mux_4_port, S => n53, Z 
                           => a_shf_5_port);
   U183 : MUX2_X1 port map( A => a_mux_57_port, B => a_mux_58_port, S => n53, Z
                           => a_shf_59_port);
   U184 : MUX2_X1 port map( A => a_mux_56_port, B => a_mux_57_port, S => n53, Z
                           => a_shf_58_port);
   U185 : MUX2_X1 port map( A => a_mux_55_port, B => a_mux_56_port, S => n53, Z
                           => a_shf_57_port);
   U186 : MUX2_X1 port map( A => a_mux_54_port, B => a_mux_55_port, S => n53, Z
                           => a_shf_56_port);
   U187 : MUX2_X1 port map( A => a_mux_53_port, B => a_mux_54_port, S => n53, Z
                           => a_shf_55_port);
   U188 : MUX2_X1 port map( A => a_mux_52_port, B => a_mux_53_port, S => n53, Z
                           => a_shf_54_port);
   U189 : MUX2_X1 port map( A => a_mux_51_port, B => a_mux_52_port, S => n53, Z
                           => a_shf_53_port);
   U190 : MUX2_X1 port map( A => a_mux_50_port, B => a_mux_51_port, S => n53, Z
                           => a_shf_52_port);
   U191 : MUX2_X1 port map( A => a_mux_49_port, B => a_mux_50_port, S => n53, Z
                           => a_shf_51_port);
   U192 : MUX2_X1 port map( A => a_mux_48_port, B => a_mux_49_port, S => n53, Z
                           => a_shf_50_port);
   U193 : MUX2_X1 port map( A => a_mux_2_port, B => a_mux_3_port, S => n53, Z 
                           => a_shf_4_port);
   U194 : MUX2_X1 port map( A => a_mux_47_port, B => a_mux_48_port, S => n53, Z
                           => a_shf_49_port);
   U195 : MUX2_X1 port map( A => a_mux_46_port, B => a_mux_47_port, S => n53, Z
                           => a_shf_48_port);
   U196 : MUX2_X1 port map( A => a_mux_45_port, B => a_mux_46_port, S => n53, Z
                           => a_shf_47_port);
   U197 : MUX2_X1 port map( A => a_mux_44_port, B => a_mux_45_port, S => n53, Z
                           => a_shf_46_port);
   U198 : MUX2_X1 port map( A => a_mux_43_port, B => a_mux_44_port, S => n53, Z
                           => a_shf_45_port);
   U199 : MUX2_X1 port map( A => a_mux_42_port, B => a_mux_43_port, S => n53, Z
                           => a_shf_44_port);
   U200 : MUX2_X1 port map( A => a_mux_41_port, B => a_mux_42_port, S => n53, Z
                           => a_shf_43_port);
   U201 : MUX2_X1 port map( A => a_mux_40_port, B => a_mux_41_port, S => n53, Z
                           => a_shf_42_port);
   U202 : MUX2_X1 port map( A => a_mux_39_port, B => a_mux_40_port, S => n53, Z
                           => a_shf_41_port);
   U203 : MUX2_X1 port map( A => a_mux_38_port, B => a_mux_39_port, S => n53, Z
                           => a_shf_40_port);
   U204 : MUX2_X1 port map( A => a_mux_1_port, B => a_mux_2_port, S => n53, Z 
                           => a_shf_3_port);
   U205 : MUX2_X1 port map( A => a_mux_37_port, B => a_mux_38_port, S => n53, Z
                           => a_shf_39_port);
   U206 : MUX2_X1 port map( A => a_mux_36_port, B => a_mux_37_port, S => n53, Z
                           => a_shf_38_port);
   U207 : MUX2_X1 port map( A => a_mux_35_port, B => a_mux_36_port, S => n53, Z
                           => a_shf_37_port);
   U208 : MUX2_X1 port map( A => a_mux_34_port, B => a_mux_35_port, S => n53, Z
                           => a_shf_36_port);
   U209 : MUX2_X1 port map( A => a_mux_33_port, B => a_mux_34_port, S => n53, Z
                           => a_shf_35_port);
   U210 : MUX2_X1 port map( A => a_mux_32_port, B => a_mux_33_port, S => n53, Z
                           => a_shf_34_port);
   U211 : MUX2_X1 port map( A => a_mux_31_port, B => a_mux_32_port, S => n53, Z
                           => a_shf_33_port);
   U212 : MUX2_X1 port map( A => a_mux_30_port, B => a_mux_31_port, S => n53, Z
                           => a_shf_32_port);
   U213 : MUX2_X1 port map( A => a_mux_29_port, B => a_mux_30_port, S => n53, Z
                           => a_shf_31_port);
   U214 : MUX2_X1 port map( A => a_mux_28_port, B => a_mux_29_port, S => n53, Z
                           => a_shf_30_port);
   U215 : MUX2_X1 port map( A => a_mux_0_port, B => a_mux_1_port, S => n53, Z 
                           => a_shf_2_port);
   U216 : MUX2_X1 port map( A => a_mux_27_port, B => a_mux_28_port, S => n53, Z
                           => a_shf_29_port);
   U217 : MUX2_X1 port map( A => a_mux_26_port, B => a_mux_27_port, S => n53, Z
                           => a_shf_28_port);
   U218 : MUX2_X1 port map( A => a_mux_25_port, B => a_mux_26_port, S => n53, Z
                           => a_shf_27_port);
   U219 : MUX2_X1 port map( A => a_mux_24_port, B => a_mux_25_port, S => n53, Z
                           => a_shf_26_port);
   U220 : MUX2_X1 port map( A => a_mux_23_port, B => a_mux_24_port, S => n53, Z
                           => a_shf_25_port);
   U221 : MUX2_X1 port map( A => a_mux_22_port, B => a_mux_23_port, S => n53, Z
                           => a_shf_24_port);
   U222 : MUX2_X1 port map( A => a_mux_21_port, B => a_mux_22_port, S => n53, Z
                           => a_shf_23_port);
   U223 : MUX2_X1 port map( A => a_mux_20_port, B => a_mux_21_port, S => n53, Z
                           => a_shf_22_port);
   U224 : MUX2_X1 port map( A => a_mux_19_port, B => a_mux_20_port, S => n53, Z
                           => a_shf_21_port);
   U225 : MUX2_X1 port map( A => a_mux_18_port, B => a_mux_19_port, S => n53, Z
                           => a_shf_20_port);
   U226 : AND2_X1 port map( A1 => n53, A2 => a_mux_0_port, ZN => a_shf_1_port);
   U227 : MUX2_X1 port map( A => a_mux_17_port, B => a_mux_18_port, S => n53, Z
                           => a_shf_19_port);
   U228 : MUX2_X1 port map( A => a_mux_16_port, B => a_mux_17_port, S => n53, Z
                           => a_shf_18_port);
   U229 : MUX2_X1 port map( A => a_mux_15_port, B => a_mux_16_port, S => n53, Z
                           => a_shf_17_port);
   U230 : MUX2_X1 port map( A => a_mux_14_port, B => a_mux_15_port, S => n53, Z
                           => a_shf_16_port);
   U231 : MUX2_X1 port map( A => a_mux_13_port, B => a_mux_14_port, S => n53, Z
                           => a_shf_15_port);
   U232 : MUX2_X1 port map( A => a_mux_12_port, B => a_mux_13_port, S => n53, Z
                           => a_shf_14_port);
   U233 : MUX2_X1 port map( A => a_mux_11_port, B => a_mux_12_port, S => n53, Z
                           => a_shf_13_port);
   U234 : MUX2_X1 port map( A => a_mux_10_port, B => a_mux_11_port, S => n53, Z
                           => a_shf_12_port);
   U235 : MUX2_X1 port map( A => a_mux_9_port, B => a_mux_10_port, S => n53, Z 
                           => a_shf_11_port);
   U236 : MUX2_X1 port map( A => a_mux_8_port, B => a_mux_9_port, S => n53, Z 
                           => a_shf_10_port);

end SYN_div_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mul_DATA_SIZE16_STAGE10 is

   port( rst, clk, en, lock, sign : in std_logic;  a, b : in std_logic_vector 
         (15 downto 0);  o : out std_logic_vector (31 downto 0));

end Mul_DATA_SIZE16_STAGE10;

architecture SYN_mul_arch_struct of Mul_DATA_SIZE16_STAGE10 is

   component BoothMul_DATA_SIZE16_STAGE10
      port( rst, clk, en, lock, sign : in std_logic;  a, b : in 
            std_logic_vector (15 downto 0);  o : out std_logic_vector (31 
            downto 0));
   end component;

begin
   
   BM0 : BoothMul_DATA_SIZE16_STAGE10 port map( rst => rst, clk => clk, en => 
                           en, lock => lock, sign => sign, a(15) => a(15), 
                           a(14) => a(14), a(13) => a(13), a(12) => a(12), 
                           a(11) => a(11), a(10) => a(10), a(9) => a(9), a(8) 
                           => a(8), a(7) => a(7), a(6) => a(6), a(5) => a(5), 
                           a(4) => a(4), a(3) => a(3), a(2) => a(2), a(1) => 
                           a(1), a(0) => a(0), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           o(31) => o(31), o(30) => o(30), o(29) => o(29), 
                           o(28) => o(28), o(27) => o(27), o(26) => o(26), 
                           o(25) => o(25), o(24) => o(24), o(23) => o(23), 
                           o(22) => o(22), o(21) => o(21), o(20) => o(20), 
                           o(19) => o(19), o(18) => o(18), o(17) => o(17), 
                           o(16) => o(16), o(15) => o(15), o(14) => o(14), 
                           o(13) => o(13), o(12) => o(12), o(11) => o(11), 
                           o(10) => o(10), o(9) => o(9), o(8) => o(8), o(7) => 
                           o(7), o(6) => o(6), o(5) => o(5), o(4) => o(4), o(3)
                           => o(3), o(2) => o(2), o(1) => o(1), o(0) => o(0));

end SYN_mul_arch_struct;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Alu_DATA_SIZE32 is

   port( f : in std_logic_vector (4 downto 0);  a, b : in std_logic_vector (31 
         downto 0);  o : out std_logic_vector (31 downto 0));

end Alu_DATA_SIZE32;

architecture SYN_alu_arch of Alu_DATA_SIZE32 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component Shifter_DATA_SIZE32
      port( l_r, l_a, s_r : in std_logic;  a, b : in std_logic_vector (31 
            downto 0);  o : out std_logic_vector (31 downto 0));
   end component;
   
   component Adder_DATA_SIZE32_6
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;
   
   signal X_Logic0_port, b_new_31_port, b_new_30_port, b_new_29_port, 
      b_new_28_port, b_new_27_port, b_new_26_port, b_new_25_port, b_new_24_port
      , b_new_23_port, b_new_22_port, b_new_21_port, b_new_20_port, 
      b_new_19_port, b_new_18_port, b_new_17_port, b_new_16_port, b_new_15_port
      , b_new_14_port, b_new_13_port, b_new_12_port, b_new_11_port, 
      b_new_10_port, b_new_9_port, b_new_8_port, b_new_7_port, b_new_6_port, 
      b_new_5_port, b_new_4_port, b_new_3_port, b_new_2_port, b_new_1_port, 
      b_new_0_port, ado_31_port, ado_30_port, ado_29_port, ado_28_port, 
      ado_27_port, ado_26_port, ado_25_port, ado_24_port, ado_23_port, 
      ado_22_port, ado_21_port, ado_20_port, ado_19_port, ado_18_port, 
      ado_17_port, ado_16_port, ado_15_port, ado_14_port, ado_13_port, 
      ado_12_port, ado_11_port, ado_10_port, ado_9_port, ado_8_port, ado_7_port
      , ado_6_port, ado_5_port, ado_4_port, ado_3_port, ado_2_port, ado_1_port,
      ado_0_port, c_f, sho_31_port, sho_30_port, sho_29_port, sho_28_port, 
      sho_27_port, sho_26_port, sho_25_port, sho_24_port, sho_23_port, 
      sho_22_port, sho_21_port, sho_20_port, sho_19_port, sho_18_port, 
      sho_17_port, sho_16_port, sho_15_port, sho_14_port, sho_13_port, 
      sho_12_port, sho_11_port, sho_10_port, sho_9_port, sho_8_port, sho_7_port
      , sho_6_port, sho_5_port, sho_4_port, sho_3_port, sho_2_port, sho_1_port,
      sho_0_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, 
      n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29
      , n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, 
      n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58
      , n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, 
      n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87
      , n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
      n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, 
      n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, 
      n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, 
      n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, 
      n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232 : 
      std_logic;

begin
   
   X_Logic0_port <= '0';
   ADD0 : Adder_DATA_SIZE32_6 port map( cin => f(4), a(31) => a(31), a(30) => 
                           a(30), a(29) => a(29), a(28) => a(28), a(27) => 
                           a(27), a(26) => a(26), a(25) => a(25), a(24) => 
                           a(24), a(23) => a(23), a(22) => a(22), a(21) => 
                           a(21), a(20) => a(20), a(19) => a(19), a(18) => 
                           a(18), a(17) => a(17), a(16) => a(16), a(15) => 
                           a(15), a(14) => a(14), a(13) => a(13), a(12) => 
                           a(12), a(11) => a(11), a(10) => a(10), a(9) => a(9),
                           a(8) => a(8), a(7) => a(7), a(6) => a(6), a(5) => 
                           a(5), a(4) => a(4), a(3) => a(3), a(2) => a(2), a(1)
                           => a(1), a(0) => a(0), b(31) => b_new_31_port, b(30)
                           => b_new_30_port, b(29) => b_new_29_port, b(28) => 
                           b_new_28_port, b(27) => b_new_27_port, b(26) => 
                           b_new_26_port, b(25) => b_new_25_port, b(24) => 
                           b_new_24_port, b(23) => b_new_23_port, b(22) => 
                           b_new_22_port, b(21) => b_new_21_port, b(20) => 
                           b_new_20_port, b(19) => b_new_19_port, b(18) => 
                           b_new_18_port, b(17) => b_new_17_port, b(16) => 
                           b_new_16_port, b(15) => b_new_15_port, b(14) => 
                           b_new_14_port, b(13) => b_new_13_port, b(12) => 
                           b_new_12_port, b(11) => b_new_11_port, b(10) => 
                           b_new_10_port, b(9) => b_new_9_port, b(8) => 
                           b_new_8_port, b(7) => b_new_7_port, b(6) => 
                           b_new_6_port, b(5) => b_new_5_port, b(4) => 
                           b_new_4_port, b(3) => b_new_3_port, b(2) => 
                           b_new_2_port, b(1) => b_new_1_port, b(0) => 
                           b_new_0_port, s(31) => ado_31_port, s(30) => 
                           ado_30_port, s(29) => ado_29_port, s(28) => 
                           ado_28_port, s(27) => ado_27_port, s(26) => 
                           ado_26_port, s(25) => ado_25_port, s(24) => 
                           ado_24_port, s(23) => ado_23_port, s(22) => 
                           ado_22_port, s(21) => ado_21_port, s(20) => 
                           ado_20_port, s(19) => ado_19_port, s(18) => 
                           ado_18_port, s(17) => ado_17_port, s(16) => 
                           ado_16_port, s(15) => ado_15_port, s(14) => 
                           ado_14_port, s(13) => ado_13_port, s(12) => 
                           ado_12_port, s(11) => ado_11_port, s(10) => 
                           ado_10_port, s(9) => ado_9_port, s(8) => ado_8_port,
                           s(7) => ado_7_port, s(6) => ado_6_port, s(5) => 
                           ado_5_port, s(4) => ado_4_port, s(3) => ado_3_port, 
                           s(2) => ado_2_port, s(1) => ado_1_port, s(0) => 
                           ado_0_port, cout => c_f);
   SHF0 : Shifter_DATA_SIZE32 port map( l_r => f(0), l_a => f(1), s_r => 
                           X_Logic0_port, a(31) => a(31), a(30) => a(30), a(29)
                           => a(29), a(28) => a(28), a(27) => a(27), a(26) => 
                           a(26), a(25) => a(25), a(24) => a(24), a(23) => 
                           a(23), a(22) => a(22), a(21) => a(21), a(20) => 
                           a(20), a(19) => a(19), a(18) => a(18), a(17) => 
                           a(17), a(16) => a(16), a(15) => a(15), a(14) => 
                           a(14), a(13) => a(13), a(12) => a(12), a(11) => 
                           a(11), a(10) => a(10), a(9) => a(9), a(8) => a(8), 
                           a(7) => a(7), a(6) => a(6), a(5) => a(5), a(4) => 
                           a(4), a(3) => a(3), a(2) => a(2), a(1) => a(1), a(0)
                           => a(0), b(31) => b(31), b(30) => b(30), b(29) => 
                           b(29), b(28) => b(28), b(27) => b(27), b(26) => 
                           b(26), b(25) => b(25), b(24) => b(24), b(23) => 
                           b(23), b(22) => b(22), b(21) => b(21), b(20) => 
                           b(20), b(19) => b(19), b(18) => b(18), b(17) => 
                           b(17), b(16) => b(16), b(15) => b(15), b(14) => 
                           b(14), b(13) => b(13), b(12) => b(12), b(11) => 
                           b(11), b(10) => b(10), b(9) => b(9), b(8) => b(8), 
                           b(7) => b(7), b(6) => b(6), b(5) => b(5), b(4) => 
                           b(4), b(3) => b(3), b(2) => b(2), b(1) => b(1), b(0)
                           => b(0), o(31) => sho_31_port, o(30) => sho_30_port,
                           o(29) => sho_29_port, o(28) => sho_28_port, o(27) =>
                           sho_27_port, o(26) => sho_26_port, o(25) => 
                           sho_25_port, o(24) => sho_24_port, o(23) => 
                           sho_23_port, o(22) => sho_22_port, o(21) => 
                           sho_21_port, o(20) => sho_20_port, o(19) => 
                           sho_19_port, o(18) => sho_18_port, o(17) => 
                           sho_17_port, o(16) => sho_16_port, o(15) => 
                           sho_15_port, o(14) => sho_14_port, o(13) => 
                           sho_13_port, o(12) => sho_12_port, o(11) => 
                           sho_11_port, o(10) => sho_10_port, o(9) => 
                           sho_9_port, o(8) => sho_8_port, o(7) => sho_7_port, 
                           o(6) => sho_6_port, o(5) => sho_5_port, o(4) => 
                           sho_4_port, o(3) => sho_3_port, o(2) => sho_2_port, 
                           o(1) => sho_1_port, o(0) => sho_0_port);
   U2 : NAND2_X4 port map( A1 => n203, A2 => f(1), ZN => n11);
   U3 : NAND2_X2 port map( A1 => n202, A2 => n203, ZN => n10);
   U4 : OR3_X1 port map( A1 => f(2), A2 => f(3), A3 => n207, ZN => n1);
   U5 : INV_X2 port map( A => n1, ZN => n2);
   U6 : OR4_X1 port map( A1 => n206, A2 => n202, A3 => f(3), A4 => f(4), ZN => 
                           n3);
   U7 : INV_X2 port map( A => n3, ZN => n4);
   U8 : INV_X1 port map( A => n5, ZN => o(9));
   U9 : AOI221_X1 port map( B1 => ado_9_port, B2 => n2, C1 => sho_9_port, C2 =>
                           n4, A => n6, ZN => n5);
   U10 : MUX2_X1 port map( A => n7, B => n8, S => a(9), Z => n6);
   U11 : NAND2_X1 port map( A1 => n9, A2 => n10, ZN => n8);
   U12 : MUX2_X1 port map( A => n11, B => n12, S => b(9), Z => n9);
   U13 : NOR2_X1 port map( A1 => n11, A2 => n13, ZN => n7);
   U14 : INV_X1 port map( A => b(9), ZN => n13);
   U15 : INV_X1 port map( A => n14, ZN => o(8));
   U16 : AOI221_X1 port map( B1 => ado_8_port, B2 => n2, C1 => sho_8_port, C2 
                           => n4, A => n15, ZN => n14);
   U17 : MUX2_X1 port map( A => n16, B => n17, S => a(8), Z => n15);
   U18 : NAND2_X1 port map( A1 => n18, A2 => n10, ZN => n17);
   U19 : MUX2_X1 port map( A => n11, B => n12, S => b(8), Z => n18);
   U20 : NOR2_X1 port map( A1 => n11, A2 => n19, ZN => n16);
   U21 : INV_X1 port map( A => b(8), ZN => n19);
   U22 : INV_X1 port map( A => n20, ZN => o(7));
   U23 : AOI221_X1 port map( B1 => ado_7_port, B2 => n2, C1 => sho_7_port, C2 
                           => n4, A => n21, ZN => n20);
   U24 : MUX2_X1 port map( A => n22, B => n23, S => a(7), Z => n21);
   U25 : NAND2_X1 port map( A1 => n24, A2 => n10, ZN => n23);
   U26 : MUX2_X1 port map( A => n11, B => n12, S => b(7), Z => n24);
   U27 : NOR2_X1 port map( A1 => n11, A2 => n25, ZN => n22);
   U28 : INV_X1 port map( A => b(7), ZN => n25);
   U29 : INV_X1 port map( A => n26, ZN => o(6));
   U30 : AOI221_X1 port map( B1 => ado_6_port, B2 => n2, C1 => sho_6_port, C2 
                           => n4, A => n27, ZN => n26);
   U31 : MUX2_X1 port map( A => n28, B => n29, S => a(6), Z => n27);
   U32 : NAND2_X1 port map( A1 => n30, A2 => n10, ZN => n29);
   U33 : MUX2_X1 port map( A => n11, B => n12, S => b(6), Z => n30);
   U34 : NOR2_X1 port map( A1 => n11, A2 => n31, ZN => n28);
   U35 : INV_X1 port map( A => b(6), ZN => n31);
   U36 : INV_X1 port map( A => n32, ZN => o(5));
   U37 : AOI221_X1 port map( B1 => ado_5_port, B2 => n2, C1 => sho_5_port, C2 
                           => n4, A => n33, ZN => n32);
   U38 : MUX2_X1 port map( A => n34, B => n35, S => a(5), Z => n33);
   U39 : NAND2_X1 port map( A1 => n36, A2 => n10, ZN => n35);
   U40 : MUX2_X1 port map( A => n11, B => n12, S => b(5), Z => n36);
   U41 : NOR2_X1 port map( A1 => n11, A2 => n37, ZN => n34);
   U42 : INV_X1 port map( A => b(5), ZN => n37);
   U43 : INV_X1 port map( A => n38, ZN => o(4));
   U44 : AOI221_X1 port map( B1 => ado_4_port, B2 => n2, C1 => sho_4_port, C2 
                           => n4, A => n39, ZN => n38);
   U45 : MUX2_X1 port map( A => n40, B => n41, S => a(4), Z => n39);
   U46 : NAND2_X1 port map( A1 => n42, A2 => n10, ZN => n41);
   U47 : MUX2_X1 port map( A => n11, B => n12, S => b(4), Z => n42);
   U48 : NOR2_X1 port map( A1 => n11, A2 => n43, ZN => n40);
   U49 : INV_X1 port map( A => b(4), ZN => n43);
   U50 : INV_X1 port map( A => n44, ZN => o(3));
   U51 : AOI221_X1 port map( B1 => ado_3_port, B2 => n2, C1 => sho_3_port, C2 
                           => n4, A => n45, ZN => n44);
   U52 : MUX2_X1 port map( A => n46, B => n47, S => a(3), Z => n45);
   U53 : NAND2_X1 port map( A1 => n48, A2 => n10, ZN => n47);
   U54 : MUX2_X1 port map( A => n11, B => n12, S => b(3), Z => n48);
   U55 : NOR2_X1 port map( A1 => n11, A2 => n49, ZN => n46);
   U56 : INV_X1 port map( A => b(3), ZN => n49);
   U57 : INV_X1 port map( A => n50, ZN => o(31));
   U58 : AOI221_X1 port map( B1 => ado_31_port, B2 => n2, C1 => sho_31_port, C2
                           => n4, A => n51, ZN => n50);
   U59 : MUX2_X1 port map( A => n52, B => n53, S => a(31), Z => n51);
   U60 : NAND2_X1 port map( A1 => n54, A2 => n10, ZN => n53);
   U61 : MUX2_X1 port map( A => n11, B => n12, S => b(31), Z => n54);
   U62 : NOR2_X1 port map( A1 => n11, A2 => n55, ZN => n52);
   U63 : INV_X1 port map( A => b(31), ZN => n55);
   U64 : INV_X1 port map( A => n56, ZN => o(30));
   U65 : AOI221_X1 port map( B1 => ado_30_port, B2 => n2, C1 => sho_30_port, C2
                           => n4, A => n57, ZN => n56);
   U66 : MUX2_X1 port map( A => n58, B => n59, S => a(30), Z => n57);
   U67 : NAND2_X1 port map( A1 => n60, A2 => n10, ZN => n59);
   U68 : MUX2_X1 port map( A => n11, B => n12, S => b(30), Z => n60);
   U69 : NOR2_X1 port map( A1 => n11, A2 => n61, ZN => n58);
   U70 : INV_X1 port map( A => b(30), ZN => n61);
   U71 : INV_X1 port map( A => n62, ZN => o(2));
   U72 : AOI221_X1 port map( B1 => ado_2_port, B2 => n2, C1 => sho_2_port, C2 
                           => n4, A => n63, ZN => n62);
   U73 : MUX2_X1 port map( A => n64, B => n65, S => a(2), Z => n63);
   U74 : NAND2_X1 port map( A1 => n66, A2 => n10, ZN => n65);
   U75 : MUX2_X1 port map( A => n11, B => n12, S => b(2), Z => n66);
   U76 : NOR2_X1 port map( A1 => n11, A2 => n67, ZN => n64);
   U77 : INV_X1 port map( A => b(2), ZN => n67);
   U78 : INV_X1 port map( A => n68, ZN => o(29));
   U79 : AOI221_X1 port map( B1 => ado_29_port, B2 => n2, C1 => sho_29_port, C2
                           => n4, A => n69, ZN => n68);
   U80 : MUX2_X1 port map( A => n70, B => n71, S => a(29), Z => n69);
   U81 : NAND2_X1 port map( A1 => n72, A2 => n10, ZN => n71);
   U82 : MUX2_X1 port map( A => n11, B => n12, S => b(29), Z => n72);
   U83 : NOR2_X1 port map( A1 => n11, A2 => n73, ZN => n70);
   U84 : INV_X1 port map( A => b(29), ZN => n73);
   U85 : INV_X1 port map( A => n74, ZN => o(28));
   U86 : AOI221_X1 port map( B1 => ado_28_port, B2 => n2, C1 => sho_28_port, C2
                           => n4, A => n75, ZN => n74);
   U87 : MUX2_X1 port map( A => n76, B => n77, S => a(28), Z => n75);
   U88 : NAND2_X1 port map( A1 => n78, A2 => n10, ZN => n77);
   U89 : MUX2_X1 port map( A => n11, B => n12, S => b(28), Z => n78);
   U90 : NOR2_X1 port map( A1 => n11, A2 => n79, ZN => n76);
   U91 : INV_X1 port map( A => b(28), ZN => n79);
   U92 : INV_X1 port map( A => n80, ZN => o(27));
   U93 : AOI221_X1 port map( B1 => ado_27_port, B2 => n2, C1 => sho_27_port, C2
                           => n4, A => n81, ZN => n80);
   U94 : MUX2_X1 port map( A => n82, B => n83, S => a(27), Z => n81);
   U95 : NAND2_X1 port map( A1 => n84, A2 => n10, ZN => n83);
   U96 : MUX2_X1 port map( A => n11, B => n12, S => b(27), Z => n84);
   U97 : NOR2_X1 port map( A1 => n11, A2 => n85, ZN => n82);
   U98 : INV_X1 port map( A => b(27), ZN => n85);
   U99 : INV_X1 port map( A => n86, ZN => o(26));
   U100 : AOI221_X1 port map( B1 => ado_26_port, B2 => n2, C1 => sho_26_port, 
                           C2 => n4, A => n87, ZN => n86);
   U101 : MUX2_X1 port map( A => n88, B => n89, S => a(26), Z => n87);
   U102 : NAND2_X1 port map( A1 => n90, A2 => n10, ZN => n89);
   U103 : MUX2_X1 port map( A => n11, B => n12, S => b(26), Z => n90);
   U104 : NOR2_X1 port map( A1 => n11, A2 => n91, ZN => n88);
   U105 : INV_X1 port map( A => b(26), ZN => n91);
   U106 : INV_X1 port map( A => n92, ZN => o(25));
   U107 : AOI221_X1 port map( B1 => ado_25_port, B2 => n2, C1 => sho_25_port, 
                           C2 => n4, A => n93, ZN => n92);
   U108 : MUX2_X1 port map( A => n94, B => n95, S => a(25), Z => n93);
   U109 : NAND2_X1 port map( A1 => n96, A2 => n10, ZN => n95);
   U110 : MUX2_X1 port map( A => n11, B => n12, S => b(25), Z => n96);
   U111 : NOR2_X1 port map( A1 => n11, A2 => n97, ZN => n94);
   U112 : INV_X1 port map( A => b(25), ZN => n97);
   U113 : INV_X1 port map( A => n98, ZN => o(24));
   U114 : AOI221_X1 port map( B1 => ado_24_port, B2 => n2, C1 => sho_24_port, 
                           C2 => n4, A => n99, ZN => n98);
   U115 : MUX2_X1 port map( A => n100, B => n101, S => a(24), Z => n99);
   U116 : NAND2_X1 port map( A1 => n102, A2 => n10, ZN => n101);
   U117 : MUX2_X1 port map( A => n11, B => n12, S => b(24), Z => n102);
   U118 : NOR2_X1 port map( A1 => n11, A2 => n103, ZN => n100);
   U119 : INV_X1 port map( A => b(24), ZN => n103);
   U120 : INV_X1 port map( A => n104, ZN => o(23));
   U121 : AOI221_X1 port map( B1 => ado_23_port, B2 => n2, C1 => sho_23_port, 
                           C2 => n4, A => n105, ZN => n104);
   U122 : MUX2_X1 port map( A => n106, B => n107, S => a(23), Z => n105);
   U123 : NAND2_X1 port map( A1 => n108, A2 => n10, ZN => n107);
   U124 : MUX2_X1 port map( A => n11, B => n12, S => b(23), Z => n108);
   U125 : NOR2_X1 port map( A1 => n11, A2 => n109, ZN => n106);
   U126 : INV_X1 port map( A => b(23), ZN => n109);
   U127 : INV_X1 port map( A => n110, ZN => o(22));
   U128 : AOI221_X1 port map( B1 => ado_22_port, B2 => n2, C1 => sho_22_port, 
                           C2 => n4, A => n111, ZN => n110);
   U129 : MUX2_X1 port map( A => n112, B => n113, S => a(22), Z => n111);
   U130 : NAND2_X1 port map( A1 => n114, A2 => n10, ZN => n113);
   U131 : MUX2_X1 port map( A => n11, B => n12, S => b(22), Z => n114);
   U132 : NOR2_X1 port map( A1 => n11, A2 => n115, ZN => n112);
   U133 : INV_X1 port map( A => b(22), ZN => n115);
   U134 : INV_X1 port map( A => n116, ZN => o(21));
   U135 : AOI221_X1 port map( B1 => ado_21_port, B2 => n2, C1 => sho_21_port, 
                           C2 => n4, A => n117, ZN => n116);
   U136 : MUX2_X1 port map( A => n118, B => n119, S => a(21), Z => n117);
   U137 : NAND2_X1 port map( A1 => n120, A2 => n10, ZN => n119);
   U138 : MUX2_X1 port map( A => n11, B => n12, S => b(21), Z => n120);
   U139 : NOR2_X1 port map( A1 => n11, A2 => n121, ZN => n118);
   U140 : INV_X1 port map( A => b(21), ZN => n121);
   U141 : INV_X1 port map( A => n122, ZN => o(20));
   U142 : AOI221_X1 port map( B1 => ado_20_port, B2 => n2, C1 => sho_20_port, 
                           C2 => n4, A => n123, ZN => n122);
   U143 : MUX2_X1 port map( A => n124, B => n125, S => a(20), Z => n123);
   U144 : NAND2_X1 port map( A1 => n126, A2 => n10, ZN => n125);
   U145 : MUX2_X1 port map( A => n11, B => n12, S => b(20), Z => n126);
   U146 : NOR2_X1 port map( A1 => n11, A2 => n127, ZN => n124);
   U147 : INV_X1 port map( A => b(20), ZN => n127);
   U148 : INV_X1 port map( A => n128, ZN => o(1));
   U149 : AOI221_X1 port map( B1 => ado_1_port, B2 => n2, C1 => sho_1_port, C2 
                           => n4, A => n129, ZN => n128);
   U150 : MUX2_X1 port map( A => n130, B => n131, S => a(1), Z => n129);
   U151 : NAND2_X1 port map( A1 => n132, A2 => n10, ZN => n131);
   U152 : MUX2_X1 port map( A => n11, B => n12, S => b(1), Z => n132);
   U153 : NOR2_X1 port map( A1 => n11, A2 => n133, ZN => n130);
   U154 : INV_X1 port map( A => b(1), ZN => n133);
   U155 : INV_X1 port map( A => n134, ZN => o(19));
   U156 : AOI221_X1 port map( B1 => ado_19_port, B2 => n2, C1 => sho_19_port, 
                           C2 => n4, A => n135, ZN => n134);
   U157 : MUX2_X1 port map( A => n136, B => n137, S => a(19), Z => n135);
   U158 : NAND2_X1 port map( A1 => n138, A2 => n10, ZN => n137);
   U159 : MUX2_X1 port map( A => n11, B => n12, S => b(19), Z => n138);
   U160 : NOR2_X1 port map( A1 => n11, A2 => n139, ZN => n136);
   U161 : INV_X1 port map( A => b(19), ZN => n139);
   U162 : INV_X1 port map( A => n140, ZN => o(18));
   U163 : AOI221_X1 port map( B1 => ado_18_port, B2 => n2, C1 => sho_18_port, 
                           C2 => n4, A => n141, ZN => n140);
   U164 : MUX2_X1 port map( A => n142, B => n143, S => a(18), Z => n141);
   U165 : NAND2_X1 port map( A1 => n144, A2 => n10, ZN => n143);
   U166 : MUX2_X1 port map( A => n11, B => n12, S => b(18), Z => n144);
   U167 : NOR2_X1 port map( A1 => n11, A2 => n145, ZN => n142);
   U168 : INV_X1 port map( A => b(18), ZN => n145);
   U169 : INV_X1 port map( A => n146, ZN => o(17));
   U170 : AOI221_X1 port map( B1 => ado_17_port, B2 => n2, C1 => sho_17_port, 
                           C2 => n4, A => n147, ZN => n146);
   U171 : MUX2_X1 port map( A => n148, B => n149, S => a(17), Z => n147);
   U172 : NAND2_X1 port map( A1 => n150, A2 => n10, ZN => n149);
   U173 : MUX2_X1 port map( A => n11, B => n12, S => b(17), Z => n150);
   U174 : NOR2_X1 port map( A1 => n11, A2 => n151, ZN => n148);
   U175 : INV_X1 port map( A => b(17), ZN => n151);
   U176 : INV_X1 port map( A => n152, ZN => o(16));
   U177 : AOI221_X1 port map( B1 => ado_16_port, B2 => n2, C1 => sho_16_port, 
                           C2 => n4, A => n153, ZN => n152);
   U178 : MUX2_X1 port map( A => n154, B => n155, S => a(16), Z => n153);
   U179 : NAND2_X1 port map( A1 => n156, A2 => n10, ZN => n155);
   U180 : MUX2_X1 port map( A => n11, B => n12, S => b(16), Z => n156);
   U181 : NOR2_X1 port map( A1 => n11, A2 => n157, ZN => n154);
   U182 : INV_X1 port map( A => b(16), ZN => n157);
   U183 : INV_X1 port map( A => n158, ZN => o(15));
   U184 : AOI221_X1 port map( B1 => ado_15_port, B2 => n2, C1 => sho_15_port, 
                           C2 => n4, A => n159, ZN => n158);
   U185 : MUX2_X1 port map( A => n160, B => n161, S => a(15), Z => n159);
   U186 : NAND2_X1 port map( A1 => n162, A2 => n10, ZN => n161);
   U187 : MUX2_X1 port map( A => n11, B => n12, S => b(15), Z => n162);
   U188 : NOR2_X1 port map( A1 => n11, A2 => n163, ZN => n160);
   U189 : INV_X1 port map( A => b(15), ZN => n163);
   U190 : INV_X1 port map( A => n164, ZN => o(14));
   U191 : AOI221_X1 port map( B1 => ado_14_port, B2 => n2, C1 => sho_14_port, 
                           C2 => n4, A => n165, ZN => n164);
   U192 : MUX2_X1 port map( A => n166, B => n167, S => a(14), Z => n165);
   U193 : NAND2_X1 port map( A1 => n168, A2 => n10, ZN => n167);
   U194 : MUX2_X1 port map( A => n11, B => n12, S => b(14), Z => n168);
   U195 : NOR2_X1 port map( A1 => n11, A2 => n169, ZN => n166);
   U196 : INV_X1 port map( A => b(14), ZN => n169);
   U197 : INV_X1 port map( A => n170, ZN => o(13));
   U198 : AOI221_X1 port map( B1 => ado_13_port, B2 => n2, C1 => sho_13_port, 
                           C2 => n4, A => n171, ZN => n170);
   U199 : MUX2_X1 port map( A => n172, B => n173, S => a(13), Z => n171);
   U200 : NAND2_X1 port map( A1 => n174, A2 => n10, ZN => n173);
   U201 : MUX2_X1 port map( A => n11, B => n12, S => b(13), Z => n174);
   U202 : NOR2_X1 port map( A1 => n11, A2 => n175, ZN => n172);
   U203 : INV_X1 port map( A => b(13), ZN => n175);
   U204 : INV_X1 port map( A => n176, ZN => o(12));
   U205 : AOI221_X1 port map( B1 => ado_12_port, B2 => n2, C1 => sho_12_port, 
                           C2 => n4, A => n177, ZN => n176);
   U206 : MUX2_X1 port map( A => n178, B => n179, S => a(12), Z => n177);
   U207 : NAND2_X1 port map( A1 => n180, A2 => n10, ZN => n179);
   U208 : MUX2_X1 port map( A => n11, B => n12, S => b(12), Z => n180);
   U209 : NOR2_X1 port map( A1 => n11, A2 => n181, ZN => n178);
   U210 : INV_X1 port map( A => b(12), ZN => n181);
   U211 : INV_X1 port map( A => n182, ZN => o(11));
   U212 : AOI221_X1 port map( B1 => ado_11_port, B2 => n2, C1 => sho_11_port, 
                           C2 => n4, A => n183, ZN => n182);
   U213 : MUX2_X1 port map( A => n184, B => n185, S => a(11), Z => n183);
   U214 : NAND2_X1 port map( A1 => n186, A2 => n10, ZN => n185);
   U215 : MUX2_X1 port map( A => n11, B => n12, S => b(11), Z => n186);
   U216 : NOR2_X1 port map( A1 => n11, A2 => n187, ZN => n184);
   U217 : INV_X1 port map( A => b(11), ZN => n187);
   U218 : INV_X1 port map( A => n188, ZN => o(10));
   U219 : AOI221_X1 port map( B1 => ado_10_port, B2 => n2, C1 => sho_10_port, 
                           C2 => n4, A => n189, ZN => n188);
   U220 : MUX2_X1 port map( A => n190, B => n191, S => a(10), Z => n189);
   U221 : NAND2_X1 port map( A1 => n192, A2 => n10, ZN => n191);
   U222 : MUX2_X1 port map( A => n11, B => n12, S => b(10), Z => n192);
   U223 : NOR2_X1 port map( A1 => n11, A2 => n193, ZN => n190);
   U224 : INV_X1 port map( A => b(10), ZN => n193);
   U225 : INV_X1 port map( A => n194, ZN => o(0));
   U226 : AOI221_X1 port map( B1 => f(4), B2 => n195, C1 => n2, C2 => 
                           ado_0_port, A => n196, ZN => n194);
   U227 : INV_X1 port map( A => n197, ZN => n196);
   U228 : AOI21_X1 port map( B1 => sho_0_port, B2 => n4, A => n198, ZN => n197)
                           ;
   U229 : MUX2_X1 port map( A => n199, B => n200, S => a(0), Z => n198);
   U230 : NAND2_X1 port map( A1 => n201, A2 => n10, ZN => n200);
   U231 : MUX2_X1 port map( A => n11, B => n12, S => b(0), Z => n201);
   U232 : NAND3_X1 port map( A1 => n203, A2 => n204, A3 => f(0), ZN => n12);
   U233 : NOR2_X1 port map( A1 => n11, A2 => n205, ZN => n199);
   U234 : INV_X1 port map( A => b(0), ZN => n205);
   U235 : NOR3_X1 port map( A1 => f(3), A2 => f(4), A3 => f(2), ZN => n203);
   U236 : INV_X1 port map( A => n208, ZN => n195);
   U237 : MUX2_X1 port map( A => n209, B => n210, S => f(3), Z => n208);
   U238 : OAI21_X1 port map( B1 => n211, B2 => n212, A => n206, ZN => n210);
   U239 : MUX2_X1 port map( A => n204, B => n202, S => n213, Z => n212);
   U240 : NOR2_X1 port map( A1 => c_f, A2 => n207, ZN => n211);
   U241 : AOI221_X1 port map( B1 => n214, B2 => n202, C1 => n215, C2 => f(0), A
                           => n216, ZN => n209);
   U242 : AOI211_X1 port map( C1 => n217, C2 => n213, A => n206, B => n207, ZN 
                           => n216);
   U243 : OR2_X1 port map( A1 => f(0), A2 => f(1), ZN => n207);
   U244 : INV_X1 port map( A => f(2), ZN => n206);
   U245 : MUX2_X1 port map( A => n218, B => n219, S => f(1), Z => n215);
   U246 : INV_X1 port map( A => n214, ZN => n219);
   U247 : AND2_X1 port map( A1 => n213, A2 => n214, ZN => n218);
   U248 : NAND2_X1 port map( A1 => n220, A2 => n221, ZN => n213);
   U249 : NOR4_X1 port map( A1 => n222, A2 => n223, A3 => n224, A4 => n225, ZN 
                           => n221);
   U250 : OR4_X1 port map( A1 => ado_24_port, A2 => ado_25_port, A3 => 
                           ado_26_port, A4 => ado_27_port, ZN => n225);
   U251 : OR4_X1 port map( A1 => ado_28_port, A2 => ado_29_port, A3 => 
                           ado_2_port, A4 => ado_30_port, ZN => n224);
   U252 : OR4_X1 port map( A1 => ado_31_port, A2 => ado_3_port, A3 => 
                           ado_4_port, A4 => ado_5_port, ZN => n223);
   U253 : OR4_X1 port map( A1 => ado_6_port, A2 => ado_7_port, A3 => ado_8_port
                           , A4 => ado_9_port, ZN => n222);
   U254 : NOR4_X1 port map( A1 => n226, A2 => n227, A3 => n228, A4 => n229, ZN 
                           => n220);
   U255 : OR4_X1 port map( A1 => ado_0_port, A2 => ado_10_port, A3 => 
                           ado_11_port, A4 => ado_12_port, ZN => n229);
   U256 : OR4_X1 port map( A1 => ado_13_port, A2 => ado_14_port, A3 => 
                           ado_15_port, A4 => ado_16_port, ZN => n228);
   U257 : OR4_X1 port map( A1 => ado_17_port, A2 => ado_18_port, A3 => 
                           ado_19_port, A4 => ado_1_port, ZN => n227);
   U258 : OR4_X1 port map( A1 => ado_20_port, A2 => ado_21_port, A3 => 
                           ado_22_port, A4 => ado_23_port, ZN => n226);
   U259 : NOR2_X1 port map( A1 => n204, A2 => f(0), ZN => n202);
   U260 : INV_X1 port map( A => f(1), ZN => n204);
   U261 : MUX2_X1 port map( A => n217, B => c_f, S => f(2), Z => n214);
   U262 : XOR2_X1 port map( A => n230, B => ado_31_port, Z => n217);
   U263 : OAI21_X1 port map( B1 => ado_31_port, B2 => a(31), A => n231, ZN => 
                           n230);
   U264 : INV_X1 port map( A => n232, ZN => n231);
   U265 : MUX2_X1 port map( A => a(31), B => ado_31_port, S => b_new_31_port, Z
                           => n232);
   U266 : XOR2_X1 port map( A => f(4), B => b(9), Z => b_new_9_port);
   U267 : XOR2_X1 port map( A => f(4), B => b(8), Z => b_new_8_port);
   U268 : XOR2_X1 port map( A => f(4), B => b(7), Z => b_new_7_port);
   U269 : XOR2_X1 port map( A => f(4), B => b(6), Z => b_new_6_port);
   U270 : XOR2_X1 port map( A => f(4), B => b(5), Z => b_new_5_port);
   U271 : XOR2_X1 port map( A => f(4), B => b(4), Z => b_new_4_port);
   U272 : XOR2_X1 port map( A => f(4), B => b(3), Z => b_new_3_port);
   U273 : XOR2_X1 port map( A => b(31), B => f(4), Z => b_new_31_port);
   U274 : XOR2_X1 port map( A => f(4), B => b(30), Z => b_new_30_port);
   U275 : XOR2_X1 port map( A => f(4), B => b(2), Z => b_new_2_port);
   U276 : XOR2_X1 port map( A => f(4), B => b(29), Z => b_new_29_port);
   U277 : XOR2_X1 port map( A => f(4), B => b(28), Z => b_new_28_port);
   U278 : XOR2_X1 port map( A => f(4), B => b(27), Z => b_new_27_port);
   U279 : XOR2_X1 port map( A => f(4), B => b(26), Z => b_new_26_port);
   U280 : XOR2_X1 port map( A => f(4), B => b(25), Z => b_new_25_port);
   U281 : XOR2_X1 port map( A => f(4), B => b(24), Z => b_new_24_port);
   U282 : XOR2_X1 port map( A => f(4), B => b(23), Z => b_new_23_port);
   U283 : XOR2_X1 port map( A => f(4), B => b(22), Z => b_new_22_port);
   U284 : XOR2_X1 port map( A => f(4), B => b(21), Z => b_new_21_port);
   U285 : XOR2_X1 port map( A => f(4), B => b(20), Z => b_new_20_port);
   U286 : XOR2_X1 port map( A => f(4), B => b(1), Z => b_new_1_port);
   U287 : XOR2_X1 port map( A => f(4), B => b(19), Z => b_new_19_port);
   U288 : XOR2_X1 port map( A => f(4), B => b(18), Z => b_new_18_port);
   U289 : XOR2_X1 port map( A => f(4), B => b(17), Z => b_new_17_port);
   U290 : XOR2_X1 port map( A => f(4), B => b(16), Z => b_new_16_port);
   U291 : XOR2_X1 port map( A => f(4), B => b(15), Z => b_new_15_port);
   U292 : XOR2_X1 port map( A => f(4), B => b(14), Z => b_new_14_port);
   U293 : XOR2_X1 port map( A => f(4), B => b(13), Z => b_new_13_port);
   U294 : XOR2_X1 port map( A => f(4), B => b(12), Z => b_new_12_port);
   U295 : XOR2_X1 port map( A => f(4), B => b(11), Z => b_new_11_port);
   U296 : XOR2_X1 port map( A => f(4), B => b(10), Z => b_new_10_port);
   U297 : XOR2_X1 port map( A => f(4), B => b(0), Z => b_new_0_port);

end SYN_alu_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE5_0 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 0); 
         dout : out std_logic_vector (4 downto 0));

end Reg_DATA_SIZE5_0;

architecture SYN_reg_arch of Reg_DATA_SIZE5_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal dout_4_port, dout_3_port, dout_2_port, dout_1_port, dout_0_port, n11,
      n12, n13, n14, n15, net108611, net108612, net108613, net108614, net108615
      : std_logic;

begin
   dout <= ( dout_4_port, dout_3_port, dout_2_port, dout_1_port, dout_0_port );
   
   dout_reg_4_inst : DFFR_X1 port map( D => n15, CK => clk, RN => rst, Q => 
                           dout_4_port, QN => net108615);
   dout_reg_3_inst : DFFR_X1 port map( D => n14, CK => clk, RN => rst, Q => 
                           dout_3_port, QN => net108614);
   dout_reg_2_inst : DFFR_X1 port map( D => n13, CK => clk, RN => rst, Q => 
                           dout_2_port, QN => net108613);
   dout_reg_1_inst : DFFR_X1 port map( D => n12, CK => clk, RN => rst, Q => 
                           dout_1_port, QN => net108612);
   dout_reg_0_inst : DFFR_X1 port map( D => n11, CK => clk, RN => rst, Q => 
                           dout_0_port, QN => net108611);
   U2 : MUX2_X1 port map( A => dout_4_port, B => din(4), S => en, Z => n15);
   U3 : MUX2_X1 port map( A => dout_3_port, B => din(3), S => en, Z => n14);
   U4 : MUX2_X1 port map( A => dout_2_port, B => din(2), S => en, Z => n13);
   U5 : MUX2_X1 port map( A => dout_1_port, B => din(1), S => en, Z => n12);
   U6 : MUX2_X1 port map( A => dout_0_port, B => din(0), S => en, Z => n11);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_0 is

   port( reg_c, reg_f, reg_ff : in std_logic_vector (31 downto 0);  addr_c, 
         addr_f, addr_ff : in std_logic_vector (4 downto 0);  valid_f, valid_ff
         , dirty_f, dirty_ff, en : in std_logic;  output : out std_logic_vector
         (31 downto 0);  match_dirty_f, match_dirty_ff : out std_logic);

end FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_0;

architecture SYN_fwd_mux_2_arch of FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X4
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X2
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N91, N92,
      N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105, 
      N106, N107, N108, N109, N110, N111, N112, n1, n2, n3, n4, n5, n6, n7, n8,
      n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
      n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38
      , n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, 
      n53, n54, n55 : std_logic;

begin
   
   match_dirty_ff_reg : DLH_X1 port map( G => en, D => N111, Q => 
                           match_dirty_ff);
   output_reg_31_inst : DLH_X1 port map( G => en, D => N110, Q => output(31));
   output_reg_30_inst : DLH_X1 port map( G => en, D => N109, Q => output(30));
   output_reg_29_inst : DLH_X1 port map( G => en, D => N108, Q => output(29));
   output_reg_28_inst : DLH_X1 port map( G => en, D => N107, Q => output(28));
   output_reg_27_inst : DLH_X1 port map( G => en, D => N106, Q => output(27));
   output_reg_26_inst : DLH_X1 port map( G => en, D => N105, Q => output(26));
   output_reg_25_inst : DLH_X1 port map( G => en, D => N104, Q => output(25));
   output_reg_24_inst : DLH_X1 port map( G => en, D => N103, Q => output(24));
   output_reg_23_inst : DLH_X1 port map( G => en, D => N102, Q => output(23));
   output_reg_22_inst : DLH_X1 port map( G => en, D => N101, Q => output(22));
   output_reg_21_inst : DLH_X1 port map( G => en, D => N100, Q => output(21));
   output_reg_20_inst : DLH_X1 port map( G => en, D => N99, Q => output(20));
   output_reg_19_inst : DLH_X1 port map( G => en, D => N98, Q => output(19));
   output_reg_18_inst : DLH_X1 port map( G => en, D => N97, Q => output(18));
   output_reg_17_inst : DLH_X1 port map( G => en, D => N96, Q => output(17));
   output_reg_16_inst : DLH_X1 port map( G => en, D => N95, Q => output(16));
   output_reg_15_inst : DLH_X1 port map( G => en, D => N94, Q => output(15));
   output_reg_14_inst : DLH_X1 port map( G => en, D => N93, Q => output(14));
   output_reg_13_inst : DLH_X1 port map( G => en, D => N92, Q => output(13));
   output_reg_12_inst : DLH_X1 port map( G => en, D => N91, Q => output(12));
   output_reg_11_inst : DLH_X1 port map( G => en, D => N90, Q => output(11));
   output_reg_10_inst : DLH_X1 port map( G => en, D => N89, Q => output(10));
   output_reg_9_inst : DLH_X1 port map( G => en, D => N88, Q => output(9));
   output_reg_8_inst : DLH_X1 port map( G => en, D => N87, Q => output(8));
   output_reg_7_inst : DLH_X1 port map( G => en, D => N86, Q => output(7));
   output_reg_6_inst : DLH_X1 port map( G => en, D => N85, Q => output(6));
   output_reg_5_inst : DLH_X1 port map( G => en, D => N84, Q => output(5));
   output_reg_4_inst : DLH_X1 port map( G => en, D => N83, Q => output(4));
   output_reg_3_inst : DLH_X1 port map( G => en, D => N82, Q => output(3));
   output_reg_2_inst : DLH_X1 port map( G => en, D => N81, Q => output(2));
   output_reg_1_inst : DLH_X1 port map( G => en, D => N80, Q => output(1));
   output_reg_0_inst : DLH_X1 port map( G => en, D => N79, Q => output(0));
   match_dirty_f_reg : DLH_X2 port map( G => en, D => N112, Q => match_dirty_f)
                           ;
   U2 : OAI21_X4 port map( B1 => n38, B2 => n39, A => n36, ZN => n2);
   U3 : AND3_X2 port map( A1 => n36, A2 => n37, A3 => n38, ZN => n4);
   U4 : AND2_X2 port map( A1 => n39, A2 => n36, ZN => n3);
   U5 : INV_X1 port map( A => n1, ZN => N99);
   U6 : AOI222_X1 port map( A1 => reg_c(20), A2 => n2, B1 => reg_f(20), B2 => 
                           n3, C1 => reg_ff(20), C2 => n4, ZN => n1);
   U7 : INV_X1 port map( A => n5, ZN => N98);
   U8 : AOI222_X1 port map( A1 => reg_c(19), A2 => n2, B1 => reg_f(19), B2 => 
                           n3, C1 => reg_ff(19), C2 => n4, ZN => n5);
   U9 : INV_X1 port map( A => n6, ZN => N97);
   U10 : AOI222_X1 port map( A1 => reg_c(18), A2 => n2, B1 => reg_f(18), B2 => 
                           n3, C1 => reg_ff(18), C2 => n4, ZN => n6);
   U11 : INV_X1 port map( A => n7, ZN => N96);
   U12 : AOI222_X1 port map( A1 => reg_c(17), A2 => n2, B1 => reg_f(17), B2 => 
                           n3, C1 => reg_ff(17), C2 => n4, ZN => n7);
   U13 : INV_X1 port map( A => n8, ZN => N95);
   U14 : AOI222_X1 port map( A1 => reg_c(16), A2 => n2, B1 => reg_f(16), B2 => 
                           n3, C1 => reg_ff(16), C2 => n4, ZN => n8);
   U15 : INV_X1 port map( A => n9, ZN => N94);
   U16 : AOI222_X1 port map( A1 => reg_c(15), A2 => n2, B1 => reg_f(15), B2 => 
                           n3, C1 => reg_ff(15), C2 => n4, ZN => n9);
   U17 : INV_X1 port map( A => n10, ZN => N93);
   U18 : AOI222_X1 port map( A1 => reg_c(14), A2 => n2, B1 => reg_f(14), B2 => 
                           n3, C1 => reg_ff(14), C2 => n4, ZN => n10);
   U19 : INV_X1 port map( A => n11, ZN => N92);
   U20 : AOI222_X1 port map( A1 => reg_c(13), A2 => n2, B1 => reg_f(13), B2 => 
                           n3, C1 => reg_ff(13), C2 => n4, ZN => n11);
   U21 : INV_X1 port map( A => n12, ZN => N91);
   U22 : AOI222_X1 port map( A1 => reg_c(12), A2 => n2, B1 => reg_f(12), B2 => 
                           n3, C1 => reg_ff(12), C2 => n4, ZN => n12);
   U23 : INV_X1 port map( A => n13, ZN => N90);
   U24 : AOI222_X1 port map( A1 => reg_c(11), A2 => n2, B1 => reg_f(11), B2 => 
                           n3, C1 => reg_ff(11), C2 => n4, ZN => n13);
   U25 : INV_X1 port map( A => n14, ZN => N89);
   U26 : AOI222_X1 port map( A1 => reg_c(10), A2 => n2, B1 => reg_f(10), B2 => 
                           n3, C1 => reg_ff(10), C2 => n4, ZN => n14);
   U27 : INV_X1 port map( A => n15, ZN => N88);
   U28 : AOI222_X1 port map( A1 => reg_c(9), A2 => n2, B1 => reg_f(9), B2 => n3
                           , C1 => reg_ff(9), C2 => n4, ZN => n15);
   U29 : INV_X1 port map( A => n16, ZN => N87);
   U30 : AOI222_X1 port map( A1 => reg_c(8), A2 => n2, B1 => reg_f(8), B2 => n3
                           , C1 => reg_ff(8), C2 => n4, ZN => n16);
   U31 : INV_X1 port map( A => n17, ZN => N86);
   U32 : AOI222_X1 port map( A1 => reg_c(7), A2 => n2, B1 => reg_f(7), B2 => n3
                           , C1 => reg_ff(7), C2 => n4, ZN => n17);
   U33 : INV_X1 port map( A => n18, ZN => N85);
   U34 : AOI222_X1 port map( A1 => reg_c(6), A2 => n2, B1 => reg_f(6), B2 => n3
                           , C1 => reg_ff(6), C2 => n4, ZN => n18);
   U35 : INV_X1 port map( A => n19, ZN => N84);
   U36 : AOI222_X1 port map( A1 => reg_c(5), A2 => n2, B1 => reg_f(5), B2 => n3
                           , C1 => reg_ff(5), C2 => n4, ZN => n19);
   U37 : INV_X1 port map( A => n20, ZN => N83);
   U38 : AOI222_X1 port map( A1 => reg_c(4), A2 => n2, B1 => reg_f(4), B2 => n3
                           , C1 => reg_ff(4), C2 => n4, ZN => n20);
   U39 : INV_X1 port map( A => n21, ZN => N82);
   U40 : AOI222_X1 port map( A1 => reg_c(3), A2 => n2, B1 => reg_f(3), B2 => n3
                           , C1 => reg_ff(3), C2 => n4, ZN => n21);
   U41 : INV_X1 port map( A => n22, ZN => N81);
   U42 : AOI222_X1 port map( A1 => reg_c(2), A2 => n2, B1 => reg_f(2), B2 => n3
                           , C1 => reg_ff(2), C2 => n4, ZN => n22);
   U43 : INV_X1 port map( A => n23, ZN => N80);
   U44 : AOI222_X1 port map( A1 => reg_c(1), A2 => n2, B1 => reg_f(1), B2 => n3
                           , C1 => reg_ff(1), C2 => n4, ZN => n23);
   U45 : INV_X1 port map( A => n24, ZN => N79);
   U46 : AOI222_X1 port map( A1 => reg_c(0), A2 => n2, B1 => reg_f(0), B2 => n3
                           , C1 => reg_ff(0), C2 => n4, ZN => n24);
   U47 : AND2_X1 port map( A1 => dirty_f, A2 => n3, ZN => N112);
   U48 : AND2_X1 port map( A1 => dirty_ff, A2 => n4, ZN => N111);
   U49 : INV_X1 port map( A => n25, ZN => N110);
   U50 : AOI222_X1 port map( A1 => reg_c(31), A2 => n2, B1 => reg_f(31), B2 => 
                           n3, C1 => reg_ff(31), C2 => n4, ZN => n25);
   U51 : INV_X1 port map( A => n26, ZN => N109);
   U52 : AOI222_X1 port map( A1 => reg_c(30), A2 => n2, B1 => reg_f(30), B2 => 
                           n3, C1 => reg_ff(30), C2 => n4, ZN => n26);
   U53 : INV_X1 port map( A => n27, ZN => N108);
   U54 : AOI222_X1 port map( A1 => reg_c(29), A2 => n2, B1 => reg_f(29), B2 => 
                           n3, C1 => reg_ff(29), C2 => n4, ZN => n27);
   U55 : INV_X1 port map( A => n28, ZN => N107);
   U56 : AOI222_X1 port map( A1 => reg_c(28), A2 => n2, B1 => reg_f(28), B2 => 
                           n3, C1 => reg_ff(28), C2 => n4, ZN => n28);
   U57 : INV_X1 port map( A => n29, ZN => N106);
   U58 : AOI222_X1 port map( A1 => reg_c(27), A2 => n2, B1 => reg_f(27), B2 => 
                           n3, C1 => reg_ff(27), C2 => n4, ZN => n29);
   U59 : INV_X1 port map( A => n30, ZN => N105);
   U60 : AOI222_X1 port map( A1 => reg_c(26), A2 => n2, B1 => reg_f(26), B2 => 
                           n3, C1 => reg_ff(26), C2 => n4, ZN => n30);
   U61 : INV_X1 port map( A => n31, ZN => N104);
   U62 : AOI222_X1 port map( A1 => reg_c(25), A2 => n2, B1 => reg_f(25), B2 => 
                           n3, C1 => reg_ff(25), C2 => n4, ZN => n31);
   U63 : INV_X1 port map( A => n32, ZN => N103);
   U64 : AOI222_X1 port map( A1 => reg_c(24), A2 => n2, B1 => reg_f(24), B2 => 
                           n3, C1 => reg_ff(24), C2 => n4, ZN => n32);
   U65 : INV_X1 port map( A => n33, ZN => N102);
   U66 : AOI222_X1 port map( A1 => reg_c(23), A2 => n2, B1 => reg_f(23), B2 => 
                           n3, C1 => reg_ff(23), C2 => n4, ZN => n33);
   U67 : INV_X1 port map( A => n34, ZN => N101);
   U68 : AOI222_X1 port map( A1 => reg_c(22), A2 => n2, B1 => reg_f(22), B2 => 
                           n3, C1 => reg_ff(22), C2 => n4, ZN => n34);
   U69 : INV_X1 port map( A => n35, ZN => N100);
   U70 : AOI222_X1 port map( A1 => reg_c(21), A2 => n2, B1 => reg_f(21), B2 => 
                           n3, C1 => reg_ff(21), C2 => n4, ZN => n35);
   U71 : NAND4_X1 port map( A1 => n40, A2 => n41, A3 => n42, A4 => n43, ZN => 
                           n36);
   U72 : NOR2_X1 port map( A1 => addr_c(1), A2 => addr_c(0), ZN => n43);
   U73 : INV_X1 port map( A => addr_c(4), ZN => n41);
   U74 : INV_X1 port map( A => n37, ZN => n39);
   U75 : NAND4_X1 port map( A1 => n44, A2 => valid_f, A3 => n45, A4 => n46, ZN 
                           => n37);
   U76 : NOR3_X1 port map( A1 => n47, A2 => n48, A3 => n49, ZN => n46);
   U77 : XOR2_X1 port map( A => addr_f(2), B => addr_c(2), Z => n49);
   U78 : XOR2_X1 port map( A => addr_f(4), B => addr_c(4), Z => n48);
   U79 : XOR2_X1 port map( A => addr_f(3), B => addr_c(3), Z => n47);
   U80 : XNOR2_X1 port map( A => addr_c(0), B => addr_f(0), ZN => n45);
   U81 : XNOR2_X1 port map( A => addr_c(1), B => addr_f(1), ZN => n44);
   U82 : AND4_X1 port map( A1 => n50, A2 => valid_ff, A3 => n51, A4 => n52, ZN 
                           => n38);
   U83 : NOR3_X1 port map( A1 => n53, A2 => n54, A3 => n55, ZN => n52);
   U84 : XOR2_X1 port map( A => addr_ff(0), B => addr_c(0), Z => n55);
   U85 : XOR2_X1 port map( A => addr_ff(1), B => addr_c(1), Z => n54);
   U86 : XOR2_X1 port map( A => addr_ff(4), B => addr_c(4), Z => n53);
   U87 : XOR2_X1 port map( A => n40, B => addr_ff(3), Z => n51);
   U88 : INV_X1 port map( A => addr_c(3), ZN => n40);
   U89 : XOR2_X1 port map( A => n42, B => addr_ff(2), Z => n50);
   U90 : INV_X1 port map( A => addr_c(2), ZN => n42);

end SYN_fwd_mux_2_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity RegisterFile_DATA_SIZE32_REG_NUM32 is

   port( clk, rst, en, rd1_en, rd2_en, wr_en, link_en : in std_logic;  rd1_addr
         , rd2_addr, wr_addr : in std_logic_vector (4 downto 0);  d_out1, 
         d_out2 : out std_logic_vector (31 downto 0);  d_in, d_link : in 
         std_logic_vector (31 downto 0));

end RegisterFile_DATA_SIZE32_REG_NUM32;

architecture SYN_register_file_arch of RegisterFile_DATA_SIZE32_REG_NUM32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal d_out1_31_port, d_out1_30_port, d_out1_29_port, d_out1_28_port, 
      d_out1_27_port, d_out1_26_port, d_out1_25_port, d_out1_24_port, 
      d_out1_23_port, d_out1_22_port, d_out1_21_port, d_out1_20_port, 
      d_out1_19_port, d_out1_18_port, d_out1_17_port, d_out1_16_port, 
      d_out1_15_port, d_out1_14_port, d_out1_13_port, d_out1_12_port, 
      d_out1_11_port, d_out1_10_port, d_out1_9_port, d_out1_8_port, 
      d_out1_7_port, d_out1_6_port, d_out1_5_port, d_out1_4_port, d_out1_3_port
      , d_out1_2_port, d_out1_1_port, d_out1_0_port, d_out2_31_port, 
      d_out2_30_port, d_out2_29_port, d_out2_28_port, d_out2_27_port, 
      d_out2_26_port, d_out2_25_port, d_out2_24_port, d_out2_23_port, 
      d_out2_22_port, d_out2_21_port, d_out2_20_port, d_out2_19_port, 
      d_out2_18_port, d_out2_17_port, d_out2_16_port, d_out2_15_port, 
      d_out2_14_port, d_out2_13_port, d_out2_12_port, d_out2_11_port, 
      d_out2_10_port, d_out2_9_port, d_out2_8_port, d_out2_7_port, 
      d_out2_6_port, d_out2_5_port, d_out2_4_port, d_out2_3_port, d_out2_2_port
      , d_out2_1_port, d_out2_0_port, registers_1_31_port, registers_1_30_port,
      registers_1_29_port, registers_1_28_port, registers_1_27_port, 
      registers_1_26_port, registers_1_25_port, registers_1_24_port, 
      registers_1_23_port, registers_1_22_port, registers_1_21_port, 
      registers_1_20_port, registers_1_19_port, registers_1_18_port, 
      registers_1_17_port, registers_1_16_port, registers_1_15_port, 
      registers_1_14_port, registers_1_13_port, registers_1_12_port, 
      registers_1_11_port, registers_1_10_port, registers_1_9_port, 
      registers_1_8_port, registers_1_7_port, registers_1_6_port, 
      registers_1_5_port, registers_1_4_port, registers_1_3_port, 
      registers_1_2_port, registers_1_1_port, registers_1_0_port, 
      registers_2_31_port, registers_2_30_port, registers_2_29_port, 
      registers_2_28_port, registers_2_27_port, registers_2_26_port, 
      registers_2_25_port, registers_2_24_port, registers_2_23_port, 
      registers_2_22_port, registers_2_21_port, registers_2_20_port, 
      registers_2_19_port, registers_2_18_port, registers_2_17_port, 
      registers_2_16_port, registers_2_15_port, registers_2_14_port, 
      registers_2_13_port, registers_2_12_port, registers_2_11_port, 
      registers_2_10_port, registers_2_9_port, registers_2_8_port, 
      registers_2_7_port, registers_2_6_port, registers_2_5_port, 
      registers_2_4_port, registers_2_3_port, registers_2_2_port, 
      registers_2_1_port, registers_2_0_port, registers_3_31_port, 
      registers_3_30_port, registers_3_29_port, registers_3_28_port, 
      registers_3_27_port, registers_3_26_port, registers_3_25_port, 
      registers_3_24_port, registers_3_23_port, registers_3_22_port, 
      registers_3_21_port, registers_3_20_port, registers_3_19_port, 
      registers_3_18_port, registers_3_17_port, registers_3_16_port, 
      registers_3_15_port, registers_3_14_port, registers_3_13_port, 
      registers_3_12_port, registers_3_11_port, registers_3_10_port, 
      registers_3_9_port, registers_3_8_port, registers_3_7_port, 
      registers_3_6_port, registers_3_5_port, registers_3_4_port, 
      registers_3_3_port, registers_3_2_port, registers_3_1_port, 
      registers_3_0_port, registers_4_31_port, registers_4_30_port, 
      registers_4_29_port, registers_4_28_port, registers_4_27_port, 
      registers_4_26_port, registers_4_25_port, registers_4_24_port, 
      registers_4_23_port, registers_4_22_port, registers_4_21_port, 
      registers_4_20_port, registers_4_19_port, registers_4_18_port, 
      registers_4_17_port, registers_4_16_port, registers_4_15_port, 
      registers_4_14_port, registers_4_13_port, registers_4_12_port, 
      registers_4_11_port, registers_4_10_port, registers_4_9_port, 
      registers_4_8_port, registers_4_7_port, registers_4_6_port, 
      registers_4_5_port, registers_4_4_port, registers_4_3_port, 
      registers_4_2_port, registers_4_1_port, registers_4_0_port, 
      registers_5_31_port, registers_5_30_port, registers_5_29_port, 
      registers_5_28_port, registers_5_27_port, registers_5_26_port, 
      registers_5_25_port, registers_5_24_port, registers_5_23_port, 
      registers_5_22_port, registers_5_21_port, registers_5_20_port, 
      registers_5_19_port, registers_5_18_port, registers_5_17_port, 
      registers_5_16_port, registers_5_15_port, registers_5_14_port, 
      registers_5_13_port, registers_5_12_port, registers_5_11_port, 
      registers_5_10_port, registers_5_9_port, registers_5_8_port, 
      registers_5_7_port, registers_5_6_port, registers_5_5_port, 
      registers_5_4_port, registers_5_3_port, registers_5_2_port, 
      registers_5_1_port, registers_5_0_port, registers_6_31_port, 
      registers_6_30_port, registers_6_29_port, registers_6_28_port, 
      registers_6_27_port, registers_6_26_port, registers_6_25_port, 
      registers_6_24_port, registers_6_23_port, registers_6_22_port, 
      registers_6_21_port, registers_6_20_port, registers_6_19_port, 
      registers_6_18_port, registers_6_17_port, registers_6_16_port, 
      registers_6_15_port, registers_6_14_port, registers_6_13_port, 
      registers_6_12_port, registers_6_11_port, registers_6_10_port, 
      registers_6_9_port, registers_6_8_port, registers_6_7_port, 
      registers_6_6_port, registers_6_5_port, registers_6_4_port, 
      registers_6_3_port, registers_6_2_port, registers_6_1_port, 
      registers_6_0_port, registers_7_31_port, registers_7_30_port, 
      registers_7_29_port, registers_7_28_port, registers_7_27_port, 
      registers_7_26_port, registers_7_25_port, registers_7_24_port, 
      registers_7_23_port, registers_7_22_port, registers_7_21_port, 
      registers_7_20_port, registers_7_19_port, registers_7_18_port, 
      registers_7_17_port, registers_7_16_port, registers_7_15_port, 
      registers_7_14_port, registers_7_13_port, registers_7_12_port, 
      registers_7_11_port, registers_7_10_port, registers_7_9_port, 
      registers_7_8_port, registers_7_7_port, registers_7_6_port, 
      registers_7_5_port, registers_7_4_port, registers_7_3_port, 
      registers_7_2_port, registers_7_1_port, registers_7_0_port, 
      registers_8_31_port, registers_8_30_port, registers_8_29_port, 
      registers_8_28_port, registers_8_27_port, registers_8_26_port, 
      registers_8_25_port, registers_8_24_port, registers_8_23_port, 
      registers_8_22_port, registers_8_21_port, registers_8_20_port, 
      registers_8_19_port, registers_8_18_port, registers_8_17_port, 
      registers_8_16_port, registers_8_15_port, registers_8_14_port, 
      registers_8_13_port, registers_8_12_port, registers_8_11_port, 
      registers_8_10_port, registers_8_9_port, registers_8_8_port, 
      registers_8_7_port, registers_8_6_port, registers_8_5_port, 
      registers_8_4_port, registers_8_3_port, registers_8_2_port, 
      registers_8_1_port, registers_8_0_port, registers_9_31_port, 
      registers_9_30_port, registers_9_29_port, registers_9_28_port, 
      registers_9_27_port, registers_9_26_port, registers_9_25_port, 
      registers_9_24_port, registers_9_23_port, registers_9_22_port, 
      registers_9_21_port, registers_9_20_port, registers_9_19_port, 
      registers_9_18_port, registers_9_17_port, registers_9_16_port, 
      registers_9_15_port, registers_9_14_port, registers_9_13_port, 
      registers_9_12_port, registers_9_11_port, registers_9_10_port, 
      registers_9_9_port, registers_9_8_port, registers_9_7_port, 
      registers_9_6_port, registers_9_5_port, registers_9_4_port, 
      registers_9_3_port, registers_9_2_port, registers_9_1_port, 
      registers_9_0_port, registers_10_31_port, registers_10_30_port, 
      registers_10_29_port, registers_10_28_port, registers_10_27_port, 
      registers_10_26_port, registers_10_25_port, registers_10_24_port, 
      registers_10_23_port, registers_10_22_port, registers_10_21_port, 
      registers_10_20_port, registers_10_19_port, registers_10_18_port, 
      registers_10_17_port, registers_10_16_port, registers_10_15_port, 
      registers_10_14_port, registers_10_13_port, registers_10_12_port, 
      registers_10_11_port, registers_10_10_port, registers_10_9_port, 
      registers_10_8_port, registers_10_7_port, registers_10_6_port, 
      registers_10_5_port, registers_10_4_port, registers_10_3_port, 
      registers_10_2_port, registers_10_1_port, registers_10_0_port, 
      registers_11_31_port, registers_11_30_port, registers_11_29_port, 
      registers_11_28_port, registers_11_27_port, registers_11_26_port, 
      registers_11_25_port, registers_11_24_port, registers_11_23_port, 
      registers_11_22_port, registers_11_21_port, registers_11_20_port, 
      registers_11_19_port, registers_11_18_port, registers_11_17_port, 
      registers_11_16_port, registers_11_15_port, registers_11_14_port, 
      registers_11_13_port, registers_11_12_port, registers_11_11_port, 
      registers_11_10_port, registers_11_9_port, registers_11_8_port, 
      registers_11_7_port, registers_11_6_port, registers_11_5_port, 
      registers_11_4_port, registers_11_3_port, registers_11_2_port, 
      registers_11_1_port, registers_11_0_port, registers_12_31_port, 
      registers_12_30_port, registers_12_29_port, registers_12_28_port, 
      registers_12_27_port, registers_12_26_port, registers_12_25_port, 
      registers_12_24_port, registers_12_23_port, registers_12_22_port, 
      registers_12_21_port, registers_12_20_port, registers_12_19_port, 
      registers_12_18_port, registers_12_17_port, registers_12_16_port, 
      registers_12_15_port, registers_12_14_port, registers_12_13_port, 
      registers_12_12_port, registers_12_11_port, registers_12_10_port, 
      registers_12_9_port, registers_12_8_port, registers_12_7_port, 
      registers_12_6_port, registers_12_5_port, registers_12_4_port, 
      registers_12_3_port, registers_12_2_port, registers_12_1_port, 
      registers_12_0_port, registers_13_31_port, registers_13_30_port, 
      registers_13_29_port, registers_13_28_port, registers_13_27_port, 
      registers_13_26_port, registers_13_25_port, registers_13_24_port, 
      registers_13_23_port, registers_13_22_port, registers_13_21_port, 
      registers_13_20_port, registers_13_19_port, registers_13_18_port, 
      registers_13_17_port, registers_13_16_port, registers_13_15_port, 
      registers_13_14_port, registers_13_13_port, registers_13_12_port, 
      registers_13_11_port, registers_13_10_port, registers_13_9_port, 
      registers_13_8_port, registers_13_7_port, registers_13_6_port, 
      registers_13_5_port, registers_13_4_port, registers_13_3_port, 
      registers_13_2_port, registers_13_1_port, registers_13_0_port, 
      registers_14_31_port, registers_14_30_port, registers_14_29_port, 
      registers_14_28_port, registers_14_27_port, registers_14_26_port, 
      registers_14_25_port, registers_14_24_port, registers_14_23_port, 
      registers_14_22_port, registers_14_21_port, registers_14_20_port, 
      registers_14_19_port, registers_14_18_port, registers_14_17_port, 
      registers_14_16_port, registers_14_15_port, registers_14_14_port, 
      registers_14_13_port, registers_14_12_port, registers_14_11_port, 
      registers_14_10_port, registers_14_9_port, registers_14_8_port, 
      registers_14_7_port, registers_14_6_port, registers_14_5_port, 
      registers_14_4_port, registers_14_3_port, registers_14_2_port, 
      registers_14_1_port, registers_14_0_port, registers_15_31_port, 
      registers_15_30_port, registers_15_29_port, registers_15_28_port, 
      registers_15_27_port, registers_15_26_port, registers_15_25_port, 
      registers_15_24_port, registers_15_23_port, registers_15_22_port, 
      registers_15_21_port, registers_15_20_port, registers_15_19_port, 
      registers_15_18_port, registers_15_17_port, registers_15_16_port, 
      registers_15_15_port, registers_15_14_port, registers_15_13_port, 
      registers_15_12_port, registers_15_11_port, registers_15_10_port, 
      registers_15_9_port, registers_15_8_port, registers_15_7_port, 
      registers_15_6_port, registers_15_5_port, registers_15_4_port, 
      registers_15_3_port, registers_15_2_port, registers_15_1_port, 
      registers_15_0_port, registers_16_31_port, registers_16_30_port, 
      registers_16_29_port, registers_16_28_port, registers_16_27_port, 
      registers_16_26_port, registers_16_25_port, registers_16_24_port, 
      registers_16_23_port, registers_16_22_port, registers_16_21_port, 
      registers_16_20_port, registers_16_19_port, registers_16_18_port, 
      registers_16_17_port, registers_16_16_port, registers_16_15_port, 
      registers_16_14_port, registers_16_13_port, registers_16_12_port, 
      registers_16_11_port, registers_16_10_port, registers_16_9_port, 
      registers_16_8_port, registers_16_7_port, registers_16_6_port, 
      registers_16_5_port, registers_16_4_port, registers_16_3_port, 
      registers_16_2_port, registers_16_1_port, registers_16_0_port, 
      registers_17_31_port, registers_17_30_port, registers_17_29_port, 
      registers_17_28_port, registers_17_27_port, registers_17_26_port, 
      registers_17_25_port, registers_17_24_port, registers_17_23_port, 
      registers_17_22_port, registers_17_21_port, registers_17_20_port, 
      registers_17_19_port, registers_17_18_port, registers_17_17_port, 
      registers_17_16_port, registers_17_15_port, registers_17_14_port, 
      registers_17_13_port, registers_17_12_port, registers_17_11_port, 
      registers_17_10_port, registers_17_9_port, registers_17_8_port, 
      registers_17_7_port, registers_17_6_port, registers_17_5_port, 
      registers_17_4_port, registers_17_3_port, registers_17_2_port, 
      registers_17_1_port, registers_17_0_port, registers_18_31_port, 
      registers_18_30_port, registers_18_29_port, registers_18_28_port, 
      registers_18_27_port, registers_18_26_port, registers_18_25_port, 
      registers_18_24_port, registers_18_23_port, registers_18_22_port, 
      registers_18_21_port, registers_18_20_port, registers_18_19_port, 
      registers_18_18_port, registers_18_17_port, registers_18_16_port, 
      registers_18_15_port, registers_18_14_port, registers_18_13_port, 
      registers_18_12_port, registers_18_11_port, registers_18_10_port, 
      registers_18_9_port, registers_18_8_port, registers_18_7_port, 
      registers_18_6_port, registers_18_5_port, registers_18_4_port, 
      registers_18_3_port, registers_18_2_port, registers_18_1_port, 
      registers_18_0_port, registers_19_31_port, registers_19_30_port, 
      registers_19_29_port, registers_19_28_port, registers_19_27_port, 
      registers_19_26_port, registers_19_25_port, registers_19_24_port, 
      registers_19_23_port, registers_19_22_port, registers_19_21_port, 
      registers_19_20_port, registers_19_19_port, registers_19_18_port, 
      registers_19_17_port, registers_19_16_port, registers_19_15_port, 
      registers_19_14_port, registers_19_13_port, registers_19_12_port, 
      registers_19_11_port, registers_19_10_port, registers_19_9_port, 
      registers_19_8_port, registers_19_7_port, registers_19_6_port, 
      registers_19_5_port, registers_19_4_port, registers_19_3_port, 
      registers_19_2_port, registers_19_1_port, registers_19_0_port, 
      registers_20_31_port, registers_20_30_port, registers_20_29_port, 
      registers_20_28_port, registers_20_27_port, registers_20_26_port, 
      registers_20_25_port, registers_20_24_port, registers_20_23_port, 
      registers_20_22_port, registers_20_21_port, registers_20_20_port, 
      registers_20_19_port, registers_20_18_port, registers_20_17_port, 
      registers_20_16_port, registers_20_15_port, registers_20_14_port, 
      registers_20_13_port, registers_20_12_port, registers_20_11_port, 
      registers_20_10_port, registers_20_9_port, registers_20_8_port, 
      registers_20_7_port, registers_20_6_port, registers_20_5_port, 
      registers_20_4_port, registers_20_3_port, registers_20_2_port, 
      registers_20_1_port, registers_20_0_port, registers_21_31_port, 
      registers_21_30_port, registers_21_29_port, registers_21_28_port, 
      registers_21_27_port, registers_21_26_port, registers_21_25_port, 
      registers_21_24_port, registers_21_23_port, registers_21_22_port, 
      registers_21_21_port, registers_21_20_port, registers_21_19_port, 
      registers_21_18_port, registers_21_17_port, registers_21_16_port, 
      registers_21_15_port, registers_21_14_port, registers_21_13_port, 
      registers_21_12_port, registers_21_11_port, registers_21_10_port, 
      registers_21_9_port, registers_21_8_port, registers_21_7_port, 
      registers_21_6_port, registers_21_5_port, registers_21_4_port, 
      registers_21_3_port, registers_21_2_port, registers_21_1_port, 
      registers_21_0_port, registers_22_31_port, registers_22_30_port, 
      registers_22_29_port, registers_22_28_port, registers_22_27_port, 
      registers_22_26_port, registers_22_25_port, registers_22_24_port, 
      registers_22_23_port, registers_22_22_port, registers_22_21_port, 
      registers_22_20_port, registers_22_19_port, registers_22_18_port, 
      registers_22_17_port, registers_22_16_port, registers_22_15_port, 
      registers_22_14_port, registers_22_13_port, registers_22_12_port, 
      registers_22_11_port, registers_22_10_port, registers_22_9_port, 
      registers_22_8_port, registers_22_7_port, registers_22_6_port, 
      registers_22_5_port, registers_22_4_port, registers_22_3_port, 
      registers_22_2_port, registers_22_1_port, registers_22_0_port, 
      registers_23_31_port, registers_23_30_port, registers_23_29_port, 
      registers_23_28_port, registers_23_27_port, registers_23_26_port, 
      registers_23_25_port, registers_23_24_port, registers_23_23_port, 
      registers_23_22_port, registers_23_21_port, registers_23_20_port, 
      registers_23_19_port, registers_23_18_port, registers_23_17_port, 
      registers_23_16_port, registers_23_15_port, registers_23_14_port, 
      registers_23_13_port, registers_23_12_port, registers_23_11_port, 
      registers_23_10_port, registers_23_9_port, registers_23_8_port, 
      registers_23_7_port, registers_23_6_port, registers_23_5_port, 
      registers_23_4_port, registers_23_3_port, registers_23_2_port, 
      registers_23_1_port, registers_23_0_port, registers_24_31_port, 
      registers_24_30_port, registers_24_29_port, registers_24_28_port, 
      registers_24_27_port, registers_24_26_port, registers_24_25_port, 
      registers_24_24_port, registers_24_23_port, registers_24_22_port, 
      registers_24_21_port, registers_24_20_port, registers_24_19_port, 
      registers_24_18_port, registers_24_17_port, registers_24_16_port, 
      registers_24_15_port, registers_24_14_port, registers_24_13_port, 
      registers_24_12_port, registers_24_11_port, registers_24_10_port, 
      registers_24_9_port, registers_24_8_port, registers_24_7_port, 
      registers_24_6_port, registers_24_5_port, registers_24_4_port, 
      registers_24_3_port, registers_24_2_port, registers_24_1_port, 
      registers_24_0_port, registers_25_31_port, registers_25_30_port, 
      registers_25_29_port, registers_25_28_port, registers_25_27_port, 
      registers_25_26_port, registers_25_25_port, registers_25_24_port, 
      registers_25_23_port, registers_25_22_port, registers_25_21_port, 
      registers_25_20_port, registers_25_19_port, registers_25_18_port, 
      registers_25_17_port, registers_25_16_port, registers_25_15_port, 
      registers_25_14_port, registers_25_13_port, registers_25_12_port, 
      registers_25_11_port, registers_25_10_port, registers_25_9_port, 
      registers_25_8_port, registers_25_7_port, registers_25_6_port, 
      registers_25_5_port, registers_25_4_port, registers_25_3_port, 
      registers_25_2_port, registers_25_1_port, registers_25_0_port, 
      registers_26_31_port, registers_26_30_port, registers_26_29_port, 
      registers_26_28_port, registers_26_27_port, registers_26_26_port, 
      registers_26_25_port, registers_26_24_port, registers_26_23_port, 
      registers_26_22_port, registers_26_21_port, registers_26_20_port, 
      registers_26_19_port, registers_26_18_port, registers_26_17_port, 
      registers_26_16_port, registers_26_15_port, registers_26_14_port, 
      registers_26_13_port, registers_26_12_port, registers_26_11_port, 
      registers_26_10_port, registers_26_9_port, registers_26_8_port, 
      registers_26_7_port, registers_26_6_port, registers_26_5_port, 
      registers_26_4_port, registers_26_3_port, registers_26_2_port, 
      registers_26_1_port, registers_26_0_port, registers_27_31_port, 
      registers_27_30_port, registers_27_29_port, registers_27_28_port, 
      registers_27_27_port, registers_27_26_port, registers_27_25_port, 
      registers_27_24_port, registers_27_23_port, registers_27_22_port, 
      registers_27_21_port, registers_27_20_port, registers_27_19_port, 
      registers_27_18_port, registers_27_17_port, registers_27_16_port, 
      registers_27_15_port, registers_27_14_port, registers_27_13_port, 
      registers_27_12_port, registers_27_11_port, registers_27_10_port, 
      registers_27_9_port, registers_27_8_port, registers_27_7_port, 
      registers_27_6_port, registers_27_5_port, registers_27_4_port, 
      registers_27_3_port, registers_27_2_port, registers_27_1_port, 
      registers_27_0_port, registers_28_31_port, registers_28_30_port, 
      registers_28_29_port, registers_28_28_port, registers_28_27_port, 
      registers_28_26_port, registers_28_25_port, registers_28_24_port, 
      registers_28_23_port, registers_28_22_port, registers_28_21_port, 
      registers_28_20_port, registers_28_19_port, registers_28_18_port, 
      registers_28_17_port, registers_28_16_port, registers_28_15_port, 
      registers_28_14_port, registers_28_13_port, registers_28_12_port, 
      registers_28_11_port, registers_28_10_port, registers_28_9_port, 
      registers_28_8_port, registers_28_7_port, registers_28_6_port, 
      registers_28_5_port, registers_28_4_port, registers_28_3_port, 
      registers_28_2_port, registers_28_1_port, registers_28_0_port, 
      registers_29_31_port, registers_29_30_port, registers_29_29_port, 
      registers_29_28_port, registers_29_27_port, registers_29_26_port, 
      registers_29_25_port, registers_29_24_port, registers_29_23_port, 
      registers_29_22_port, registers_29_21_port, registers_29_20_port, 
      registers_29_19_port, registers_29_18_port, registers_29_17_port, 
      registers_29_16_port, registers_29_15_port, registers_29_14_port, 
      registers_29_13_port, registers_29_12_port, registers_29_11_port, 
      registers_29_10_port, registers_29_9_port, registers_29_8_port, 
      registers_29_7_port, registers_29_6_port, registers_29_5_port, 
      registers_29_4_port, registers_29_3_port, registers_29_2_port, 
      registers_29_1_port, registers_29_0_port, registers_30_31_port, 
      registers_30_30_port, registers_30_29_port, registers_30_28_port, 
      registers_30_27_port, registers_30_26_port, registers_30_25_port, 
      registers_30_24_port, registers_30_23_port, registers_30_22_port, 
      registers_30_21_port, registers_30_20_port, registers_30_19_port, 
      registers_30_18_port, registers_30_17_port, registers_30_16_port, 
      registers_30_15_port, registers_30_14_port, registers_30_13_port, 
      registers_30_12_port, registers_30_11_port, registers_30_10_port, 
      registers_30_9_port, registers_30_8_port, registers_30_7_port, 
      registers_30_6_port, registers_30_5_port, registers_30_4_port, 
      registers_30_3_port, registers_30_2_port, registers_30_1_port, 
      registers_30_0_port, registers_31_30_port, registers_31_29_port, 
      registers_31_28_port, registers_31_27_port, registers_31_26_port, 
      registers_31_25_port, registers_31_24_port, registers_31_23_port, 
      registers_31_22_port, registers_31_21_port, registers_31_20_port, 
      registers_31_19_port, registers_31_18_port, registers_31_17_port, 
      registers_31_16_port, registers_31_15_port, registers_31_14_port, 
      registers_31_13_port, registers_31_12_port, registers_31_11_port, 
      registers_31_10_port, registers_31_9_port, registers_31_8_port, 
      registers_31_7_port, registers_31_6_port, registers_31_5_port, 
      registers_31_4_port, registers_31_3_port, registers_31_2_port, 
      registers_31_1_port, registers_31_0_port, N18, n2919, n2920, n2921, n2922
      , n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, 
      n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, 
      n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2951, n2952, n2953, 
      n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, 
      n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, 
      n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, 
      n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, 
      n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, 
      n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, 
      n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, 
      n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, 
      n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, 
      n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, 
      n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, 
      n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, 
      n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, 
      n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, 
      n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, 
      n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, 
      n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, 
      n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, 
      n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, 
      n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, 
      n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, 
      n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, 
      n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, 
      n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, 
      n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, 
      n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, 
      n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, 
      n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, 
      n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, 
      n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, 
      n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, 
      n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, 
      n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, 
      n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, 
      n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, 
      n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, 
      n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, 
      n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, 
      n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, 
      n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, 
      n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, 
      n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, 
      n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, 
      n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, 
      n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, 
      n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, 
      n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, 
      n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, 
      n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, 
      n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, 
      n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, 
      n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, 
      n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, 
      n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, 
      n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, 
      n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, 
      n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, 
      n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, 
      n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, 
      n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, 
      n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, 
      n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, 
      n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, 
      n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, 
      n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, 
      n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, 
      n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, 
      n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, 
      n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, 
      n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, 
      n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, 
      n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, 
      n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, 
      n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, 
      n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, 
      n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, 
      n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, 
      n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, 
      n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, 
      n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, 
      n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, 
      n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, 
      n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, 
      n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, 
      n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, 
      n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, 
      n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, 
      n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, 
      n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, 
      n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, 
      n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, 
      n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, 
      n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, 
      n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, 
      n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, 
      n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, 
      n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, 
      n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, 
      n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, 
      n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, 
      n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, 
      n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, 
      n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, 
      n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, 
      n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, 
      n4004, n4005, n4006, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18_port, n19, n20, n21, n22, n23, n24, n25, n26
      , n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, 
      n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55
      , n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, 
      n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84
      , n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, 
      n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, 
      n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, 
      n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, 
      n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, 
      n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, 
      n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, 
      n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, 
      n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, 
      n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, 
      n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, 
      n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, 
      n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, 
      n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, 
      n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, 
      n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, 
      n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, 
      n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, 
      n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, 
      n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, 
      n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, 
      n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, 
      n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, 
      n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, 
      n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, 
      n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, 
      n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, 
      n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, 
      n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, 
      n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, 
      n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, 
      n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, 
      n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, 
      n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, 
      n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, 
      n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, 
      n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, 
      n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, 
      n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, 
      n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, 
      n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, 
      n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, 
      n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, 
      n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, 
      n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, 
      n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, 
      n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, 
      n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, 
      n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, 
      n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, 
      n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, 
      n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, 
      n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, 
      n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, 
      n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, 
      n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, 
      n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, 
      n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, 
      n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, 
      n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, 
      n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, 
      n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, 
      n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, 
      n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, 
      n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, 
      n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, 
      n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, 
      n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, 
      n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, 
      n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, 
      n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, 
      n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, 
      n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, 
      n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, 
      n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, 
      n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, 
      n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, 
      n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, 
      n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, 
      n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, 
      n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, 
      n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, 
      n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, 
      n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, 
      n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, 
      n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, 
      n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, 
      n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, 
      n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, 
      n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, 
      n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, 
      n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, 
      n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, 
      n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, 
      n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, 
      n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, 
      n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, 
      n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, 
      n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, 
      n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, 
      n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, 
      n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, 
      n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, 
      n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, 
      n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, 
      n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, 
      n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, 
      n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, 
      n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, 
      n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, 
      n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, 
      n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, 
      n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, 
      n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, 
      n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, 
      n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, 
      n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, 
      n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, 
      n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, 
      n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, 
      n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, 
      n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, 
      n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, 
      n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, 
      n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, 
      n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, 
      n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, 
      n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, 
      n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, 
      n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, 
      n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, 
      n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, 
      n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, 
      n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, 
      n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, 
      n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, 
      n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, 
      n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, 
      n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, 
      n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, 
      n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, 
      n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, 
      n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, 
      n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, 
      n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, 
      n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, 
      n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, 
      n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, 
      n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, 
      n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, 
      n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, 
      n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, 
      n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, 
      n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, 
      n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, 
      n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, 
      n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, 
      n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, 
      n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, 
      n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, 
      n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, 
      n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, 
      n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, 
      n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, 
      n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, 
      n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, 
      n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, 
      n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, 
      n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, 
      n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, 
      n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, 
      n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, 
      n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, 
      n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, 
      n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, 
      n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, 
      n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, 
      n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, 
      n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, 
      n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, 
      n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, 
      n2049, net108129, net108130, net108131, net108132, net108133, net108134, 
      net108135, net108136, net108137, net108138, net108139, net108140, 
      net108141, net108142, net108143, net108144, net108145, net108146, 
      net108147, net108148, net108149, net108150, net108151, net108152, 
      net108153, net108154, net108155, net108156, net108157, net108158, 
      net108159, net108160, net108161, net108162, net108163, net108164, 
      net108165, net108166, net108167, net108168, net108169, net108170, 
      net108171, net108172, net108173, net108174, net108175, net108176, 
      net108177, net108178, net108179, net108180, net108181, net108182, 
      net108183, net108184, net108185, net108186, net108187, net108188, 
      net108189, net108190, net108191, net108192, net108193, net108194, 
      net108195, net108196, net108197, net108198, net108199, net108200, 
      net108201, net108202, net108203, net108204, net108205, net108206, 
      net108207, net108208, net108209, net108210, net108211, net108212, 
      net108213, net108214, net108215, net108216, net108217, net108218, 
      net108219, net108220, net108221, net108222, net108223, net108224, 
      net108225, net108226, net108227, net108228, net108229, net108230, 
      net108231, net108232, net108233, net108234, net108235, net108236, 
      net108237, net108238, net108239, net108240, net108241, net108242, 
      net108243, net108244, net108245, net108246, net108247, net108248, 
      net108249, net108250, net108251, net108252, net108253, net108254, 
      net108255, net108256, net108257, net108258, net108259, net108260, 
      net108261, net108262, net108263, net108264, net108265, net108266, 
      net108267, net108268, net108269, net108270, net108271, net108272, 
      net108273, net108274, net108275, net108276, net108277, net108278, 
      net108279, net108280, net108281, net108282, net108283, net108284, 
      net108285, net108286, net108287, net108288, net108289, net108290, 
      net108291, net108292, net108293, net108294, net108295, net108296, 
      net108297, net108298, net108299, net108300, net108301, net108302, 
      net108303, net108304, net108305, net108306, net108307, net108308, 
      net108309, net108310, net108311, net108312, net108313, net108314, 
      net108315, net108316, net108317, net108318, net108319, net108320, 
      net108321, net108322, net108323, net108324, net108325, net108326, 
      net108327, net108328, net108329, net108330, net108331, net108332, 
      net108333, net108334, net108335, net108336, net108337, net108338, 
      net108339, net108340, net108341, net108342, net108343, net108344, 
      net108345, net108346, net108347, net108348, net108349, net108350, 
      net108351, net108352, net108353, net108354, net108355, net108356, 
      net108357, net108358, net108359, net108360, net108361, net108362, 
      net108363, net108364, net108365, net108366, net108367, net108368, 
      net108369, net108370, net108371, net108372, net108373, net108374, 
      net108375, net108376, net108377, net108378, net108379, net108380, 
      net108381, net108382, net108383, net108384, net108385, net108386, 
      net108387, net108388, net108389, net108390, net108391, net108392, 
      net108393, net108394, net108395, net108396, net108397, net108398, 
      net108399, net108400, net108401, net108402, net108403, net108404, 
      net108405, net108406, net108407, net108408, net108409, net108410, 
      net108411, net108412, net108413, net108414, net108415, net108416, 
      net108417, net108418, net108419, net108420, net108421, net108422, 
      net108423, net108424, net108425, net108426, net108427, net108428, 
      net108429, net108430, net108431, net108432, net108433, net108434, 
      net108435, net108436, net108437, net108438, net108439, net108440, 
      net108441, net108442, net108443, net108444, net108445, net108446, 
      net108447, net108448, net108449, net108450, net108451, net108452, 
      net108453, net108454, net108455, net108456, net108457, net108458, 
      net108459, net108460, net108461, net108462, net108463, net108464, 
      net108465, net108466, net108467, net108468, net108469, net108470, 
      net108471, net108472, net108473, net108474, net108475, net108476, 
      net108477, net108478, net108479, net108480, net108481, net108482, 
      net108483, net108484, net108485, net108486, net108487, net108488, 
      net108489, net108490, net108491, net108492, net108493, net108494, 
      net108495, net108496, net108497, net108498, net108499, net108500, 
      net108501, net108502, net108503, net108504, net108505, net108506, 
      net108507, net108508, net108509, net108510, net108511, net108512, 
      net108513, net108514, net108515, net108516, net108517, net108518, 
      net108519, net108520, net108521, net108522, net108523, net108524, 
      net108525, net108526, net108527, net108528, net108529, net108530, 
      net108531, net108532, net108533, net108534, net108535, net108536, 
      net108537, net108538, net108539, net108540, net108541, net108542, 
      net108543, net108544, net108545, net108546, net108547, net108548, 
      net108549, net108550, net108551, net108552, net108553, net108554, 
      net108555, net108556, net108557, net108558, net108559, net108560, 
      net108561, net108562, net108563, net108564, net108565, net108566, 
      net108567, net108568, net108569, net108570, net108571, net108572, 
      net108573, net108574, net108575, net108576, net108577, net108578, 
      net108579, net108580, net108581, net108582, net108583, net108584, 
      net108585, net108586, net108587, net108588, net108589, net108590, 
      net108591, net108592, net108593, net108594, net108595, net108596, 
      net108597, net108598, net108599, net108600, net108601, net108602, 
      net108603, net108604, net108605, net108606, net108607, net108608, 
      net108609, net108610 : std_logic;

begin
   d_out1 <= ( d_out1_31_port, d_out1_30_port, d_out1_29_port, d_out1_28_port, 
      d_out1_27_port, d_out1_26_port, d_out1_25_port, d_out1_24_port, 
      d_out1_23_port, d_out1_22_port, d_out1_21_port, d_out1_20_port, 
      d_out1_19_port, d_out1_18_port, d_out1_17_port, d_out1_16_port, 
      d_out1_15_port, d_out1_14_port, d_out1_13_port, d_out1_12_port, 
      d_out1_11_port, d_out1_10_port, d_out1_9_port, d_out1_8_port, 
      d_out1_7_port, d_out1_6_port, d_out1_5_port, d_out1_4_port, d_out1_3_port
      , d_out1_2_port, d_out1_1_port, d_out1_0_port );
   d_out2 <= ( d_out2_31_port, d_out2_30_port, d_out2_29_port, d_out2_28_port, 
      d_out2_27_port, d_out2_26_port, d_out2_25_port, d_out2_24_port, 
      d_out2_23_port, d_out2_22_port, d_out2_21_port, d_out2_20_port, 
      d_out2_19_port, d_out2_18_port, d_out2_17_port, d_out2_16_port, 
      d_out2_15_port, d_out2_14_port, d_out2_13_port, d_out2_12_port, 
      d_out2_11_port, d_out2_10_port, d_out2_9_port, d_out2_8_port, 
      d_out2_7_port, d_out2_6_port, d_out2_5_port, d_out2_4_port, d_out2_3_port
      , d_out2_2_port, d_out2_1_port, d_out2_0_port );
   
   registers_reg_1_31_inst : DFFR_X1 port map( D => n4006, CK => n569, RN => 
                           rst, Q => registers_1_31_port, QN => n541);
   registers_reg_1_30_inst : DFFR_X1 port map( D => n4005, CK => n572, RN => 
                           rst, Q => registers_1_30_port, QN => n353);
   registers_reg_1_29_inst : DFFR_X1 port map( D => n4004, CK => n574, RN => 
                           rst, Q => registers_1_29_port, QN => n355);
   registers_reg_1_28_inst : DFFR_X1 port map( D => n4003, CK => n577, RN => 
                           rst, Q => registers_1_28_port, QN => n357);
   registers_reg_1_27_inst : DFFR_X1 port map( D => n4002, CK => n584, RN => 
                           rst, Q => registers_1_27_port, QN => n359);
   registers_reg_1_26_inst : DFFR_X1 port map( D => n4001, CK => n550, RN => 
                           rst, Q => registers_1_26_port, QN => n361);
   registers_reg_1_25_inst : DFFR_X1 port map( D => n4000, CK => n565, RN => 
                           rst, Q => registers_1_25_port, QN => n363);
   registers_reg_1_24_inst : DFFR_X1 port map( D => n3999, CK => n587, RN => 
                           rst, Q => registers_1_24_port, QN => n365);
   registers_reg_1_23_inst : DFFR_X1 port map( D => n3998, CK => n552, RN => 
                           rst, Q => registers_1_23_port, QN => n367);
   registers_reg_1_22_inst : DFFR_X1 port map( D => n3997, CK => n568, RN => 
                           rst, Q => registers_1_22_port, QN => n369);
   registers_reg_1_21_inst : DFFR_X1 port map( D => n3996, CK => n623, RN => 
                           rst, Q => registers_1_21_port, QN => n371);
   registers_reg_1_20_inst : DFFR_X1 port map( D => n3995, CK => n555, RN => 
                           rst, Q => registers_1_20_port, QN => n373);
   registers_reg_1_19_inst : DFFR_X1 port map( D => n3994, CK => n617, RN => 
                           rst, Q => registers_1_19_port, QN => n375);
   registers_reg_1_18_inst : DFFR_X1 port map( D => n3993, CK => n557, RN => 
                           rst, Q => registers_1_18_port, QN => n377);
   registers_reg_1_17_inst : DFFR_X1 port map( D => n3992, CK => n630, RN => 
                           rst, Q => registers_1_17_port, QN => n379);
   registers_reg_1_16_inst : DFFR_X1 port map( D => n3991, CK => n634, RN => 
                           rst, Q => registers_1_16_port, QN => n381);
   registers_reg_1_15_inst : DFFR_X1 port map( D => n3990, CK => n559, RN => 
                           rst, Q => registers_1_15_port, QN => n383);
   registers_reg_1_14_inst : DFFR_X1 port map( D => n3989, CK => n599, RN => 
                           rst, Q => registers_1_14_port, QN => n385);
   registers_reg_1_13_inst : DFFR_X1 port map( D => n3988, CK => n602, RN => 
                           rst, Q => registers_1_13_port, QN => n387);
   registers_reg_1_12_inst : DFFR_X1 port map( D => n3987, CK => n627, RN => 
                           rst, Q => registers_1_12_port, QN => n389);
   registers_reg_1_11_inst : DFFR_X1 port map( D => n3986, CK => n594, RN => 
                           rst, Q => registers_1_11_port, QN => n391);
   registers_reg_1_10_inst : DFFR_X1 port map( D => n3985, CK => n611, RN => 
                           rst, Q => registers_1_10_port, QN => n393);
   registers_reg_1_9_inst : DFFR_X1 port map( D => n3984, CK => n590, RN => rst
                           , Q => registers_1_9_port, QN => n395);
   registers_reg_1_8_inst : DFFR_X1 port map( D => n3983, CK => n562, RN => rst
                           , Q => registers_1_8_port, QN => n397);
   registers_reg_1_7_inst : DFFR_X1 port map( D => n3982, CK => n547, RN => rst
                           , Q => registers_1_7_port, QN => n399);
   registers_reg_1_6_inst : DFFR_X1 port map( D => n3981, CK => n597, RN => rst
                           , Q => registers_1_6_port, QN => n401);
   registers_reg_1_5_inst : DFFR_X1 port map( D => n3980, CK => n581, RN => rst
                           , Q => registers_1_5_port, QN => n403);
   registers_reg_1_4_inst : DFFR_X1 port map( D => n3979, CK => n620, RN => rst
                           , Q => registers_1_4_port, QN => n405);
   registers_reg_1_3_inst : DFFR_X1 port map( D => n3978, CK => n613, RN => rst
                           , Q => registers_1_3_port, QN => n407);
   registers_reg_1_2_inst : DFFR_X1 port map( D => n3977, CK => n608, RN => rst
                           , Q => registers_1_2_port, QN => n409);
   registers_reg_1_1_inst : DFFR_X1 port map( D => n3976, CK => n615, RN => rst
                           , Q => registers_1_1_port, QN => n411);
   registers_reg_1_0_inst : DFFR_X1 port map( D => n3975, CK => n592, RN => rst
                           , Q => registers_1_0_port, QN => n413);
   registers_reg_2_31_inst : DFFR_X1 port map( D => n3974, CK => n569, RN => 
                           rst, Q => registers_2_31_port, QN => n543);
   registers_reg_2_30_inst : DFFR_X1 port map( D => n3973, CK => n571, RN => 
                           rst, Q => registers_2_30_port, QN => n480);
   registers_reg_2_29_inst : DFFR_X1 port map( D => n3972, CK => n574, RN => 
                           rst, Q => registers_2_29_port, QN => n482);
   registers_reg_2_28_inst : DFFR_X1 port map( D => n3971, CK => n577, RN => 
                           rst, Q => registers_2_28_port, QN => n484);
   registers_reg_2_27_inst : DFFR_X1 port map( D => n3970, CK => n584, RN => 
                           rst, Q => registers_2_27_port, QN => n486);
   registers_reg_2_26_inst : DFFR_X1 port map( D => n3969, CK => n550, RN => 
                           rst, Q => registers_2_26_port, QN => n488);
   registers_reg_2_25_inst : DFFR_X1 port map( D => n3968, CK => n565, RN => 
                           rst, Q => registers_2_25_port, QN => n490);
   registers_reg_2_24_inst : DFFR_X1 port map( D => n3967, CK => n587, RN => 
                           rst, Q => registers_2_24_port, QN => n492);
   registers_reg_2_23_inst : DFFR_X1 port map( D => n3966, CK => n552, RN => 
                           rst, Q => registers_2_23_port, QN => n494);
   registers_reg_2_22_inst : DFFR_X1 port map( D => n3965, CK => n568, RN => 
                           rst, Q => registers_2_22_port, QN => n496);
   registers_reg_2_21_inst : DFFR_X1 port map( D => n3964, CK => n623, RN => 
                           rst, Q => registers_2_21_port, QN => n498);
   registers_reg_2_20_inst : DFFR_X1 port map( D => n3963, CK => n555, RN => 
                           rst, Q => registers_2_20_port, QN => n500);
   registers_reg_2_19_inst : DFFR_X1 port map( D => n3962, CK => n617, RN => 
                           rst, Q => registers_2_19_port, QN => n502);
   registers_reg_2_18_inst : DFFR_X1 port map( D => n3961, CK => n557, RN => 
                           rst, Q => registers_2_18_port, QN => n504);
   registers_reg_2_17_inst : DFFR_X1 port map( D => n3960, CK => n630, RN => 
                           rst, Q => registers_2_17_port, QN => n506);
   registers_reg_2_16_inst : DFFR_X1 port map( D => n3959, CK => n634, RN => 
                           rst, Q => registers_2_16_port, QN => n508);
   registers_reg_2_15_inst : DFFR_X1 port map( D => n3958, CK => n559, RN => 
                           rst, Q => registers_2_15_port, QN => n510);
   registers_reg_2_14_inst : DFFR_X1 port map( D => n3957, CK => n599, RN => 
                           rst, Q => registers_2_14_port, QN => n512);
   registers_reg_2_13_inst : DFFR_X1 port map( D => n3956, CK => n602, RN => 
                           rst, Q => registers_2_13_port, QN => n514);
   registers_reg_2_12_inst : DFFR_X1 port map( D => n3955, CK => n627, RN => 
                           rst, Q => registers_2_12_port, QN => n516);
   registers_reg_2_11_inst : DFFR_X1 port map( D => n3954, CK => n594, RN => 
                           rst, Q => registers_2_11_port, QN => n518);
   registers_reg_2_10_inst : DFFR_X1 port map( D => n3953, CK => n611, RN => 
                           rst, Q => registers_2_10_port, QN => n520);
   registers_reg_2_9_inst : DFFR_X1 port map( D => n3952, CK => n590, RN => rst
                           , Q => registers_2_9_port, QN => n522);
   registers_reg_2_8_inst : DFFR_X1 port map( D => n3951, CK => n562, RN => rst
                           , Q => registers_2_8_port, QN => n524);
   registers_reg_2_7_inst : DFFR_X1 port map( D => n3950, CK => n547, RN => rst
                           , Q => registers_2_7_port, QN => n526);
   registers_reg_2_6_inst : DFFR_X1 port map( D => n3949, CK => n597, RN => rst
                           , Q => registers_2_6_port, QN => n528);
   registers_reg_2_5_inst : DFFR_X1 port map( D => n3948, CK => n581, RN => rst
                           , Q => registers_2_5_port, QN => n530);
   registers_reg_2_4_inst : DFFR_X1 port map( D => n3947, CK => n620, RN => rst
                           , Q => registers_2_4_port, QN => n532);
   registers_reg_2_3_inst : DFFR_X1 port map( D => n3946, CK => n613, RN => rst
                           , Q => registers_2_3_port, QN => n534);
   registers_reg_2_2_inst : DFFR_X1 port map( D => n3945, CK => n608, RN => rst
                           , Q => registers_2_2_port, QN => n536);
   registers_reg_2_1_inst : DFFR_X1 port map( D => n3944, CK => n615, RN => rst
                           , Q => registers_2_1_port, QN => n538);
   registers_reg_2_0_inst : DFFR_X1 port map( D => n3943, CK => n545, RN => rst
                           , Q => registers_2_0_port, QN => n540);
   registers_reg_3_31_inst : DFFR_X1 port map( D => n3942, CK => n569, RN => 
                           rst, Q => registers_3_31_port, QN => net108610);
   registers_reg_3_30_inst : DFFR_X1 port map( D => n3941, CK => n571, RN => 
                           rst, Q => registers_3_30_port, QN => net108609);
   registers_reg_3_29_inst : DFFR_X1 port map( D => n3940, CK => n574, RN => 
                           rst, Q => registers_3_29_port, QN => net108608);
   registers_reg_3_28_inst : DFFR_X1 port map( D => n3939, CK => n577, RN => 
                           rst, Q => registers_3_28_port, QN => net108607);
   registers_reg_3_27_inst : DFFR_X1 port map( D => n3938, CK => n584, RN => 
                           rst, Q => registers_3_27_port, QN => net108606);
   registers_reg_3_26_inst : DFFR_X1 port map( D => n3937, CK => n549, RN => 
                           rst, Q => registers_3_26_port, QN => net108605);
   registers_reg_3_25_inst : DFFR_X1 port map( D => n3936, CK => n565, RN => 
                           rst, Q => registers_3_25_port, QN => net108604);
   registers_reg_3_24_inst : DFFR_X1 port map( D => n3935, CK => n587, RN => 
                           rst, Q => registers_3_24_port, QN => net108603);
   registers_reg_3_23_inst : DFFR_X1 port map( D => n3934, CK => n552, RN => 
                           rst, Q => registers_3_23_port, QN => net108602);
   registers_reg_3_22_inst : DFFR_X1 port map( D => n3933, CK => n568, RN => 
                           rst, Q => registers_3_22_port, QN => net108601);
   registers_reg_3_21_inst : DFFR_X1 port map( D => n3932, CK => n623, RN => 
                           rst, Q => registers_3_21_port, QN => net108600);
   registers_reg_3_20_inst : DFFR_X1 port map( D => n3931, CK => n555, RN => 
                           rst, Q => registers_3_20_port, QN => net108599);
   registers_reg_3_19_inst : DFFR_X1 port map( D => n3930, CK => n617, RN => 
                           rst, Q => registers_3_19_port, QN => net108598);
   registers_reg_3_18_inst : DFFR_X1 port map( D => n3929, CK => n557, RN => 
                           rst, Q => registers_3_18_port, QN => net108597);
   registers_reg_3_17_inst : DFFR_X1 port map( D => n3928, CK => n630, RN => 
                           rst, Q => registers_3_17_port, QN => net108596);
   registers_reg_3_16_inst : DFFR_X1 port map( D => n3927, CK => n632, RN => 
                           rst, Q => registers_3_16_port, QN => net108595);
   registers_reg_3_15_inst : DFFR_X1 port map( D => n3926, CK => n559, RN => 
                           rst, Q => registers_3_15_port, QN => net108594);
   registers_reg_3_14_inst : DFFR_X1 port map( D => n3925, CK => n599, RN => 
                           rst, Q => registers_3_14_port, QN => net108593);
   registers_reg_3_13_inst : DFFR_X1 port map( D => n3924, CK => n602, RN => 
                           rst, Q => registers_3_13_port, QN => net108592);
   registers_reg_3_12_inst : DFFR_X1 port map( D => n3923, CK => n627, RN => 
                           rst, Q => registers_3_12_port, QN => net108591);
   registers_reg_3_11_inst : DFFR_X1 port map( D => n3922, CK => n594, RN => 
                           rst, Q => registers_3_11_port, QN => net108590);
   registers_reg_3_10_inst : DFFR_X1 port map( D => n3921, CK => n611, RN => 
                           rst, Q => registers_3_10_port, QN => net108589);
   registers_reg_3_9_inst : DFFR_X1 port map( D => n3920, CK => n589, RN => rst
                           , Q => registers_3_9_port, QN => net108588);
   registers_reg_3_8_inst : DFFR_X1 port map( D => n3919, CK => n562, RN => rst
                           , Q => registers_3_8_port, QN => net108587);
   registers_reg_3_7_inst : DFFR_X1 port map( D => n3918, CK => n547, RN => rst
                           , Q => registers_3_7_port, QN => net108586);
   registers_reg_3_6_inst : DFFR_X1 port map( D => n3917, CK => n596, RN => rst
                           , Q => registers_3_6_port, QN => net108585);
   registers_reg_3_5_inst : DFFR_X1 port map( D => n3916, CK => n581, RN => rst
                           , Q => registers_3_5_port, QN => net108584);
   registers_reg_3_4_inst : DFFR_X1 port map( D => n3915, CK => n620, RN => rst
                           , Q => registers_3_4_port, QN => net108583);
   registers_reg_3_3_inst : DFFR_X1 port map( D => n3914, CK => n613, RN => rst
                           , Q => registers_3_3_port, QN => net108582);
   registers_reg_3_2_inst : DFFR_X1 port map( D => n3913, CK => n608, RN => rst
                           , Q => registers_3_2_port, QN => net108581);
   registers_reg_3_1_inst : DFFR_X1 port map( D => n3912, CK => n614, RN => rst
                           , Q => registers_3_1_port, QN => net108580);
   registers_reg_3_0_inst : DFFR_X1 port map( D => n3911, CK => n580, RN => rst
                           , Q => registers_3_0_port, QN => net108579);
   registers_reg_4_31_inst : DFFR_X1 port map( D => n3910, CK => n569, RN => 
                           rst, Q => registers_4_31_port, QN => net108578);
   registers_reg_4_30_inst : DFFR_X1 port map( D => n3909, CK => n571, RN => 
                           rst, Q => registers_4_30_port, QN => net108577);
   registers_reg_4_29_inst : DFFR_X1 port map( D => n3908, CK => n574, RN => 
                           rst, Q => registers_4_29_port, QN => net108576);
   registers_reg_4_28_inst : DFFR_X1 port map( D => n3907, CK => n577, RN => 
                           rst, Q => registers_4_28_port, QN => net108575);
   registers_reg_4_27_inst : DFFR_X1 port map( D => n3906, CK => n584, RN => 
                           rst, Q => registers_4_27_port, QN => net108574);
   registers_reg_4_26_inst : DFFR_X1 port map( D => n3905, CK => n549, RN => 
                           rst, Q => registers_4_26_port, QN => net108573);
   registers_reg_4_25_inst : DFFR_X1 port map( D => n3904, CK => n565, RN => 
                           rst, Q => registers_4_25_port, QN => net108572);
   registers_reg_4_24_inst : DFFR_X1 port map( D => n3903, CK => n587, RN => 
                           rst, Q => registers_4_24_port, QN => net108571);
   registers_reg_4_23_inst : DFFR_X1 port map( D => n3902, CK => n552, RN => 
                           rst, Q => registers_4_23_port, QN => net108570);
   registers_reg_4_22_inst : DFFR_X1 port map( D => n3901, CK => n567, RN => 
                           rst, Q => registers_4_22_port, QN => net108569);
   registers_reg_4_21_inst : DFFR_X1 port map( D => n3900, CK => n623, RN => 
                           rst, Q => registers_4_21_port, QN => net108568);
   registers_reg_4_20_inst : DFFR_X1 port map( D => n3899, CK => n555, RN => 
                           rst, Q => registers_4_20_port, QN => net108567);
   registers_reg_4_19_inst : DFFR_X1 port map( D => n3898, CK => n617, RN => 
                           rst, Q => registers_4_19_port, QN => net108566);
   registers_reg_4_18_inst : DFFR_X1 port map( D => n3897, CK => n556, RN => 
                           rst, Q => registers_4_18_port, QN => net108565);
   registers_reg_4_17_inst : DFFR_X1 port map( D => n3896, CK => n630, RN => 
                           rst, Q => registers_4_17_port, QN => net108564);
   registers_reg_4_16_inst : DFFR_X1 port map( D => n3895, CK => n633, RN => 
                           rst, Q => registers_4_16_port, QN => net108563);
   registers_reg_4_15_inst : DFFR_X1 port map( D => n3894, CK => n559, RN => 
                           rst, Q => registers_4_15_port, QN => net108562);
   registers_reg_4_14_inst : DFFR_X1 port map( D => n3893, CK => n599, RN => 
                           rst, Q => registers_4_14_port, QN => net108561);
   registers_reg_4_13_inst : DFFR_X1 port map( D => n3892, CK => n602, RN => 
                           rst, Q => registers_4_13_port, QN => net108560);
   registers_reg_4_12_inst : DFFR_X1 port map( D => n3891, CK => n627, RN => 
                           rst, Q => registers_4_12_port, QN => net108559);
   registers_reg_4_11_inst : DFFR_X1 port map( D => n3890, CK => n594, RN => 
                           rst, Q => registers_4_11_port, QN => net108558);
   registers_reg_4_10_inst : DFFR_X1 port map( D => n3889, CK => n611, RN => 
                           rst, Q => registers_4_10_port, QN => net108557);
   registers_reg_4_9_inst : DFFR_X1 port map( D => n3888, CK => n589, RN => rst
                           , Q => registers_4_9_port, QN => net108556);
   registers_reg_4_8_inst : DFFR_X1 port map( D => n3887, CK => n562, RN => rst
                           , Q => registers_4_8_port, QN => net108555);
   registers_reg_4_7_inst : DFFR_X1 port map( D => n3886, CK => n547, RN => rst
                           , Q => registers_4_7_port, QN => net108554);
   registers_reg_4_6_inst : DFFR_X1 port map( D => n3885, CK => n596, RN => rst
                           , Q => registers_4_6_port, QN => net108553);
   registers_reg_4_5_inst : DFFR_X1 port map( D => n3884, CK => n581, RN => rst
                           , Q => registers_4_5_port, QN => net108552);
   registers_reg_4_4_inst : DFFR_X1 port map( D => n3883, CK => n620, RN => rst
                           , Q => registers_4_4_port, QN => net108551);
   registers_reg_4_3_inst : DFFR_X1 port map( D => n3882, CK => n613, RN => rst
                           , Q => registers_4_3_port, QN => net108550);
   registers_reg_4_2_inst : DFFR_X1 port map( D => n3881, CK => n608, RN => rst
                           , Q => registers_4_2_port, QN => net108549);
   registers_reg_4_1_inst : DFFR_X1 port map( D => n3880, CK => n614, RN => rst
                           , Q => registers_4_1_port, QN => net108548);
   registers_reg_4_0_inst : DFFR_X1 port map( D => n3879, CK => n580, RN => rst
                           , Q => registers_4_0_port, QN => net108547);
   registers_reg_5_31_inst : DFFR_X1 port map( D => n3878, CK => n568, RN => 
                           rst, Q => registers_5_31_port, QN => n290);
   registers_reg_5_30_inst : DFFR_X1 port map( D => n3877, CK => n571, RN => 
                           rst, Q => registers_5_30_port, QN => n291);
   registers_reg_5_29_inst : DFFR_X1 port map( D => n3876, CK => n574, RN => 
                           rst, Q => registers_5_29_port, QN => n292);
   registers_reg_5_28_inst : DFFR_X1 port map( D => n3875, CK => n577, RN => 
                           rst, Q => registers_5_28_port, QN => n293);
   registers_reg_5_27_inst : DFFR_X1 port map( D => n3874, CK => n584, RN => 
                           rst, Q => registers_5_27_port, QN => n294);
   registers_reg_5_26_inst : DFFR_X1 port map( D => n3873, CK => n549, RN => 
                           rst, Q => registers_5_26_port, QN => n295);
   registers_reg_5_25_inst : DFFR_X1 port map( D => n3872, CK => n565, RN => 
                           rst, Q => registers_5_25_port, QN => n296);
   registers_reg_5_24_inst : DFFR_X1 port map( D => n3871, CK => n587, RN => 
                           rst, Q => registers_5_24_port, QN => n297);
   registers_reg_5_23_inst : DFFR_X1 port map( D => n3870, CK => n552, RN => 
                           rst, Q => registers_5_23_port, QN => n298);
   registers_reg_5_22_inst : DFFR_X1 port map( D => n3869, CK => n567, RN => 
                           rst, Q => registers_5_22_port, QN => n299);
   registers_reg_5_21_inst : DFFR_X1 port map( D => n3868, CK => n623, RN => 
                           rst, Q => registers_5_21_port, QN => n300);
   registers_reg_5_20_inst : DFFR_X1 port map( D => n3867, CK => n555, RN => 
                           rst, Q => registers_5_20_port, QN => n301);
   registers_reg_5_19_inst : DFFR_X1 port map( D => n3866, CK => n617, RN => 
                           rst, Q => registers_5_19_port, QN => n302);
   registers_reg_5_18_inst : DFFR_X1 port map( D => n3865, CK => n556, RN => 
                           rst, Q => registers_5_18_port, QN => n303);
   registers_reg_5_17_inst : DFFR_X1 port map( D => n3864, CK => n629, RN => 
                           rst, Q => registers_5_17_port, QN => n304);
   registers_reg_5_16_inst : DFFR_X1 port map( D => n3863, CK => n633, RN => 
                           rst, Q => registers_5_16_port, QN => n305);
   registers_reg_5_15_inst : DFFR_X1 port map( D => n3862, CK => n559, RN => 
                           rst, Q => registers_5_15_port, QN => n306);
   registers_reg_5_14_inst : DFFR_X1 port map( D => n3861, CK => n599, RN => 
                           rst, Q => registers_5_14_port, QN => n307);
   registers_reg_5_13_inst : DFFR_X1 port map( D => n3860, CK => n602, RN => 
                           rst, Q => registers_5_13_port, QN => n308);
   registers_reg_5_12_inst : DFFR_X1 port map( D => n3859, CK => n627, RN => 
                           rst, Q => registers_5_12_port, QN => n309);
   registers_reg_5_11_inst : DFFR_X1 port map( D => n3858, CK => n594, RN => 
                           rst, Q => registers_5_11_port, QN => n310);
   registers_reg_5_10_inst : DFFR_X1 port map( D => n3857, CK => n610, RN => 
                           rst, Q => registers_5_10_port, QN => n311);
   registers_reg_5_9_inst : DFFR_X1 port map( D => n3856, CK => n589, RN => rst
                           , Q => registers_5_9_port, QN => n312);
   registers_reg_5_8_inst : DFFR_X1 port map( D => n3855, CK => n562, RN => rst
                           , Q => registers_5_8_port, QN => n313);
   registers_reg_5_7_inst : DFFR_X1 port map( D => n3854, CK => n547, RN => rst
                           , Q => registers_5_7_port, QN => n314);
   registers_reg_5_6_inst : DFFR_X1 port map( D => n3853, CK => n596, RN => rst
                           , Q => registers_5_6_port, QN => n315);
   registers_reg_5_5_inst : DFFR_X1 port map( D => n3852, CK => n581, RN => rst
                           , Q => registers_5_5_port, QN => n316);
   registers_reg_5_4_inst : DFFR_X1 port map( D => n3851, CK => n620, RN => rst
                           , Q => registers_5_4_port, QN => n317);
   registers_reg_5_3_inst : DFFR_X1 port map( D => n3850, CK => n613, RN => rst
                           , Q => registers_5_3_port, QN => n318);
   registers_reg_5_2_inst : DFFR_X1 port map( D => n3849, CK => n608, RN => rst
                           , Q => registers_5_2_port, QN => n319);
   registers_reg_5_1_inst : DFFR_X1 port map( D => n3848, CK => n614, RN => rst
                           , Q => registers_5_1_port, QN => n320);
   registers_reg_5_0_inst : DFFR_X1 port map( D => n3847, CK => n580, RN => rst
                           , Q => registers_5_0_port, QN => n321);
   registers_reg_6_31_inst : DFFR_X1 port map( D => n3846, CK => n568, RN => 
                           rst, Q => registers_6_31_port, QN => net108546);
   registers_reg_6_30_inst : DFFR_X1 port map( D => n3845, CK => n571, RN => 
                           rst, Q => registers_6_30_port, QN => net108545);
   registers_reg_6_29_inst : DFFR_X1 port map( D => n3844, CK => n574, RN => 
                           rst, Q => registers_6_29_port, QN => net108544);
   registers_reg_6_28_inst : DFFR_X1 port map( D => n3843, CK => n577, RN => 
                           rst, Q => registers_6_28_port, QN => net108543);
   registers_reg_6_27_inst : DFFR_X1 port map( D => n3842, CK => n584, RN => 
                           rst, Q => registers_6_27_port, QN => net108542);
   registers_reg_6_26_inst : DFFR_X1 port map( D => n3841, CK => n549, RN => 
                           rst, Q => registers_6_26_port, QN => net108541);
   registers_reg_6_25_inst : DFFR_X1 port map( D => n3840, CK => n565, RN => 
                           rst, Q => registers_6_25_port, QN => net108540);
   registers_reg_6_24_inst : DFFR_X1 port map( D => n3839, CK => n586, RN => 
                           rst, Q => registers_6_24_port, QN => net108539);
   registers_reg_6_23_inst : DFFR_X1 port map( D => n3838, CK => n552, RN => 
                           rst, Q => registers_6_23_port, QN => net108538);
   registers_reg_6_22_inst : DFFR_X1 port map( D => n3837, CK => n567, RN => 
                           rst, Q => registers_6_22_port, QN => net108537);
   registers_reg_6_21_inst : DFFR_X1 port map( D => n3836, CK => n622, RN => 
                           rst, Q => registers_6_21_port, QN => net108536);
   registers_reg_6_20_inst : DFFR_X1 port map( D => n3835, CK => n555, RN => 
                           rst, Q => registers_6_20_port, QN => net108535);
   registers_reg_6_19_inst : DFFR_X1 port map( D => n3834, CK => n617, RN => 
                           rst, Q => registers_6_19_port, QN => net108534);
   registers_reg_6_18_inst : DFFR_X1 port map( D => n3833, CK => n562, RN => 
                           rst, Q => registers_6_18_port, QN => net108533);
   registers_reg_6_17_inst : DFFR_X1 port map( D => n3832, CK => n629, RN => 
                           rst, Q => registers_6_17_port, QN => net108532);
   registers_reg_6_16_inst : DFFR_X1 port map( D => n3831, CK => n633, RN => 
                           rst, Q => registers_6_16_port, QN => net108531);
   registers_reg_6_15_inst : DFFR_X1 port map( D => n3830, CK => n559, RN => 
                           rst, Q => registers_6_15_port, QN => net108530);
   registers_reg_6_14_inst : DFFR_X1 port map( D => n3829, CK => n599, RN => 
                           rst, Q => registers_6_14_port, QN => net108529);
   registers_reg_6_13_inst : DFFR_X1 port map( D => n3828, CK => n602, RN => 
                           rst, Q => registers_6_13_port, QN => net108528);
   registers_reg_6_12_inst : DFFR_X1 port map( D => n3827, CK => n627, RN => 
                           rst, Q => registers_6_12_port, QN => net108527);
   registers_reg_6_11_inst : DFFR_X1 port map( D => n3826, CK => n593, RN => 
                           rst, Q => registers_6_11_port, QN => net108526);
   registers_reg_6_10_inst : DFFR_X1 port map( D => n3825, CK => n610, RN => 
                           rst, Q => registers_6_10_port, QN => net108525);
   registers_reg_6_9_inst : DFFR_X1 port map( D => n3824, CK => n589, RN => rst
                           , Q => registers_6_9_port, QN => net108524);
   registers_reg_6_8_inst : DFFR_X1 port map( D => n3823, CK => n562, RN => rst
                           , Q => registers_6_8_port, QN => net108523);
   registers_reg_6_7_inst : DFFR_X1 port map( D => n3822, CK => n546, RN => rst
                           , Q => registers_6_7_port, QN => net108522);
   registers_reg_6_6_inst : DFFR_X1 port map( D => n3821, CK => n596, RN => rst
                           , Q => registers_6_6_port, QN => net108521);
   registers_reg_6_5_inst : DFFR_X1 port map( D => n3820, CK => n581, RN => rst
                           , Q => registers_6_5_port, QN => net108520);
   registers_reg_6_4_inst : DFFR_X1 port map( D => n3819, CK => n620, RN => rst
                           , Q => registers_6_4_port, QN => net108519);
   registers_reg_6_3_inst : DFFR_X1 port map( D => n3818, CK => n613, RN => rst
                           , Q => registers_6_3_port, QN => net108518);
   registers_reg_6_2_inst : DFFR_X1 port map( D => n3817, CK => n608, RN => rst
                           , Q => registers_6_2_port, QN => net108517);
   registers_reg_6_1_inst : DFFR_X1 port map( D => n3816, CK => n614, RN => rst
                           , Q => registers_6_1_port, QN => net108516);
   registers_reg_6_0_inst : DFFR_X1 port map( D => n3815, CK => n580, RN => rst
                           , Q => registers_6_0_port, QN => net108515);
   registers_reg_7_31_inst : DFFR_X1 port map( D => n3814, CK => n568, RN => 
                           rst, Q => registers_7_31_port, QN => n162);
   registers_reg_7_30_inst : DFFR_X1 port map( D => n3813, CK => n571, RN => 
                           rst, Q => registers_7_30_port, QN => n98);
   registers_reg_7_29_inst : DFFR_X1 port map( D => n3812, CK => n574, RN => 
                           rst, Q => registers_7_29_port, QN => n100);
   registers_reg_7_28_inst : DFFR_X1 port map( D => n3811, CK => n577, RN => 
                           rst, Q => registers_7_28_port, QN => n102);
   registers_reg_7_27_inst : DFFR_X1 port map( D => n3810, CK => n584, RN => 
                           rst, Q => registers_7_27_port, QN => n104);
   registers_reg_7_26_inst : DFFR_X1 port map( D => n3809, CK => n549, RN => 
                           rst, Q => registers_7_26_port, QN => n106);
   registers_reg_7_25_inst : DFFR_X1 port map( D => n3808, CK => n564, RN => 
                           rst, Q => registers_7_25_port, QN => n108);
   registers_reg_7_24_inst : DFFR_X1 port map( D => n3807, CK => n586, RN => 
                           rst, Q => registers_7_24_port, QN => n110);
   registers_reg_7_23_inst : DFFR_X1 port map( D => n3806, CK => n552, RN => 
                           rst, Q => registers_7_23_port, QN => n112);
   registers_reg_7_22_inst : DFFR_X1 port map( D => n3805, CK => n567, RN => 
                           rst, Q => registers_7_22_port, QN => n114);
   registers_reg_7_21_inst : DFFR_X1 port map( D => n3804, CK => n622, RN => 
                           rst, Q => registers_7_21_port, QN => n116);
   registers_reg_7_20_inst : DFFR_X1 port map( D => n3803, CK => n555, RN => 
                           rst, Q => registers_7_20_port, QN => n118);
   registers_reg_7_19_inst : DFFR_X1 port map( D => n3802, CK => n617, RN => 
                           rst, Q => registers_7_19_port, QN => n120);
   registers_reg_7_18_inst : DFFR_X1 port map( D => n3801, CK => n568, RN => 
                           rst, Q => registers_7_18_port, QN => n122);
   registers_reg_7_17_inst : DFFR_X1 port map( D => n3800, CK => n629, RN => 
                           rst, Q => registers_7_17_port, QN => n124);
   registers_reg_7_16_inst : DFFR_X1 port map( D => n3799, CK => n633, RN => 
                           rst, Q => registers_7_16_port, QN => n126);
   registers_reg_7_15_inst : DFFR_X1 port map( D => n3798, CK => n559, RN => 
                           rst, Q => registers_7_15_port, QN => n128);
   registers_reg_7_14_inst : DFFR_X1 port map( D => n3797, CK => n599, RN => 
                           rst, Q => registers_7_14_port, QN => n130);
   registers_reg_7_13_inst : DFFR_X1 port map( D => n3796, CK => n602, RN => 
                           rst, Q => registers_7_13_port, QN => n132);
   registers_reg_7_12_inst : DFFR_X1 port map( D => n3795, CK => n627, RN => 
                           rst, Q => registers_7_12_port, QN => n134);
   registers_reg_7_11_inst : DFFR_X1 port map( D => n3794, CK => n593, RN => 
                           rst, Q => registers_7_11_port, QN => n136);
   registers_reg_7_10_inst : DFFR_X1 port map( D => n3793, CK => n610, RN => 
                           rst, Q => registers_7_10_port, QN => n138);
   registers_reg_7_9_inst : DFFR_X1 port map( D => n3792, CK => n589, RN => rst
                           , Q => registers_7_9_port, QN => n140);
   registers_reg_7_8_inst : DFFR_X1 port map( D => n3791, CK => n562, RN => rst
                           , Q => registers_7_8_port, QN => n142);
   registers_reg_7_7_inst : DFFR_X1 port map( D => n3790, CK => n546, RN => rst
                           , Q => registers_7_7_port, QN => n144);
   registers_reg_7_6_inst : DFFR_X1 port map( D => n3789, CK => n596, RN => rst
                           , Q => registers_7_6_port, QN => n146);
   registers_reg_7_5_inst : DFFR_X1 port map( D => n3788, CK => n581, RN => rst
                           , Q => registers_7_5_port, QN => n148);
   registers_reg_7_4_inst : DFFR_X1 port map( D => n3787, CK => n620, RN => rst
                           , Q => registers_7_4_port, QN => n150);
   registers_reg_7_3_inst : DFFR_X1 port map( D => n3786, CK => n613, RN => rst
                           , Q => registers_7_3_port, QN => n152);
   registers_reg_7_2_inst : DFFR_X1 port map( D => n3785, CK => n607, RN => rst
                           , Q => registers_7_2_port, QN => n154);
   registers_reg_7_1_inst : DFFR_X1 port map( D => n3784, CK => n614, RN => rst
                           , Q => registers_7_1_port, QN => n156);
   registers_reg_7_0_inst : DFFR_X1 port map( D => n3783, CK => n579, RN => rst
                           , Q => registers_7_0_port, QN => n158);
   registers_reg_8_31_inst : DFFR_X1 port map( D => n3782, CK => n568, RN => 
                           rst, Q => registers_8_31_port, QN => n65);
   registers_reg_8_30_inst : DFFR_X1 port map( D => n3781, CK => n571, RN => 
                           rst, Q => registers_8_30_port, QN => n66);
   registers_reg_8_29_inst : DFFR_X1 port map( D => n3780, CK => n574, RN => 
                           rst, Q => registers_8_29_port, QN => n67);
   registers_reg_8_28_inst : DFFR_X1 port map( D => n3779, CK => n576, RN => 
                           rst, Q => registers_8_28_port, QN => n68);
   registers_reg_8_27_inst : DFFR_X1 port map( D => n3778, CK => n583, RN => 
                           rst, Q => registers_8_27_port, QN => n69);
   registers_reg_8_26_inst : DFFR_X1 port map( D => n3777, CK => n549, RN => 
                           rst, Q => registers_8_26_port, QN => n70);
   registers_reg_8_25_inst : DFFR_X1 port map( D => n3776, CK => n564, RN => 
                           rst, Q => registers_8_25_port, QN => n71);
   registers_reg_8_24_inst : DFFR_X1 port map( D => n3775, CK => n586, RN => 
                           rst, Q => registers_8_24_port, QN => n72);
   registers_reg_8_23_inst : DFFR_X1 port map( D => n3774, CK => n552, RN => 
                           rst, Q => registers_8_23_port, QN => n73);
   registers_reg_8_22_inst : DFFR_X1 port map( D => n3773, CK => n567, RN => 
                           rst, Q => registers_8_22_port, QN => n74);
   registers_reg_8_21_inst : DFFR_X1 port map( D => n3772, CK => n622, RN => 
                           rst, Q => registers_8_21_port, QN => n75);
   registers_reg_8_20_inst : DFFR_X1 port map( D => n3771, CK => n555, RN => 
                           rst, Q => registers_8_20_port, QN => n76);
   registers_reg_8_19_inst : DFFR_X1 port map( D => n3770, CK => n617, RN => 
                           rst, Q => registers_8_19_port, QN => n77);
   registers_reg_8_18_inst : DFFR_X1 port map( D => n3769, CK => n625, RN => 
                           rst, Q => registers_8_18_port, QN => n78);
   registers_reg_8_17_inst : DFFR_X1 port map( D => n3768, CK => n629, RN => 
                           rst, Q => registers_8_17_port, QN => n79);
   registers_reg_8_16_inst : DFFR_X1 port map( D => n3767, CK => n632, RN => 
                           rst, Q => registers_8_16_port, QN => n80);
   registers_reg_8_15_inst : DFFR_X1 port map( D => n3766, CK => n559, RN => 
                           rst, Q => registers_8_15_port, QN => n81);
   registers_reg_8_14_inst : DFFR_X1 port map( D => n3765, CK => n599, RN => 
                           rst, Q => registers_8_14_port, QN => n82);
   registers_reg_8_13_inst : DFFR_X1 port map( D => n3764, CK => n602, RN => 
                           rst, Q => registers_8_13_port, QN => n83);
   registers_reg_8_12_inst : DFFR_X1 port map( D => n3763, CK => n626, RN => 
                           rst, Q => registers_8_12_port, QN => n84);
   registers_reg_8_11_inst : DFFR_X1 port map( D => n3762, CK => n593, RN => 
                           rst, Q => registers_8_11_port, QN => n85);
   registers_reg_8_10_inst : DFFR_X1 port map( D => n3761, CK => n610, RN => 
                           rst, Q => registers_8_10_port, QN => n86);
   registers_reg_8_9_inst : DFFR_X1 port map( D => n3760, CK => n589, RN => rst
                           , Q => registers_8_9_port, QN => n87);
   registers_reg_8_8_inst : DFFR_X1 port map( D => n3759, CK => n562, RN => rst
                           , Q => registers_8_8_port, QN => n88);
   registers_reg_8_7_inst : DFFR_X1 port map( D => n3758, CK => n546, RN => rst
                           , Q => registers_8_7_port, QN => n89);
   registers_reg_8_6_inst : DFFR_X1 port map( D => n3757, CK => n596, RN => rst
                           , Q => registers_8_6_port, QN => n90);
   registers_reg_8_5_inst : DFFR_X1 port map( D => n3756, CK => n581, RN => rst
                           , Q => registers_8_5_port, QN => n91);
   registers_reg_8_4_inst : DFFR_X1 port map( D => n3755, CK => n620, RN => rst
                           , Q => registers_8_4_port, QN => n92);
   registers_reg_8_3_inst : DFFR_X1 port map( D => n3754, CK => n613, RN => rst
                           , Q => registers_8_3_port, QN => n93);
   registers_reg_8_2_inst : DFFR_X1 port map( D => n3753, CK => n607, RN => rst
                           , Q => registers_8_2_port, QN => n94);
   registers_reg_8_1_inst : DFFR_X1 port map( D => n3752, CK => n614, RN => rst
                           , Q => registers_8_1_port, QN => n95);
   registers_reg_8_0_inst : DFFR_X1 port map( D => n3751, CK => n579, RN => rst
                           , Q => registers_8_0_port, QN => n96);
   registers_reg_9_31_inst : DFFR_X1 port map( D => n3750, CK => n574, RN => 
                           rst, Q => registers_9_31_port, QN => net108514);
   registers_reg_9_30_inst : DFFR_X1 port map( D => n3749, CK => n571, RN => 
                           rst, Q => registers_9_30_port, QN => net108513);
   registers_reg_9_29_inst : DFFR_X1 port map( D => n3748, CK => n574, RN => 
                           rst, Q => registers_9_29_port, QN => net108512);
   registers_reg_9_28_inst : DFFR_X1 port map( D => n3747, CK => n576, RN => 
                           rst, Q => registers_9_28_port, QN => net108511);
   registers_reg_9_27_inst : DFFR_X1 port map( D => n3746, CK => n583, RN => 
                           rst, Q => registers_9_27_port, QN => net108510);
   registers_reg_9_26_inst : DFFR_X1 port map( D => n3745, CK => n549, RN => 
                           rst, Q => registers_9_26_port, QN => net108509);
   registers_reg_9_25_inst : DFFR_X1 port map( D => n3744, CK => n564, RN => 
                           rst, Q => registers_9_25_port, QN => net108508);
   registers_reg_9_24_inst : DFFR_X1 port map( D => n3743, CK => n586, RN => 
                           rst, Q => registers_9_24_port, QN => net108507);
   registers_reg_9_23_inst : DFFR_X1 port map( D => n3742, CK => n552, RN => 
                           rst, Q => registers_9_23_port, QN => net108506);
   registers_reg_9_22_inst : DFFR_X1 port map( D => n3741, CK => n567, RN => 
                           rst, Q => registers_9_22_port, QN => net108505);
   registers_reg_9_21_inst : DFFR_X1 port map( D => n3740, CK => n622, RN => 
                           rst, Q => registers_9_21_port, QN => net108504);
   registers_reg_9_20_inst : DFFR_X1 port map( D => n3739, CK => n554, RN => 
                           rst, Q => registers_9_20_port, QN => net108503);
   registers_reg_9_19_inst : DFFR_X1 port map( D => n3738, CK => n617, RN => 
                           rst, Q => registers_9_19_port, QN => net108502);
   registers_reg_9_18_inst : DFFR_X1 port map( D => n3737, CK => n625, RN => 
                           rst, Q => registers_9_18_port, QN => net108501);
   registers_reg_9_17_inst : DFFR_X1 port map( D => n3736, CK => n629, RN => 
                           rst, Q => registers_9_17_port, QN => net108500);
   registers_reg_9_16_inst : DFFR_X1 port map( D => n3735, CK => n633, RN => 
                           rst, Q => registers_9_16_port, QN => net108499);
   registers_reg_9_15_inst : DFFR_X1 port map( D => n3734, CK => n559, RN => 
                           rst, Q => registers_9_15_port, QN => net108498);
   registers_reg_9_14_inst : DFFR_X1 port map( D => n3733, CK => n599, RN => 
                           rst, Q => registers_9_14_port, QN => net108497);
   registers_reg_9_13_inst : DFFR_X1 port map( D => n3732, CK => n601, RN => 
                           rst, Q => registers_9_13_port, QN => net108496);
   registers_reg_9_12_inst : DFFR_X1 port map( D => n3731, CK => n626, RN => 
                           rst, Q => registers_9_12_port, QN => net108495);
   registers_reg_9_11_inst : DFFR_X1 port map( D => n3730, CK => n593, RN => 
                           rst, Q => registers_9_11_port, QN => net108494);
   registers_reg_9_10_inst : DFFR_X1 port map( D => n3729, CK => n610, RN => 
                           rst, Q => registers_9_10_port, QN => net108493);
   registers_reg_9_9_inst : DFFR_X1 port map( D => n3728, CK => n589, RN => rst
                           , Q => registers_9_9_port, QN => net108492);
   registers_reg_9_8_inst : DFFR_X1 port map( D => n3727, CK => n561, RN => rst
                           , Q => registers_9_8_port, QN => net108491);
   registers_reg_9_7_inst : DFFR_X1 port map( D => n3726, CK => n546, RN => rst
                           , Q => registers_9_7_port, QN => net108490);
   registers_reg_9_6_inst : DFFR_X1 port map( D => n3725, CK => n596, RN => rst
                           , Q => registers_9_6_port, QN => net108489);
   registers_reg_9_5_inst : DFFR_X1 port map( D => n3724, CK => n581, RN => rst
                           , Q => registers_9_5_port, QN => net108488);
   registers_reg_9_4_inst : DFFR_X1 port map( D => n3723, CK => n619, RN => rst
                           , Q => registers_9_4_port, QN => net108487);
   registers_reg_9_3_inst : DFFR_X1 port map( D => n3722, CK => n613, RN => rst
                           , Q => registers_9_3_port, QN => net108486);
   registers_reg_9_2_inst : DFFR_X1 port map( D => n3721, CK => n607, RN => rst
                           , Q => registers_9_2_port, QN => net108485);
   registers_reg_9_1_inst : DFFR_X1 port map( D => n3720, CK => n619, RN => rst
                           , Q => registers_9_1_port, QN => net108484);
   registers_reg_9_0_inst : DFFR_X1 port map( D => n3719, CK => n579, RN => rst
                           , Q => registers_9_0_port, QN => net108483);
   registers_reg_10_31_inst : DFFR_X1 port map( D => n3718, CK => n592, RN => 
                           rst, Q => registers_10_31_port, QN => n544);
   registers_reg_10_30_inst : DFFR_X1 port map( D => n3717, CK => n571, RN => 
                           rst, Q => registers_10_30_port, QN => n354);
   registers_reg_10_29_inst : DFFR_X1 port map( D => n3716, CK => n573, RN => 
                           rst, Q => registers_10_29_port, QN => n356);
   registers_reg_10_28_inst : DFFR_X1 port map( D => n3715, CK => n576, RN => 
                           rst, Q => registers_10_28_port, QN => n358);
   registers_reg_10_27_inst : DFFR_X1 port map( D => n3714, CK => n583, RN => 
                           rst, Q => registers_10_27_port, QN => n360);
   registers_reg_10_26_inst : DFFR_X1 port map( D => n3713, CK => n549, RN => 
                           rst, Q => registers_10_26_port, QN => n362);
   registers_reg_10_25_inst : DFFR_X1 port map( D => n3712, CK => n564, RN => 
                           rst, Q => registers_10_25_port, QN => n364);
   registers_reg_10_24_inst : DFFR_X1 port map( D => n3711, CK => n586, RN => 
                           rst, Q => registers_10_24_port, QN => n366);
   registers_reg_10_23_inst : DFFR_X1 port map( D => n3710, CK => n552, RN => 
                           rst, Q => registers_10_23_port, QN => n368);
   registers_reg_10_22_inst : DFFR_X1 port map( D => n3709, CK => n567, RN => 
                           rst, Q => registers_10_22_port, QN => n370);
   registers_reg_10_21_inst : DFFR_X1 port map( D => n3708, CK => n622, RN => 
                           rst, Q => registers_10_21_port, QN => n372);
   registers_reg_10_20_inst : DFFR_X1 port map( D => n3707, CK => n554, RN => 
                           rst, Q => registers_10_20_port, QN => n374);
   registers_reg_10_19_inst : DFFR_X1 port map( D => n3706, CK => n617, RN => 
                           rst, Q => registers_10_19_port, QN => n376);
   registers_reg_10_18_inst : DFFR_X1 port map( D => n3705, CK => n625, RN => 
                           rst, Q => registers_10_18_port, QN => n378);
   registers_reg_10_17_inst : DFFR_X1 port map( D => n3704, CK => n629, RN => 
                           rst, Q => registers_10_17_port, QN => n380);
   registers_reg_10_16_inst : DFFR_X1 port map( D => n3703, CK => n633, RN => 
                           rst, Q => registers_10_16_port, QN => n382);
   registers_reg_10_15_inst : DFFR_X1 port map( D => n3702, CK => n559, RN => 
                           rst, Q => registers_10_15_port, QN => n384);
   registers_reg_10_14_inst : DFFR_X1 port map( D => n3701, CK => n599, RN => 
                           rst, Q => registers_10_14_port, QN => n386);
   registers_reg_10_13_inst : DFFR_X1 port map( D => n3700, CK => n601, RN => 
                           rst, Q => registers_10_13_port, QN => n388);
   registers_reg_10_12_inst : DFFR_X1 port map( D => n3699, CK => n626, RN => 
                           rst, Q => registers_10_12_port, QN => n390);
   registers_reg_10_11_inst : DFFR_X1 port map( D => n3698, CK => n593, RN => 
                           rst, Q => registers_10_11_port, QN => n392);
   registers_reg_10_10_inst : DFFR_X1 port map( D => n3697, CK => n610, RN => 
                           rst, Q => registers_10_10_port, QN => n394);
   registers_reg_10_9_inst : DFFR_X1 port map( D => n3696, CK => n589, RN => 
                           rst, Q => registers_10_9_port, QN => n396);
   registers_reg_10_8_inst : DFFR_X1 port map( D => n3695, CK => n561, RN => 
                           rst, Q => registers_10_8_port, QN => n398);
   registers_reg_10_7_inst : DFFR_X1 port map( D => n3694, CK => n546, RN => 
                           rst, Q => registers_10_7_port, QN => n400);
   registers_reg_10_6_inst : DFFR_X1 port map( D => n3693, CK => n596, RN => 
                           rst, Q => registers_10_6_port, QN => n402);
   registers_reg_10_5_inst : DFFR_X1 port map( D => n3692, CK => n581, RN => 
                           rst, Q => registers_10_5_port, QN => n404);
   registers_reg_10_4_inst : DFFR_X1 port map( D => n3691, CK => n619, RN => 
                           rst, Q => registers_10_4_port, QN => n406);
   registers_reg_10_3_inst : DFFR_X1 port map( D => n3690, CK => n613, RN => 
                           rst, Q => registers_10_3_port, QN => n408);
   registers_reg_10_2_inst : DFFR_X1 port map( D => n3689, CK => n607, RN => 
                           rst, Q => registers_10_2_port, QN => n410);
   registers_reg_10_1_inst : DFFR_X1 port map( D => n3688, CK => n631, RN => 
                           rst, Q => registers_10_1_port, QN => n412);
   registers_reg_10_0_inst : DFFR_X1 port map( D => n3687, CK => n579, RN => 
                           rst, Q => registers_10_0_port, QN => n414);
   registers_reg_11_31_inst : DFFR_X1 port map( D => n3686, CK => n591, RN => 
                           rst, Q => registers_11_31_port, QN => net108482);
   registers_reg_11_30_inst : DFFR_X1 port map( D => n3685, CK => n571, RN => 
                           rst, Q => registers_11_30_port, QN => net108481);
   registers_reg_11_29_inst : DFFR_X1 port map( D => n3684, CK => n573, RN => 
                           rst, Q => registers_11_29_port, QN => net108480);
   registers_reg_11_28_inst : DFFR_X1 port map( D => n3683, CK => n576, RN => 
                           rst, Q => registers_11_28_port, QN => net108479);
   registers_reg_11_27_inst : DFFR_X1 port map( D => n3682, CK => n583, RN => 
                           rst, Q => registers_11_27_port, QN => net108478);
   registers_reg_11_26_inst : DFFR_X1 port map( D => n3681, CK => n549, RN => 
                           rst, Q => registers_11_26_port, QN => net108477);
   registers_reg_11_25_inst : DFFR_X1 port map( D => n3680, CK => n564, RN => 
                           rst, Q => registers_11_25_port, QN => net108476);
   registers_reg_11_24_inst : DFFR_X1 port map( D => n3679, CK => n586, RN => 
                           rst, Q => registers_11_24_port, QN => net108475);
   registers_reg_11_23_inst : DFFR_X1 port map( D => n3678, CK => n552, RN => 
                           rst, Q => registers_11_23_port, QN => net108474);
   registers_reg_11_22_inst : DFFR_X1 port map( D => n3677, CK => n567, RN => 
                           rst, Q => registers_11_22_port, QN => net108473);
   registers_reg_11_21_inst : DFFR_X1 port map( D => n3676, CK => n622, RN => 
                           rst, Q => registers_11_21_port, QN => net108472);
   registers_reg_11_20_inst : DFFR_X1 port map( D => n3675, CK => n554, RN => 
                           rst, Q => registers_11_20_port, QN => net108471);
   registers_reg_11_19_inst : DFFR_X1 port map( D => n3674, CK => n616, RN => 
                           rst, Q => registers_11_19_port, QN => net108470);
   registers_reg_11_18_inst : DFFR_X1 port map( D => n3673, CK => n625, RN => 
                           rst, Q => registers_11_18_port, QN => net108469);
   registers_reg_11_17_inst : DFFR_X1 port map( D => n3672, CK => n629, RN => 
                           rst, Q => registers_11_17_port, QN => net108468);
   registers_reg_11_16_inst : DFFR_X1 port map( D => n3671, CK => n632, RN => 
                           rst, Q => registers_11_16_port, QN => net108467);
   registers_reg_11_15_inst : DFFR_X1 port map( D => n3670, CK => n559, RN => 
                           rst, Q => registers_11_15_port, QN => net108466);
   registers_reg_11_14_inst : DFFR_X1 port map( D => n3669, CK => n599, RN => 
                           rst, Q => registers_11_14_port, QN => net108465);
   registers_reg_11_13_inst : DFFR_X1 port map( D => n3668, CK => n601, RN => 
                           rst, Q => registers_11_13_port, QN => net108464);
   registers_reg_11_12_inst : DFFR_X1 port map( D => n3667, CK => n626, RN => 
                           rst, Q => registers_11_12_port, QN => net108463);
   registers_reg_11_11_inst : DFFR_X1 port map( D => n3666, CK => n593, RN => 
                           rst, Q => registers_11_11_port, QN => net108462);
   registers_reg_11_10_inst : DFFR_X1 port map( D => n3665, CK => n610, RN => 
                           rst, Q => registers_11_10_port, QN => net108461);
   registers_reg_11_9_inst : DFFR_X1 port map( D => n3664, CK => n589, RN => 
                           rst, Q => registers_11_9_port, QN => net108460);
   registers_reg_11_8_inst : DFFR_X1 port map( D => n3663, CK => n561, RN => 
                           rst, Q => registers_11_8_port, QN => net108459);
   registers_reg_11_7_inst : DFFR_X1 port map( D => n3662, CK => n546, RN => 
                           rst, Q => registers_11_7_port, QN => net108458);
   registers_reg_11_6_inst : DFFR_X1 port map( D => n3661, CK => n596, RN => 
                           rst, Q => registers_11_6_port, QN => net108457);
   registers_reg_11_5_inst : DFFR_X1 port map( D => n3660, CK => n580, RN => 
                           rst, Q => registers_11_5_port, QN => net108456);
   registers_reg_11_4_inst : DFFR_X1 port map( D => n3659, CK => n619, RN => 
                           rst, Q => registers_11_4_port, QN => net108455);
   registers_reg_11_3_inst : DFFR_X1 port map( D => n3658, CK => n613, RN => 
                           rst, Q => registers_11_3_port, QN => net108454);
   registers_reg_11_2_inst : DFFR_X1 port map( D => n3657, CK => n607, RN => 
                           rst, Q => registers_11_2_port, QN => net108453);
   registers_reg_11_1_inst : DFFR_X1 port map( D => n3656, CK => n631, RN => 
                           rst, Q => registers_11_1_port, QN => net108452);
   registers_reg_11_0_inst : DFFR_X1 port map( D => n3655, CK => n579, RN => 
                           rst, Q => registers_11_0_port, QN => net108451);
   registers_reg_12_31_inst : DFFR_X1 port map( D => n3654, CK => n591, RN => 
                           rst, Q => registers_12_31_port, QN => net108450);
   registers_reg_12_30_inst : DFFR_X1 port map( D => n3653, CK => n571, RN => 
                           rst, Q => registers_12_30_port, QN => net108449);
   registers_reg_12_29_inst : DFFR_X1 port map( D => n3652, CK => n573, RN => 
                           rst, Q => registers_12_29_port, QN => net108448);
   registers_reg_12_28_inst : DFFR_X1 port map( D => n3651, CK => n576, RN => 
                           rst, Q => registers_12_28_port, QN => net108447);
   registers_reg_12_27_inst : DFFR_X1 port map( D => n3650, CK => n583, RN => 
                           rst, Q => registers_12_27_port, QN => net108446);
   registers_reg_12_26_inst : DFFR_X1 port map( D => n3649, CK => n549, RN => 
                           rst, Q => registers_12_26_port, QN => net108445);
   registers_reg_12_25_inst : DFFR_X1 port map( D => n3648, CK => n564, RN => 
                           rst, Q => registers_12_25_port, QN => net108444);
   registers_reg_12_24_inst : DFFR_X1 port map( D => n3647, CK => n586, RN => 
                           rst, Q => registers_12_24_port, QN => net108443);
   registers_reg_12_23_inst : DFFR_X1 port map( D => n3646, CK => n551, RN => 
                           rst, Q => registers_12_23_port, QN => net108442);
   registers_reg_12_22_inst : DFFR_X1 port map( D => n3645, CK => n567, RN => 
                           rst, Q => registers_12_22_port, QN => net108441);
   registers_reg_12_21_inst : DFFR_X1 port map( D => n3644, CK => n622, RN => 
                           rst, Q => registers_12_21_port, QN => net108440);
   registers_reg_12_20_inst : DFFR_X1 port map( D => n3643, CK => n554, RN => 
                           rst, Q => registers_12_20_port, QN => net108439);
   registers_reg_12_19_inst : DFFR_X1 port map( D => n3642, CK => n616, RN => 
                           rst, Q => registers_12_19_port, QN => net108438);
   registers_reg_12_18_inst : DFFR_X1 port map( D => n3641, CK => n625, RN => 
                           rst, Q => registers_12_18_port, QN => net108437);
   registers_reg_12_17_inst : DFFR_X1 port map( D => n3640, CK => n629, RN => 
                           rst, Q => registers_12_17_port, QN => net108436);
   registers_reg_12_16_inst : DFFR_X1 port map( D => n3639, CK => n632, RN => 
                           rst, Q => registers_12_16_port, QN => net108435);
   registers_reg_12_15_inst : DFFR_X1 port map( D => n3638, CK => n558, RN => 
                           rst, Q => registers_12_15_port, QN => net108434);
   registers_reg_12_14_inst : DFFR_X1 port map( D => n3637, CK => n598, RN => 
                           rst, Q => registers_12_14_port, QN => net108433);
   registers_reg_12_13_inst : DFFR_X1 port map( D => n3636, CK => n601, RN => 
                           rst, Q => registers_12_13_port, QN => net108432);
   registers_reg_12_12_inst : DFFR_X1 port map( D => n3635, CK => n626, RN => 
                           rst, Q => registers_12_12_port, QN => net108431);
   registers_reg_12_11_inst : DFFR_X1 port map( D => n3634, CK => n593, RN => 
                           rst, Q => registers_12_11_port, QN => net108430);
   registers_reg_12_10_inst : DFFR_X1 port map( D => n3633, CK => n610, RN => 
                           rst, Q => registers_12_10_port, QN => net108429);
   registers_reg_12_9_inst : DFFR_X1 port map( D => n3632, CK => n589, RN => 
                           rst, Q => registers_12_9_port, QN => net108428);
   registers_reg_12_8_inst : DFFR_X1 port map( D => n3631, CK => n561, RN => 
                           rst, Q => registers_12_8_port, QN => net108427);
   registers_reg_12_7_inst : DFFR_X1 port map( D => n3630, CK => n546, RN => 
                           rst, Q => registers_12_7_port, QN => net108426);
   registers_reg_12_6_inst : DFFR_X1 port map( D => n3629, CK => n596, RN => 
                           rst, Q => registers_12_6_port, QN => net108425);
   registers_reg_12_5_inst : DFFR_X1 port map( D => n3628, CK => n580, RN => 
                           rst, Q => registers_12_5_port, QN => net108424);
   registers_reg_12_4_inst : DFFR_X1 port map( D => n3627, CK => n619, RN => 
                           rst, Q => registers_12_4_port, QN => net108423);
   registers_reg_12_3_inst : DFFR_X1 port map( D => n3626, CK => n612, RN => 
                           rst, Q => registers_12_3_port, QN => net108422);
   registers_reg_12_2_inst : DFFR_X1 port map( D => n3625, CK => n607, RN => 
                           rst, Q => registers_12_2_port, QN => net108421);
   registers_reg_12_1_inst : DFFR_X1 port map( D => n3624, CK => n632, RN => 
                           rst, Q => registers_12_1_port, QN => net108420);
   registers_reg_12_0_inst : DFFR_X1 port map( D => n3623, CK => n579, RN => 
                           rst, Q => registers_12_0_port, QN => net108419);
   registers_reg_13_31_inst : DFFR_X1 port map( D => n3622, CK => n591, RN => 
                           rst, Q => registers_13_31_port, QN => n415);
   registers_reg_13_30_inst : DFFR_X1 port map( D => n3621, CK => n570, RN => 
                           rst, Q => registers_13_30_port, QN => n417);
   registers_reg_13_29_inst : DFFR_X1 port map( D => n3620, CK => n573, RN => 
                           rst, Q => registers_13_29_port, QN => n419);
   registers_reg_13_28_inst : DFFR_X1 port map( D => n3619, CK => n576, RN => 
                           rst, Q => registers_13_28_port, QN => n421);
   registers_reg_13_27_inst : DFFR_X1 port map( D => n3618, CK => n583, RN => 
                           rst, Q => registers_13_27_port, QN => n423);
   registers_reg_13_26_inst : DFFR_X1 port map( D => n3617, CK => n549, RN => 
                           rst, Q => registers_13_26_port, QN => n425);
   registers_reg_13_25_inst : DFFR_X1 port map( D => n3616, CK => n564, RN => 
                           rst, Q => registers_13_25_port, QN => n427);
   registers_reg_13_24_inst : DFFR_X1 port map( D => n3615, CK => n586, RN => 
                           rst, Q => registers_13_24_port, QN => n429);
   registers_reg_13_23_inst : DFFR_X1 port map( D => n3614, CK => n551, RN => 
                           rst, Q => registers_13_23_port, QN => n431);
   registers_reg_13_22_inst : DFFR_X1 port map( D => n3613, CK => n567, RN => 
                           rst, Q => registers_13_22_port, QN => n433);
   registers_reg_13_21_inst : DFFR_X1 port map( D => n3612, CK => n622, RN => 
                           rst, Q => registers_13_21_port, QN => n435);
   registers_reg_13_20_inst : DFFR_X1 port map( D => n3611, CK => n554, RN => 
                           rst, Q => registers_13_20_port, QN => n437);
   registers_reg_13_19_inst : DFFR_X1 port map( D => n3610, CK => n616, RN => 
                           rst, Q => registers_13_19_port, QN => n439);
   registers_reg_13_18_inst : DFFR_X1 port map( D => n3609, CK => n625, RN => 
                           rst, Q => registers_13_18_port, QN => n441);
   registers_reg_13_17_inst : DFFR_X1 port map( D => n3608, CK => n629, RN => 
                           rst, Q => registers_13_17_port, QN => n443);
   registers_reg_13_16_inst : DFFR_X1 port map( D => n3607, CK => n632, RN => 
                           rst, Q => registers_13_16_port, QN => n445);
   registers_reg_13_15_inst : DFFR_X1 port map( D => n3606, CK => n558, RN => 
                           rst, Q => registers_13_15_port, QN => n447);
   registers_reg_13_14_inst : DFFR_X1 port map( D => n3605, CK => n598, RN => 
                           rst, Q => registers_13_14_port, QN => n449);
   registers_reg_13_13_inst : DFFR_X1 port map( D => n3604, CK => n601, RN => 
                           rst, Q => registers_13_13_port, QN => n451);
   registers_reg_13_12_inst : DFFR_X1 port map( D => n3603, CK => n626, RN => 
                           rst, Q => registers_13_12_port, QN => n453);
   registers_reg_13_11_inst : DFFR_X1 port map( D => n3602, CK => n593, RN => 
                           rst, Q => registers_13_11_port, QN => n455);
   registers_reg_13_10_inst : DFFR_X1 port map( D => n3601, CK => n610, RN => 
                           rst, Q => registers_13_10_port, QN => n457);
   registers_reg_13_9_inst : DFFR_X1 port map( D => n3600, CK => n589, RN => 
                           rst, Q => registers_13_9_port, QN => n459);
   registers_reg_13_8_inst : DFFR_X1 port map( D => n3599, CK => n561, RN => 
                           rst, Q => registers_13_8_port, QN => n461);
   registers_reg_13_7_inst : DFFR_X1 port map( D => n3598, CK => n546, RN => 
                           rst, Q => registers_13_7_port, QN => n463);
   registers_reg_13_6_inst : DFFR_X1 port map( D => n3597, CK => n596, RN => 
                           rst, Q => registers_13_6_port, QN => n465);
   registers_reg_13_5_inst : DFFR_X1 port map( D => n3596, CK => n580, RN => 
                           rst, Q => registers_13_5_port, QN => n467);
   registers_reg_13_4_inst : DFFR_X1 port map( D => n3595, CK => n619, RN => 
                           rst, Q => registers_13_4_port, QN => n469);
   registers_reg_13_3_inst : DFFR_X1 port map( D => n3594, CK => n612, RN => 
                           rst, Q => registers_13_3_port, QN => n471);
   registers_reg_13_2_inst : DFFR_X1 port map( D => n3593, CK => n607, RN => 
                           rst, Q => registers_13_2_port, QN => n473);
   registers_reg_13_1_inst : DFFR_X1 port map( D => n3592, CK => n632, RN => 
                           rst, Q => registers_13_1_port, QN => n475);
   registers_reg_13_0_inst : DFFR_X1 port map( D => n3591, CK => n579, RN => 
                           rst, Q => registers_13_0_port, QN => n477);
   registers_reg_14_31_inst : DFFR_X1 port map( D => n3590, CK => n591, RN => 
                           rst, Q => registers_14_31_port, QN => net108418);
   registers_reg_14_30_inst : DFFR_X1 port map( D => n3589, CK => n570, RN => 
                           rst, Q => registers_14_30_port, QN => net108417);
   registers_reg_14_29_inst : DFFR_X1 port map( D => n3588, CK => n573, RN => 
                           rst, Q => registers_14_29_port, QN => net108416);
   registers_reg_14_28_inst : DFFR_X1 port map( D => n3587, CK => n576, RN => 
                           rst, Q => registers_14_28_port, QN => net108415);
   registers_reg_14_27_inst : DFFR_X1 port map( D => n3586, CK => n583, RN => 
                           rst, Q => registers_14_27_port, QN => net108414);
   registers_reg_14_26_inst : DFFR_X1 port map( D => n3585, CK => n548, RN => 
                           rst, Q => registers_14_26_port, QN => net108413);
   registers_reg_14_25_inst : DFFR_X1 port map( D => n3584, CK => n564, RN => 
                           rst, Q => registers_14_25_port, QN => net108412);
   registers_reg_14_24_inst : DFFR_X1 port map( D => n3583, CK => n586, RN => 
                           rst, Q => registers_14_24_port, QN => net108411);
   registers_reg_14_23_inst : DFFR_X1 port map( D => n3582, CK => n551, RN => 
                           rst, Q => registers_14_23_port, QN => net108410);
   registers_reg_14_22_inst : DFFR_X1 port map( D => n3581, CK => n567, RN => 
                           rst, Q => registers_14_22_port, QN => net108409);
   registers_reg_14_21_inst : DFFR_X1 port map( D => n3580, CK => n622, RN => 
                           rst, Q => registers_14_21_port, QN => net108408);
   registers_reg_14_20_inst : DFFR_X1 port map( D => n3579, CK => n554, RN => 
                           rst, Q => registers_14_20_port, QN => net108407);
   registers_reg_14_19_inst : DFFR_X1 port map( D => n3578, CK => n616, RN => 
                           rst, Q => registers_14_19_port, QN => net108406);
   registers_reg_14_18_inst : DFFR_X1 port map( D => n3577, CK => n624, RN => 
                           rst, Q => registers_14_18_port, QN => net108405);
   registers_reg_14_17_inst : DFFR_X1 port map( D => n3576, CK => n629, RN => 
                           rst, Q => registers_14_17_port, QN => net108404);
   registers_reg_14_16_inst : DFFR_X1 port map( D => n3575, CK => n631, RN => 
                           rst, Q => registers_14_16_port, QN => net108403);
   registers_reg_14_15_inst : DFFR_X1 port map( D => n3574, CK => n558, RN => 
                           rst, Q => registers_14_15_port, QN => net108402);
   registers_reg_14_14_inst : DFFR_X1 port map( D => n3573, CK => n598, RN => 
                           rst, Q => registers_14_14_port, QN => net108401);
   registers_reg_14_13_inst : DFFR_X1 port map( D => n3572, CK => n601, RN => 
                           rst, Q => registers_14_13_port, QN => net108400);
   registers_reg_14_12_inst : DFFR_X1 port map( D => n3571, CK => n626, RN => 
                           rst, Q => registers_14_12_port, QN => net108399);
   registers_reg_14_11_inst : DFFR_X1 port map( D => n3570, CK => n593, RN => 
                           rst, Q => registers_14_11_port, QN => net108398);
   registers_reg_14_10_inst : DFFR_X1 port map( D => n3569, CK => n610, RN => 
                           rst, Q => registers_14_10_port, QN => net108397);
   registers_reg_14_9_inst : DFFR_X1 port map( D => n3568, CK => n588, RN => 
                           rst, Q => registers_14_9_port, QN => net108396);
   registers_reg_14_8_inst : DFFR_X1 port map( D => n3567, CK => n561, RN => 
                           rst, Q => registers_14_8_port, QN => net108395);
   registers_reg_14_7_inst : DFFR_X1 port map( D => n3566, CK => n546, RN => 
                           rst, Q => registers_14_7_port, QN => net108394);
   registers_reg_14_6_inst : DFFR_X1 port map( D => n3565, CK => n595, RN => 
                           rst, Q => registers_14_6_port, QN => net108393);
   registers_reg_14_5_inst : DFFR_X1 port map( D => n3564, CK => n580, RN => 
                           rst, Q => registers_14_5_port, QN => net108392);
   registers_reg_14_4_inst : DFFR_X1 port map( D => n3563, CK => n619, RN => 
                           rst, Q => registers_14_4_port, QN => net108391);
   registers_reg_14_3_inst : DFFR_X1 port map( D => n3562, CK => n612, RN => 
                           rst, Q => registers_14_3_port, QN => net108390);
   registers_reg_14_2_inst : DFFR_X1 port map( D => n3561, CK => n607, RN => 
                           rst, Q => registers_14_2_port, QN => net108389);
   registers_reg_14_1_inst : DFFR_X1 port map( D => n3560, CK => n633, RN => 
                           rst, Q => registers_14_1_port, QN => net108388);
   registers_reg_14_0_inst : DFFR_X1 port map( D => n3559, CK => n579, RN => 
                           rst, Q => registers_14_0_port, QN => net108387);
   registers_reg_15_31_inst : DFFR_X1 port map( D => n3558, CK => n591, RN => 
                           rst, Q => registers_15_31_port, QN => net108386);
   registers_reg_15_30_inst : DFFR_X1 port map( D => n3557, CK => n570, RN => 
                           rst, Q => registers_15_30_port, QN => net108385);
   registers_reg_15_29_inst : DFFR_X1 port map( D => n3556, CK => n573, RN => 
                           rst, Q => registers_15_29_port, QN => net108384);
   registers_reg_15_28_inst : DFFR_X1 port map( D => n3555, CK => n576, RN => 
                           rst, Q => registers_15_28_port, QN => net108383);
   registers_reg_15_27_inst : DFFR_X1 port map( D => n3554, CK => n583, RN => 
                           rst, Q => registers_15_27_port, QN => net108382);
   registers_reg_15_26_inst : DFFR_X1 port map( D => n3553, CK => n548, RN => 
                           rst, Q => registers_15_26_port, QN => net108381);
   registers_reg_15_25_inst : DFFR_X1 port map( D => n3552, CK => n564, RN => 
                           rst, Q => registers_15_25_port, QN => net108380);
   registers_reg_15_24_inst : DFFR_X1 port map( D => n3551, CK => n586, RN => 
                           rst, Q => registers_15_24_port, QN => net108379);
   registers_reg_15_23_inst : DFFR_X1 port map( D => n3550, CK => n551, RN => 
                           rst, Q => registers_15_23_port, QN => net108378);
   registers_reg_15_22_inst : DFFR_X1 port map( D => n3549, CK => n566, RN => 
                           rst, Q => registers_15_22_port, QN => net108377);
   registers_reg_15_21_inst : DFFR_X1 port map( D => n3548, CK => n622, RN => 
                           rst, Q => registers_15_21_port, QN => net108376);
   registers_reg_15_20_inst : DFFR_X1 port map( D => n3547, CK => n554, RN => 
                           rst, Q => registers_15_20_port, QN => net108375);
   registers_reg_15_19_inst : DFFR_X1 port map( D => n3546, CK => n616, RN => 
                           rst, Q => registers_15_19_port, QN => net108374);
   registers_reg_15_18_inst : DFFR_X1 port map( D => n3545, CK => n624, RN => 
                           rst, Q => registers_15_18_port, QN => net108373);
   registers_reg_15_17_inst : DFFR_X1 port map( D => n3544, CK => n629, RN => 
                           rst, Q => registers_15_17_port, QN => net108372);
   registers_reg_15_16_inst : DFFR_X1 port map( D => n3543, CK => n632, RN => 
                           rst, Q => registers_15_16_port, QN => net108371);
   registers_reg_15_15_inst : DFFR_X1 port map( D => n3542, CK => n558, RN => 
                           rst, Q => registers_15_15_port, QN => net108370);
   registers_reg_15_14_inst : DFFR_X1 port map( D => n3541, CK => n598, RN => 
                           rst, Q => registers_15_14_port, QN => net108369);
   registers_reg_15_13_inst : DFFR_X1 port map( D => n3540, CK => n601, RN => 
                           rst, Q => registers_15_13_port, QN => net108368);
   registers_reg_15_12_inst : DFFR_X1 port map( D => n3539, CK => n626, RN => 
                           rst, Q => registers_15_12_port, QN => net108367);
   registers_reg_15_11_inst : DFFR_X1 port map( D => n3538, CK => n593, RN => 
                           rst, Q => registers_15_11_port, QN => net108366);
   registers_reg_15_10_inst : DFFR_X1 port map( D => n3537, CK => n610, RN => 
                           rst, Q => registers_15_10_port, QN => net108365);
   registers_reg_15_9_inst : DFFR_X1 port map( D => n3536, CK => n588, RN => 
                           rst, Q => registers_15_9_port, QN => net108364);
   registers_reg_15_8_inst : DFFR_X1 port map( D => n3535, CK => n561, RN => 
                           rst, Q => registers_15_8_port, QN => net108363);
   registers_reg_15_7_inst : DFFR_X1 port map( D => n3534, CK => n546, RN => 
                           rst, Q => registers_15_7_port, QN => net108362);
   registers_reg_15_6_inst : DFFR_X1 port map( D => n3533, CK => n595, RN => 
                           rst, Q => registers_15_6_port, QN => net108361);
   registers_reg_15_5_inst : DFFR_X1 port map( D => n3532, CK => n580, RN => 
                           rst, Q => registers_15_5_port, QN => net108360);
   registers_reg_15_4_inst : DFFR_X1 port map( D => n3531, CK => n619, RN => 
                           rst, Q => registers_15_4_port, QN => net108359);
   registers_reg_15_3_inst : DFFR_X1 port map( D => n3530, CK => n612, RN => 
                           rst, Q => registers_15_3_port, QN => net108358);
   registers_reg_15_2_inst : DFFR_X1 port map( D => n3529, CK => n607, RN => 
                           rst, Q => registers_15_2_port, QN => net108357);
   registers_reg_15_1_inst : DFFR_X1 port map( D => n3528, CK => n633, RN => 
                           rst, Q => registers_15_1_port, QN => net108356);
   registers_reg_15_0_inst : DFFR_X1 port map( D => n3527, CK => n579, RN => 
                           rst, Q => registers_15_0_port, QN => net108355);
   registers_reg_16_31_inst : DFFR_X1 port map( D => n3526, CK => n591, RN => 
                           rst, Q => registers_16_31_port, QN => n225);
   registers_reg_16_30_inst : DFFR_X1 port map( D => n3525, CK => n570, RN => 
                           rst, Q => registers_16_30_port, QN => n227);
   registers_reg_16_29_inst : DFFR_X1 port map( D => n3524, CK => n573, RN => 
                           rst, Q => registers_16_29_port, QN => n229);
   registers_reg_16_28_inst : DFFR_X1 port map( D => n3523, CK => n576, RN => 
                           rst, Q => registers_16_28_port, QN => n231);
   registers_reg_16_27_inst : DFFR_X1 port map( D => n3522, CK => n583, RN => 
                           rst, Q => registers_16_27_port, QN => n233);
   registers_reg_16_26_inst : DFFR_X1 port map( D => n3521, CK => n548, RN => 
                           rst, Q => registers_16_26_port, QN => n235);
   registers_reg_16_25_inst : DFFR_X1 port map( D => n3520, CK => n564, RN => 
                           rst, Q => registers_16_25_port, QN => n237);
   registers_reg_16_24_inst : DFFR_X1 port map( D => n3519, CK => n585, RN => 
                           rst, Q => registers_16_24_port, QN => n239);
   registers_reg_16_23_inst : DFFR_X1 port map( D => n3518, CK => n551, RN => 
                           rst, Q => registers_16_23_port, QN => n241);
   registers_reg_16_22_inst : DFFR_X1 port map( D => n3517, CK => n566, RN => 
                           rst, Q => registers_16_22_port, QN => n243);
   registers_reg_16_21_inst : DFFR_X1 port map( D => n3516, CK => n622, RN => 
                           rst, Q => registers_16_21_port, QN => n245);
   registers_reg_16_20_inst : DFFR_X1 port map( D => n3515, CK => n554, RN => 
                           rst, Q => registers_16_20_port, QN => n247);
   registers_reg_16_19_inst : DFFR_X1 port map( D => n3514, CK => n616, RN => 
                           rst, Q => registers_16_19_port, QN => n249);
   registers_reg_16_18_inst : DFFR_X1 port map( D => n3513, CK => n624, RN => 
                           rst, Q => registers_16_18_port, QN => n251);
   registers_reg_16_17_inst : DFFR_X1 port map( D => n3512, CK => n628, RN => 
                           rst, Q => registers_16_17_port, QN => n253);
   registers_reg_16_16_inst : DFFR_X1 port map( D => n3511, CK => n632, RN => 
                           rst, Q => registers_16_16_port, QN => n255);
   registers_reg_16_15_inst : DFFR_X1 port map( D => n3510, CK => n558, RN => 
                           rst, Q => registers_16_15_port, QN => n257);
   registers_reg_16_14_inst : DFFR_X1 port map( D => n3509, CK => n598, RN => 
                           rst, Q => registers_16_14_port, QN => n259);
   registers_reg_16_13_inst : DFFR_X1 port map( D => n3508, CK => n601, RN => 
                           rst, Q => registers_16_13_port, QN => n261);
   registers_reg_16_12_inst : DFFR_X1 port map( D => n3507, CK => n626, RN => 
                           rst, Q => registers_16_12_port, QN => n263);
   registers_reg_16_11_inst : DFFR_X1 port map( D => n3506, CK => n593, RN => 
                           rst, Q => registers_16_11_port, QN => n265);
   registers_reg_16_10_inst : DFFR_X1 port map( D => n3505, CK => n609, RN => 
                           rst, Q => registers_16_10_port, QN => n267);
   registers_reg_16_9_inst : DFFR_X1 port map( D => n3504, CK => n588, RN => 
                           rst, Q => registers_16_9_port, QN => n269);
   registers_reg_16_8_inst : DFFR_X1 port map( D => n3503, CK => n561, RN => 
                           rst, Q => registers_16_8_port, QN => n271);
   registers_reg_16_7_inst : DFFR_X1 port map( D => n3502, CK => n546, RN => 
                           rst, Q => registers_16_7_port, QN => n273);
   registers_reg_16_6_inst : DFFR_X1 port map( D => n3501, CK => n595, RN => 
                           rst, Q => registers_16_6_port, QN => n275);
   registers_reg_16_5_inst : DFFR_X1 port map( D => n3500, CK => n580, RN => 
                           rst, Q => registers_16_5_port, QN => n277);
   registers_reg_16_4_inst : DFFR_X1 port map( D => n3499, CK => n619, RN => 
                           rst, Q => registers_16_4_port, QN => n279);
   registers_reg_16_3_inst : DFFR_X1 port map( D => n3498, CK => n612, RN => 
                           rst, Q => registers_16_3_port, QN => n281);
   registers_reg_16_2_inst : DFFR_X1 port map( D => n3497, CK => n607, RN => 
                           rst, Q => registers_16_2_port, QN => n283);
   registers_reg_16_1_inst : DFFR_X1 port map( D => n3496, CK => n632, RN => 
                           rst, Q => registers_16_1_port, QN => n285);
   registers_reg_16_0_inst : DFFR_X1 port map( D => n3495, CK => n579, RN => 
                           rst, Q => registers_16_0_port, QN => n287);
   registers_reg_17_31_inst : DFFR_X1 port map( D => n3494, CK => n591, RN => 
                           rst, Q => registers_17_31_port, QN => n1);
   registers_reg_17_30_inst : DFFR_X1 port map( D => n3493, CK => n570, RN => 
                           rst, Q => registers_17_30_port, QN => n3);
   registers_reg_17_29_inst : DFFR_X1 port map( D => n3492, CK => n573, RN => 
                           rst, Q => registers_17_29_port, QN => n5);
   registers_reg_17_28_inst : DFFR_X1 port map( D => n3491, CK => n576, RN => 
                           rst, Q => registers_17_28_port, QN => n7);
   registers_reg_17_27_inst : DFFR_X1 port map( D => n3490, CK => n583, RN => 
                           rst, Q => registers_17_27_port, QN => n9);
   registers_reg_17_26_inst : DFFR_X1 port map( D => n3489, CK => n548, RN => 
                           rst, Q => registers_17_26_port, QN => n11);
   registers_reg_17_25_inst : DFFR_X1 port map( D => n3488, CK => n564, RN => 
                           rst, Q => registers_17_25_port, QN => n13);
   registers_reg_17_24_inst : DFFR_X1 port map( D => n3487, CK => n585, RN => 
                           rst, Q => registers_17_24_port, QN => n15);
   registers_reg_17_23_inst : DFFR_X1 port map( D => n3486, CK => n551, RN => 
                           rst, Q => registers_17_23_port, QN => n17);
   registers_reg_17_22_inst : DFFR_X1 port map( D => n3485, CK => n566, RN => 
                           rst, Q => registers_17_22_port, QN => n19);
   registers_reg_17_21_inst : DFFR_X1 port map( D => n3484, CK => n621, RN => 
                           rst, Q => registers_17_21_port, QN => n21);
   registers_reg_17_20_inst : DFFR_X1 port map( D => n3483, CK => n554, RN => 
                           rst, Q => registers_17_20_port, QN => n23);
   registers_reg_17_19_inst : DFFR_X1 port map( D => n3482, CK => n616, RN => 
                           rst, Q => registers_17_19_port, QN => n25);
   registers_reg_17_18_inst : DFFR_X1 port map( D => n3481, CK => n624, RN => 
                           rst, Q => registers_17_18_port, QN => n27);
   registers_reg_17_17_inst : DFFR_X1 port map( D => n3480, CK => n628, RN => 
                           rst, Q => registers_17_17_port, QN => n29);
   registers_reg_17_16_inst : DFFR_X1 port map( D => n3479, CK => n631, RN => 
                           rst, Q => registers_17_16_port, QN => n31);
   registers_reg_17_15_inst : DFFR_X1 port map( D => n3478, CK => n558, RN => 
                           rst, Q => registers_17_15_port, QN => n33);
   registers_reg_17_14_inst : DFFR_X1 port map( D => n3477, CK => n598, RN => 
                           rst, Q => registers_17_14_port, QN => n35);
   registers_reg_17_13_inst : DFFR_X1 port map( D => n3476, CK => n601, RN => 
                           rst, Q => registers_17_13_port, QN => n37);
   registers_reg_17_12_inst : DFFR_X1 port map( D => n3475, CK => n626, RN => 
                           rst, Q => registers_17_12_port, QN => n39);
   registers_reg_17_11_inst : DFFR_X1 port map( D => n3474, CK => n592, RN => 
                           rst, Q => registers_17_11_port, QN => n41);
   registers_reg_17_10_inst : DFFR_X1 port map( D => n3473, CK => n609, RN => 
                           rst, Q => registers_17_10_port, QN => n43);
   registers_reg_17_9_inst : DFFR_X1 port map( D => n3472, CK => n588, RN => 
                           rst, Q => registers_17_9_port, QN => n45);
   registers_reg_17_8_inst : DFFR_X1 port map( D => n3471, CK => n561, RN => 
                           rst, Q => registers_17_8_port, QN => n47);
   registers_reg_17_7_inst : DFFR_X1 port map( D => n3470, CK => n545, RN => 
                           rst, Q => registers_17_7_port, QN => n49);
   registers_reg_17_6_inst : DFFR_X1 port map( D => n3469, CK => n595, RN => 
                           rst, Q => registers_17_6_port, QN => n51);
   registers_reg_17_5_inst : DFFR_X1 port map( D => n3468, CK => n580, RN => 
                           rst, Q => registers_17_5_port, QN => n53);
   registers_reg_17_4_inst : DFFR_X1 port map( D => n3467, CK => n619, RN => 
                           rst, Q => registers_17_4_port, QN => n55);
   registers_reg_17_3_inst : DFFR_X1 port map( D => n3466, CK => n612, RN => 
                           rst, Q => registers_17_3_port, QN => n57);
   registers_reg_17_2_inst : DFFR_X1 port map( D => n3465, CK => n607, RN => 
                           rst, Q => registers_17_2_port, QN => n59);
   registers_reg_17_1_inst : DFFR_X1 port map( D => n3464, CK => n634, RN => 
                           rst, Q => registers_17_1_port, QN => n61);
   registers_reg_17_0_inst : DFFR_X1 port map( D => n3463, CK => n579, RN => 
                           rst, Q => registers_17_0_port, QN => n63);
   registers_reg_18_31_inst : DFFR_X1 port map( D => n3462, CK => n591, RN => 
                           rst, Q => registers_18_31_port, QN => n159);
   registers_reg_18_30_inst : DFFR_X1 port map( D => n3461, CK => n570, RN => 
                           rst, Q => registers_18_30_port, QN => n97);
   registers_reg_18_29_inst : DFFR_X1 port map( D => n3460, CK => n573, RN => 
                           rst, Q => registers_18_29_port, QN => n99);
   registers_reg_18_28_inst : DFFR_X1 port map( D => n3459, CK => n576, RN => 
                           rst, Q => registers_18_28_port, QN => n101);
   registers_reg_18_27_inst : DFFR_X1 port map( D => n3458, CK => n583, RN => 
                           rst, Q => registers_18_27_port, QN => n103);
   registers_reg_18_26_inst : DFFR_X1 port map( D => n3457, CK => n548, RN => 
                           rst, Q => registers_18_26_port, QN => n105);
   registers_reg_18_25_inst : DFFR_X1 port map( D => n3456, CK => n563, RN => 
                           rst, Q => registers_18_25_port, QN => n107);
   registers_reg_18_24_inst : DFFR_X1 port map( D => n3455, CK => n585, RN => 
                           rst, Q => registers_18_24_port, QN => n109);
   registers_reg_18_23_inst : DFFR_X1 port map( D => n3454, CK => n551, RN => 
                           rst, Q => registers_18_23_port, QN => n111);
   registers_reg_18_22_inst : DFFR_X1 port map( D => n3453, CK => n566, RN => 
                           rst, Q => registers_18_22_port, QN => n113);
   registers_reg_18_21_inst : DFFR_X1 port map( D => n3452, CK => n621, RN => 
                           rst, Q => registers_18_21_port, QN => n115);
   registers_reg_18_20_inst : DFFR_X1 port map( D => n3451, CK => n554, RN => 
                           rst, Q => registers_18_20_port, QN => n117);
   registers_reg_18_19_inst : DFFR_X1 port map( D => n3450, CK => n616, RN => 
                           rst, Q => registers_18_19_port, QN => n119);
   registers_reg_18_18_inst : DFFR_X1 port map( D => n3449, CK => n624, RN => 
                           rst, Q => registers_18_18_port, QN => n121);
   registers_reg_18_17_inst : DFFR_X1 port map( D => n3448, CK => n628, RN => 
                           rst, Q => registers_18_17_port, QN => n123);
   registers_reg_18_16_inst : DFFR_X1 port map( D => n3447, CK => n631, RN => 
                           rst, Q => registers_18_16_port, QN => n125);
   registers_reg_18_15_inst : DFFR_X1 port map( D => n3446, CK => n558, RN => 
                           rst, Q => registers_18_15_port, QN => n127);
   registers_reg_18_14_inst : DFFR_X1 port map( D => n3445, CK => n598, RN => 
                           rst, Q => registers_18_14_port, QN => n129);
   registers_reg_18_13_inst : DFFR_X1 port map( D => n3444, CK => n601, RN => 
                           rst, Q => registers_18_13_port, QN => n131);
   registers_reg_18_12_inst : DFFR_X1 port map( D => n3443, CK => n626, RN => 
                           rst, Q => registers_18_12_port, QN => n133);
   registers_reg_18_11_inst : DFFR_X1 port map( D => n3442, CK => n592, RN => 
                           rst, Q => registers_18_11_port, QN => n135);
   registers_reg_18_10_inst : DFFR_X1 port map( D => n3441, CK => n609, RN => 
                           rst, Q => registers_18_10_port, QN => n137);
   registers_reg_18_9_inst : DFFR_X1 port map( D => n3440, CK => n588, RN => 
                           rst, Q => registers_18_9_port, QN => n139);
   registers_reg_18_8_inst : DFFR_X1 port map( D => n3439, CK => n561, RN => 
                           rst, Q => registers_18_8_port, QN => n141);
   registers_reg_18_7_inst : DFFR_X1 port map( D => n3438, CK => n545, RN => 
                           rst, Q => registers_18_7_port, QN => n143);
   registers_reg_18_6_inst : DFFR_X1 port map( D => n3437, CK => n595, RN => 
                           rst, Q => registers_18_6_port, QN => n145);
   registers_reg_18_5_inst : DFFR_X1 port map( D => n3436, CK => n586, RN => 
                           rst, Q => registers_18_5_port, QN => n147);
   registers_reg_18_4_inst : DFFR_X1 port map( D => n3435, CK => n619, RN => 
                           rst, Q => registers_18_4_port, QN => n149);
   registers_reg_18_3_inst : DFFR_X1 port map( D => n3434, CK => n612, RN => 
                           rst, Q => registers_18_3_port, QN => n151);
   registers_reg_18_2_inst : DFFR_X1 port map( D => n3433, CK => n606, RN => 
                           rst, Q => registers_18_2_port, QN => n153);
   registers_reg_18_1_inst : DFFR_X1 port map( D => n3432, CK => n633, RN => 
                           rst, Q => registers_18_1_port, QN => n155);
   registers_reg_18_0_inst : DFFR_X1 port map( D => n3431, CK => n578, RN => 
                           rst, Q => registers_18_0_port, QN => n157);
   registers_reg_19_31_inst : DFFR_X1 port map( D => n3430, CK => n591, RN => 
                           rst, Q => registers_19_31_port, QN => net108354);
   registers_reg_19_30_inst : DFFR_X1 port map( D => n3429, CK => n570, RN => 
                           rst, Q => registers_19_30_port, QN => net108353);
   registers_reg_19_29_inst : DFFR_X1 port map( D => n3428, CK => n573, RN => 
                           rst, Q => registers_19_29_port, QN => net108352);
   registers_reg_19_28_inst : DFFR_X1 port map( D => n3427, CK => n575, RN => 
                           rst, Q => registers_19_28_port, QN => net108351);
   registers_reg_19_27_inst : DFFR_X1 port map( D => n3426, CK => n582, RN => 
                           rst, Q => registers_19_27_port, QN => net108350);
   registers_reg_19_26_inst : DFFR_X1 port map( D => n3425, CK => n548, RN => 
                           rst, Q => registers_19_26_port, QN => net108349);
   registers_reg_19_25_inst : DFFR_X1 port map( D => n3424, CK => n563, RN => 
                           rst, Q => registers_19_25_port, QN => net108348);
   registers_reg_19_24_inst : DFFR_X1 port map( D => n3423, CK => n585, RN => 
                           rst, Q => registers_19_24_port, QN => net108347);
   registers_reg_19_23_inst : DFFR_X1 port map( D => n3422, CK => n551, RN => 
                           rst, Q => registers_19_23_port, QN => net108346);
   registers_reg_19_22_inst : DFFR_X1 port map( D => n3421, CK => n566, RN => 
                           rst, Q => registers_19_22_port, QN => net108345);
   registers_reg_19_21_inst : DFFR_X1 port map( D => n3420, CK => n621, RN => 
                           rst, Q => registers_19_21_port, QN => net108344);
   registers_reg_19_20_inst : DFFR_X1 port map( D => n3419, CK => n554, RN => 
                           rst, Q => registers_19_20_port, QN => net108343);
   registers_reg_19_19_inst : DFFR_X1 port map( D => n3418, CK => n616, RN => 
                           rst, Q => registers_19_19_port, QN => net108342);
   registers_reg_19_18_inst : DFFR_X1 port map( D => n3417, CK => n624, RN => 
                           rst, Q => registers_19_18_port, QN => net108341);
   registers_reg_19_17_inst : DFFR_X1 port map( D => n3416, CK => n628, RN => 
                           rst, Q => registers_19_17_port, QN => net108340);
   registers_reg_19_16_inst : DFFR_X1 port map( D => n3415, CK => n631, RN => 
                           rst, Q => registers_19_16_port, QN => net108339);
   registers_reg_19_15_inst : DFFR_X1 port map( D => n3414, CK => n558, RN => 
                           rst, Q => registers_19_15_port, QN => net108338);
   registers_reg_19_14_inst : DFFR_X1 port map( D => n3413, CK => n598, RN => 
                           rst, Q => registers_19_14_port, QN => net108337);
   registers_reg_19_13_inst : DFFR_X1 port map( D => n3412, CK => n601, RN => 
                           rst, Q => registers_19_13_port, QN => net108336);
   registers_reg_19_12_inst : DFFR_X1 port map( D => n3411, CK => n625, RN => 
                           rst, Q => registers_19_12_port, QN => net108335);
   registers_reg_19_11_inst : DFFR_X1 port map( D => n3410, CK => n592, RN => 
                           rst, Q => registers_19_11_port, QN => net108334);
   registers_reg_19_10_inst : DFFR_X1 port map( D => n3409, CK => n609, RN => 
                           rst, Q => registers_19_10_port, QN => net108333);
   registers_reg_19_9_inst : DFFR_X1 port map( D => n3408, CK => n588, RN => 
                           rst, Q => registers_19_9_port, QN => net108332);
   registers_reg_19_8_inst : DFFR_X1 port map( D => n3407, CK => n561, RN => 
                           rst, Q => registers_19_8_port, QN => net108331);
   registers_reg_19_7_inst : DFFR_X1 port map( D => n3406, CK => n545, RN => 
                           rst, Q => registers_19_7_port, QN => net108330);
   registers_reg_19_6_inst : DFFR_X1 port map( D => n3405, CK => n595, RN => 
                           rst, Q => registers_19_6_port, QN => net108329);
   registers_reg_19_5_inst : DFFR_X1 port map( D => n3404, CK => n556, RN => 
                           rst, Q => registers_19_5_port, QN => net108328);
   registers_reg_19_4_inst : DFFR_X1 port map( D => n3403, CK => n618, RN => 
                           rst, Q => registers_19_4_port, QN => net108327);
   registers_reg_19_3_inst : DFFR_X1 port map( D => n3402, CK => n612, RN => 
                           rst, Q => registers_19_3_port, QN => net108326);
   registers_reg_19_2_inst : DFFR_X1 port map( D => n3401, CK => n606, RN => 
                           rst, Q => registers_19_2_port, QN => net108325);
   registers_reg_19_1_inst : DFFR_X1 port map( D => n3400, CK => n635, RN => 
                           rst, Q => registers_19_1_port, QN => net108324);
   registers_reg_19_0_inst : DFFR_X1 port map( D => n3399, CK => n578, RN => 
                           rst, Q => registers_19_0_port, QN => net108323);
   registers_reg_20_31_inst : DFFR_X1 port map( D => n3398, CK => n591, RN => 
                           rst, Q => registers_20_31_port, QN => net108322);
   registers_reg_20_30_inst : DFFR_X1 port map( D => n3397, CK => n570, RN => 
                           rst, Q => registers_20_30_port, QN => net108321);
   registers_reg_20_29_inst : DFFR_X1 port map( D => n3396, CK => n573, RN => 
                           rst, Q => registers_20_29_port, QN => net108320);
   registers_reg_20_28_inst : DFFR_X1 port map( D => n3395, CK => n575, RN => 
                           rst, Q => registers_20_28_port, QN => net108319);
   registers_reg_20_27_inst : DFFR_X1 port map( D => n3394, CK => n582, RN => 
                           rst, Q => registers_20_27_port, QN => net108318);
   registers_reg_20_26_inst : DFFR_X1 port map( D => n3393, CK => n548, RN => 
                           rst, Q => registers_20_26_port, QN => net108317);
   registers_reg_20_25_inst : DFFR_X1 port map( D => n3392, CK => n563, RN => 
                           rst, Q => registers_20_25_port, QN => net108316);
   registers_reg_20_24_inst : DFFR_X1 port map( D => n3391, CK => n585, RN => 
                           rst, Q => registers_20_24_port, QN => net108315);
   registers_reg_20_23_inst : DFFR_X1 port map( D => n3390, CK => n551, RN => 
                           rst, Q => registers_20_23_port, QN => net108314);
   registers_reg_20_22_inst : DFFR_X1 port map( D => n3389, CK => n566, RN => 
                           rst, Q => registers_20_22_port, QN => net108313);
   registers_reg_20_21_inst : DFFR_X1 port map( D => n3388, CK => n621, RN => 
                           rst, Q => registers_20_21_port, QN => net108312);
   registers_reg_20_20_inst : DFFR_X1 port map( D => n3387, CK => n553, RN => 
                           rst, Q => registers_20_20_port, QN => net108311);
   registers_reg_20_19_inst : DFFR_X1 port map( D => n3386, CK => n616, RN => 
                           rst, Q => registers_20_19_port, QN => net108310);
   registers_reg_20_18_inst : DFFR_X1 port map( D => n3385, CK => n624, RN => 
                           rst, Q => registers_20_18_port, QN => net108309);
   registers_reg_20_17_inst : DFFR_X1 port map( D => n3384, CK => n628, RN => 
                           rst, Q => registers_20_17_port, QN => net108308);
   registers_reg_20_16_inst : DFFR_X1 port map( D => n3383, CK => n631, RN => 
                           rst, Q => registers_20_16_port, QN => net108307);
   registers_reg_20_15_inst : DFFR_X1 port map( D => n3382, CK => n558, RN => 
                           rst, Q => registers_20_15_port, QN => net108306);
   registers_reg_20_14_inst : DFFR_X1 port map( D => n3381, CK => n598, RN => 
                           rst, Q => registers_20_14_port, QN => net108305);
   registers_reg_20_13_inst : DFFR_X1 port map( D => n3380, CK => n600, RN => 
                           rst, Q => registers_20_13_port, QN => net108304);
   registers_reg_20_12_inst : DFFR_X1 port map( D => n3379, CK => n625, RN => 
                           rst, Q => registers_20_12_port, QN => net108303);
   registers_reg_20_11_inst : DFFR_X1 port map( D => n3378, CK => n592, RN => 
                           rst, Q => registers_20_11_port, QN => net108302);
   registers_reg_20_10_inst : DFFR_X1 port map( D => n3377, CK => n609, RN => 
                           rst, Q => registers_20_10_port, QN => net108301);
   registers_reg_20_9_inst : DFFR_X1 port map( D => n3376, CK => n588, RN => 
                           rst, Q => registers_20_9_port, QN => net108300);
   registers_reg_20_8_inst : DFFR_X1 port map( D => n3375, CK => n560, RN => 
                           rst, Q => registers_20_8_port, QN => net108299);
   registers_reg_20_7_inst : DFFR_X1 port map( D => n3374, CK => n545, RN => 
                           rst, Q => registers_20_7_port, QN => net108298);
   registers_reg_20_6_inst : DFFR_X1 port map( D => n3373, CK => n595, RN => 
                           rst, Q => registers_20_6_port, QN => net108297);
   registers_reg_20_5_inst : DFFR_X1 port map( D => n3372, CK => n556, RN => 
                           rst, Q => registers_20_5_port, QN => net108296);
   registers_reg_20_4_inst : DFFR_X1 port map( D => n3371, CK => n618, RN => 
                           rst, Q => registers_20_4_port, QN => net108295);
   registers_reg_20_3_inst : DFFR_X1 port map( D => n3370, CK => n612, RN => 
                           rst, Q => registers_20_3_port, QN => net108294);
   registers_reg_20_2_inst : DFFR_X1 port map( D => n3369, CK => n606, RN => 
                           rst, Q => registers_20_2_port, QN => net108293);
   registers_reg_20_1_inst : DFFR_X1 port map( D => n3368, CK => n635, RN => 
                           rst, Q => registers_20_1_port, QN => net108292);
   registers_reg_20_0_inst : DFFR_X1 port map( D => n3367, CK => n578, RN => 
                           rst, Q => registers_20_0_port, QN => net108291);
   registers_reg_21_31_inst : DFFR_X1 port map( D => n3366, CK => n591, RN => 
                           rst, Q => registers_21_31_port, QN => n226);
   registers_reg_21_30_inst : DFFR_X1 port map( D => n3365, CK => n570, RN => 
                           rst, Q => registers_21_30_port, QN => n228);
   registers_reg_21_29_inst : DFFR_X1 port map( D => n3364, CK => n572, RN => 
                           rst, Q => registers_21_29_port, QN => n230);
   registers_reg_21_28_inst : DFFR_X1 port map( D => n3363, CK => n575, RN => 
                           rst, Q => registers_21_28_port, QN => n232);
   registers_reg_21_27_inst : DFFR_X1 port map( D => n3362, CK => n582, RN => 
                           rst, Q => registers_21_27_port, QN => n234);
   registers_reg_21_26_inst : DFFR_X1 port map( D => n3361, CK => n548, RN => 
                           rst, Q => registers_21_26_port, QN => n236);
   registers_reg_21_25_inst : DFFR_X1 port map( D => n3360, CK => n563, RN => 
                           rst, Q => registers_21_25_port, QN => n238);
   registers_reg_21_24_inst : DFFR_X1 port map( D => n3359, CK => n585, RN => 
                           rst, Q => registers_21_24_port, QN => n240);
   registers_reg_21_23_inst : DFFR_X1 port map( D => n3358, CK => n551, RN => 
                           rst, Q => registers_21_23_port, QN => n242);
   registers_reg_21_22_inst : DFFR_X1 port map( D => n3357, CK => n566, RN => 
                           rst, Q => registers_21_22_port, QN => n244);
   registers_reg_21_21_inst : DFFR_X1 port map( D => n3356, CK => n621, RN => 
                           rst, Q => registers_21_21_port, QN => n246);
   registers_reg_21_20_inst : DFFR_X1 port map( D => n3355, CK => n553, RN => 
                           rst, Q => registers_21_20_port, QN => n248);
   registers_reg_21_19_inst : DFFR_X1 port map( D => n3354, CK => n616, RN => 
                           rst, Q => registers_21_19_port, QN => n250);
   registers_reg_21_18_inst : DFFR_X1 port map( D => n3353, CK => n624, RN => 
                           rst, Q => registers_21_18_port, QN => n252);
   registers_reg_21_17_inst : DFFR_X1 port map( D => n3352, CK => n628, RN => 
                           rst, Q => registers_21_17_port, QN => n254);
   registers_reg_21_16_inst : DFFR_X1 port map( D => n3351, CK => n631, RN => 
                           rst, Q => registers_21_16_port, QN => n256);
   registers_reg_21_15_inst : DFFR_X1 port map( D => n3350, CK => n558, RN => 
                           rst, Q => registers_21_15_port, QN => n258);
   registers_reg_21_14_inst : DFFR_X1 port map( D => n3349, CK => n598, RN => 
                           rst, Q => registers_21_14_port, QN => n260);
   registers_reg_21_13_inst : DFFR_X1 port map( D => n3348, CK => n600, RN => 
                           rst, Q => registers_21_13_port, QN => n262);
   registers_reg_21_12_inst : DFFR_X1 port map( D => n3347, CK => n625, RN => 
                           rst, Q => registers_21_12_port, QN => n264);
   registers_reg_21_11_inst : DFFR_X1 port map( D => n3346, CK => n592, RN => 
                           rst, Q => registers_21_11_port, QN => n266);
   registers_reg_21_10_inst : DFFR_X1 port map( D => n3345, CK => n609, RN => 
                           rst, Q => registers_21_10_port, QN => n268);
   registers_reg_21_9_inst : DFFR_X1 port map( D => n3344, CK => n588, RN => 
                           rst, Q => registers_21_9_port, QN => n270);
   registers_reg_21_8_inst : DFFR_X1 port map( D => n3343, CK => n560, RN => 
                           rst, Q => registers_21_8_port, QN => n272);
   registers_reg_21_7_inst : DFFR_X1 port map( D => n3342, CK => n545, RN => 
                           rst, Q => registers_21_7_port, QN => n274);
   registers_reg_21_6_inst : DFFR_X1 port map( D => n3341, CK => n595, RN => 
                           rst, Q => registers_21_6_port, QN => n276);
   registers_reg_21_5_inst : DFFR_X1 port map( D => n3340, CK => n556, RN => 
                           rst, Q => registers_21_5_port, QN => n278);
   registers_reg_21_4_inst : DFFR_X1 port map( D => n3339, CK => n618, RN => 
                           rst, Q => registers_21_4_port, QN => n280);
   registers_reg_21_3_inst : DFFR_X1 port map( D => n3338, CK => n612, RN => 
                           rst, Q => registers_21_3_port, QN => n282);
   registers_reg_21_2_inst : DFFR_X1 port map( D => n3337, CK => n606, RN => 
                           rst, Q => registers_21_2_port, QN => n284);
   registers_reg_21_1_inst : DFFR_X1 port map( D => n3336, CK => n633, RN => 
                           rst, Q => registers_21_1_port, QN => n286);
   registers_reg_21_0_inst : DFFR_X1 port map( D => n3335, CK => n578, RN => 
                           rst, Q => registers_21_0_port, QN => n288);
   registers_reg_22_31_inst : DFFR_X1 port map( D => n3334, CK => n590, RN => 
                           rst, Q => registers_22_31_port, QN => net108290);
   registers_reg_22_30_inst : DFFR_X1 port map( D => n3333, CK => n570, RN => 
                           rst, Q => registers_22_30_port, QN => net108289);
   registers_reg_22_29_inst : DFFR_X1 port map( D => n3332, CK => n572, RN => 
                           rst, Q => registers_22_29_port, QN => net108288);
   registers_reg_22_28_inst : DFFR_X1 port map( D => n3331, CK => n575, RN => 
                           rst, Q => registers_22_28_port, QN => net108287);
   registers_reg_22_27_inst : DFFR_X1 port map( D => n3330, CK => n582, RN => 
                           rst, Q => registers_22_27_port, QN => net108286);
   registers_reg_22_26_inst : DFFR_X1 port map( D => n3329, CK => n548, RN => 
                           rst, Q => registers_22_26_port, QN => net108285);
   registers_reg_22_25_inst : DFFR_X1 port map( D => n3328, CK => n563, RN => 
                           rst, Q => registers_22_25_port, QN => net108284);
   registers_reg_22_24_inst : DFFR_X1 port map( D => n3327, CK => n585, RN => 
                           rst, Q => registers_22_24_port, QN => net108283);
   registers_reg_22_23_inst : DFFR_X1 port map( D => n3326, CK => n551, RN => 
                           rst, Q => registers_22_23_port, QN => net108282);
   registers_reg_22_22_inst : DFFR_X1 port map( D => n3325, CK => n566, RN => 
                           rst, Q => registers_22_22_port, QN => net108281);
   registers_reg_22_21_inst : DFFR_X1 port map( D => n3324, CK => n621, RN => 
                           rst, Q => registers_22_21_port, QN => net108280);
   registers_reg_22_20_inst : DFFR_X1 port map( D => n3323, CK => n553, RN => 
                           rst, Q => registers_22_20_port, QN => net108279);
   registers_reg_22_19_inst : DFFR_X1 port map( D => n3322, CK => n615, RN => 
                           rst, Q => registers_22_19_port, QN => net108278);
   registers_reg_22_18_inst : DFFR_X1 port map( D => n3321, CK => n624, RN => 
                           rst, Q => registers_22_18_port, QN => net108277);
   registers_reg_22_17_inst : DFFR_X1 port map( D => n3320, CK => n628, RN => 
                           rst, Q => registers_22_17_port, QN => net108276);
   registers_reg_22_16_inst : DFFR_X1 port map( D => n3319, CK => n631, RN => 
                           rst, Q => registers_22_16_port, QN => net108275);
   registers_reg_22_15_inst : DFFR_X1 port map( D => n3318, CK => n558, RN => 
                           rst, Q => registers_22_15_port, QN => net108274);
   registers_reg_22_14_inst : DFFR_X1 port map( D => n3317, CK => n598, RN => 
                           rst, Q => registers_22_14_port, QN => net108273);
   registers_reg_22_13_inst : DFFR_X1 port map( D => n3316, CK => n600, RN => 
                           rst, Q => registers_22_13_port, QN => net108272);
   registers_reg_22_12_inst : DFFR_X1 port map( D => n3315, CK => n625, RN => 
                           rst, Q => registers_22_12_port, QN => net108271);
   registers_reg_22_11_inst : DFFR_X1 port map( D => n3314, CK => n592, RN => 
                           rst, Q => registers_22_11_port, QN => net108270);
   registers_reg_22_10_inst : DFFR_X1 port map( D => n3313, CK => n609, RN => 
                           rst, Q => registers_22_10_port, QN => net108269);
   registers_reg_22_9_inst : DFFR_X1 port map( D => n3312, CK => n588, RN => 
                           rst, Q => registers_22_9_port, QN => net108268);
   registers_reg_22_8_inst : DFFR_X1 port map( D => n3311, CK => n560, RN => 
                           rst, Q => registers_22_8_port, QN => net108267);
   registers_reg_22_7_inst : DFFR_X1 port map( D => n3310, CK => n545, RN => 
                           rst, Q => registers_22_7_port, QN => net108266);
   registers_reg_22_6_inst : DFFR_X1 port map( D => n3309, CK => n595, RN => 
                           rst, Q => registers_22_6_port, QN => net108265);
   registers_reg_22_5_inst : DFFR_X1 port map( D => n3308, CK => n556, RN => 
                           rst, Q => registers_22_5_port, QN => net108264);
   registers_reg_22_4_inst : DFFR_X1 port map( D => n3307, CK => n618, RN => 
                           rst, Q => registers_22_4_port, QN => net108263);
   registers_reg_22_3_inst : DFFR_X1 port map( D => n3306, CK => n612, RN => 
                           rst, Q => registers_22_3_port, QN => net108262);
   registers_reg_22_2_inst : DFFR_X1 port map( D => n3305, CK => n606, RN => 
                           rst, Q => registers_22_2_port, QN => net108261);
   registers_reg_22_1_inst : DFFR_X1 port map( D => n3304, CK => n634, RN => 
                           rst, Q => registers_22_1_port, QN => net108260);
   registers_reg_22_0_inst : DFFR_X1 port map( D => n3303, CK => n578, RN => 
                           rst, Q => registers_22_0_port, QN => net108259);
   registers_reg_23_31_inst : DFFR_X1 port map( D => n3302, CK => n590, RN => 
                           rst, Q => registers_23_31_port, QN => n542);
   registers_reg_23_30_inst : DFFR_X1 port map( D => n3301, CK => n570, RN => 
                           rst, Q => registers_23_30_port, QN => n479);
   registers_reg_23_29_inst : DFFR_X1 port map( D => n3300, CK => n572, RN => 
                           rst, Q => registers_23_29_port, QN => n481);
   registers_reg_23_28_inst : DFFR_X1 port map( D => n3299, CK => n575, RN => 
                           rst, Q => registers_23_28_port, QN => n483);
   registers_reg_23_27_inst : DFFR_X1 port map( D => n3298, CK => n582, RN => 
                           rst, Q => registers_23_27_port, QN => n485);
   registers_reg_23_26_inst : DFFR_X1 port map( D => n3297, CK => n548, RN => 
                           rst, Q => registers_23_26_port, QN => n487);
   registers_reg_23_25_inst : DFFR_X1 port map( D => n3296, CK => n563, RN => 
                           rst, Q => registers_23_25_port, QN => n489);
   registers_reg_23_24_inst : DFFR_X1 port map( D => n3295, CK => n585, RN => 
                           rst, Q => registers_23_24_port, QN => n491);
   registers_reg_23_23_inst : DFFR_X1 port map( D => n3294, CK => n550, RN => 
                           rst, Q => registers_23_23_port, QN => n493);
   registers_reg_23_22_inst : DFFR_X1 port map( D => n3293, CK => n566, RN => 
                           rst, Q => registers_23_22_port, QN => n495);
   registers_reg_23_21_inst : DFFR_X1 port map( D => n3292, CK => n621, RN => 
                           rst, Q => registers_23_21_port, QN => n497);
   registers_reg_23_20_inst : DFFR_X1 port map( D => n3291, CK => n553, RN => 
                           rst, Q => registers_23_20_port, QN => n499);
   registers_reg_23_19_inst : DFFR_X1 port map( D => n3290, CK => n615, RN => 
                           rst, Q => registers_23_19_port, QN => n501);
   registers_reg_23_18_inst : DFFR_X1 port map( D => n3289, CK => n624, RN => 
                           rst, Q => registers_23_18_port, QN => n503);
   registers_reg_23_17_inst : DFFR_X1 port map( D => n3288, CK => n628, RN => 
                           rst, Q => registers_23_17_port, QN => n505);
   registers_reg_23_16_inst : DFFR_X1 port map( D => n3287, CK => n631, RN => 
                           rst, Q => registers_23_16_port, QN => n507);
   registers_reg_23_15_inst : DFFR_X1 port map( D => n3286, CK => n557, RN => 
                           rst, Q => registers_23_15_port, QN => n509);
   registers_reg_23_14_inst : DFFR_X1 port map( D => n3285, CK => n597, RN => 
                           rst, Q => registers_23_14_port, QN => n511);
   registers_reg_23_13_inst : DFFR_X1 port map( D => n3284, CK => n600, RN => 
                           rst, Q => registers_23_13_port, QN => n513);
   registers_reg_23_12_inst : DFFR_X1 port map( D => n3283, CK => n625, RN => 
                           rst, Q => registers_23_12_port, QN => n515);
   registers_reg_23_11_inst : DFFR_X1 port map( D => n3282, CK => n592, RN => 
                           rst, Q => registers_23_11_port, QN => n517);
   registers_reg_23_10_inst : DFFR_X1 port map( D => n3281, CK => n609, RN => 
                           rst, Q => registers_23_10_port, QN => n519);
   registers_reg_23_9_inst : DFFR_X1 port map( D => n3280, CK => n588, RN => 
                           rst, Q => registers_23_9_port, QN => n521);
   registers_reg_23_8_inst : DFFR_X1 port map( D => n3279, CK => n560, RN => 
                           rst, Q => registers_23_8_port, QN => n523);
   registers_reg_23_7_inst : DFFR_X1 port map( D => n3278, CK => n545, RN => 
                           rst, Q => registers_23_7_port, QN => n525);
   registers_reg_23_6_inst : DFFR_X1 port map( D => n3277, CK => n595, RN => 
                           rst, Q => registers_23_6_port, QN => n527);
   registers_reg_23_5_inst : DFFR_X1 port map( D => n3276, CK => n556, RN => 
                           rst, Q => registers_23_5_port, QN => n529);
   registers_reg_23_4_inst : DFFR_X1 port map( D => n3275, CK => n618, RN => 
                           rst, Q => registers_23_4_port, QN => n531);
   registers_reg_23_3_inst : DFFR_X1 port map( D => n3274, CK => n614, RN => 
                           rst, Q => registers_23_3_port, QN => n533);
   registers_reg_23_2_inst : DFFR_X1 port map( D => n3273, CK => n606, RN => 
                           rst, Q => registers_23_2_port, QN => n535);
   registers_reg_23_1_inst : DFFR_X1 port map( D => n3272, CK => n634, RN => 
                           rst, Q => registers_23_1_port, QN => n537);
   registers_reg_23_0_inst : DFFR_X1 port map( D => n3271, CK => n578, RN => 
                           rst, Q => registers_23_0_port, QN => n539);
   registers_reg_24_31_inst : DFFR_X1 port map( D => n3270, CK => n590, RN => 
                           rst, Q => registers_24_31_port, QN => n160);
   registers_reg_24_30_inst : DFFR_X1 port map( D => n3269, CK => n569, RN => 
                           rst, Q => registers_24_30_port, QN => n163);
   registers_reg_24_29_inst : DFFR_X1 port map( D => n3268, CK => n572, RN => 
                           rst, Q => registers_24_29_port, QN => n165);
   registers_reg_24_28_inst : DFFR_X1 port map( D => n3267, CK => n575, RN => 
                           rst, Q => registers_24_28_port, QN => n167);
   registers_reg_24_27_inst : DFFR_X1 port map( D => n3266, CK => n582, RN => 
                           rst, Q => registers_24_27_port, QN => n169);
   registers_reg_24_26_inst : DFFR_X1 port map( D => n3265, CK => n548, RN => 
                           rst, Q => registers_24_26_port, QN => n171);
   registers_reg_24_25_inst : DFFR_X1 port map( D => n3264, CK => n563, RN => 
                           rst, Q => registers_24_25_port, QN => n173);
   registers_reg_24_24_inst : DFFR_X1 port map( D => n3263, CK => n585, RN => 
                           rst, Q => registers_24_24_port, QN => n175);
   registers_reg_24_23_inst : DFFR_X1 port map( D => n3262, CK => n550, RN => 
                           rst, Q => registers_24_23_port, QN => n177);
   registers_reg_24_22_inst : DFFR_X1 port map( D => n3261, CK => n566, RN => 
                           rst, Q => registers_24_22_port, QN => n179);
   registers_reg_24_21_inst : DFFR_X1 port map( D => n3260, CK => n621, RN => 
                           rst, Q => registers_24_21_port, QN => n181);
   registers_reg_24_20_inst : DFFR_X1 port map( D => n3259, CK => n553, RN => 
                           rst, Q => registers_24_20_port, QN => n183);
   registers_reg_24_19_inst : DFFR_X1 port map( D => n3258, CK => n615, RN => 
                           rst, Q => registers_24_19_port, QN => n185);
   registers_reg_24_18_inst : DFFR_X1 port map( D => n3257, CK => n624, RN => 
                           rst, Q => registers_24_18_port, QN => n187);
   registers_reg_24_17_inst : DFFR_X1 port map( D => n3256, CK => n628, RN => 
                           rst, Q => registers_24_17_port, QN => n189);
   registers_reg_24_16_inst : DFFR_X1 port map( D => n3255, CK => n630, RN => 
                           rst, Q => registers_24_16_port, QN => n191);
   registers_reg_24_15_inst : DFFR_X1 port map( D => n3254, CK => n557, RN => 
                           rst, Q => registers_24_15_port, QN => n193);
   registers_reg_24_14_inst : DFFR_X1 port map( D => n3253, CK => n597, RN => 
                           rst, Q => registers_24_14_port, QN => n195);
   registers_reg_24_13_inst : DFFR_X1 port map( D => n3252, CK => n600, RN => 
                           rst, Q => registers_24_13_port, QN => n197);
   registers_reg_24_12_inst : DFFR_X1 port map( D => n3251, CK => n631, RN => 
                           rst, Q => registers_24_12_port, QN => n199);
   registers_reg_24_11_inst : DFFR_X1 port map( D => n3250, CK => n592, RN => 
                           rst, Q => registers_24_11_port, QN => n201);
   registers_reg_24_10_inst : DFFR_X1 port map( D => n3249, CK => n609, RN => 
                           rst, Q => registers_24_10_port, QN => n203);
   registers_reg_24_9_inst : DFFR_X1 port map( D => n3248, CK => n588, RN => 
                           rst, Q => registers_24_9_port, QN => n205);
   registers_reg_24_8_inst : DFFR_X1 port map( D => n3247, CK => n560, RN => 
                           rst, Q => registers_24_8_port, QN => n207);
   registers_reg_24_7_inst : DFFR_X1 port map( D => n3246, CK => n545, RN => 
                           rst, Q => registers_24_7_port, QN => n209);
   registers_reg_24_6_inst : DFFR_X1 port map( D => n3245, CK => n595, RN => 
                           rst, Q => registers_24_6_port, QN => n211);
   registers_reg_24_5_inst : DFFR_X1 port map( D => n3244, CK => n556, RN => 
                           rst, Q => registers_24_5_port, QN => n213);
   registers_reg_24_4_inst : DFFR_X1 port map( D => n3243, CK => n618, RN => 
                           rst, Q => registers_24_4_port, QN => n215);
   registers_reg_24_3_inst : DFFR_X1 port map( D => n3242, CK => n611, RN => 
                           rst, Q => registers_24_3_port, QN => n217);
   registers_reg_24_2_inst : DFFR_X1 port map( D => n3241, CK => n606, RN => 
                           rst, Q => registers_24_2_port, QN => n219);
   registers_reg_24_1_inst : DFFR_X1 port map( D => n3240, CK => n634, RN => 
                           rst, Q => registers_24_1_port, QN => n221);
   registers_reg_24_0_inst : DFFR_X1 port map( D => n3239, CK => n578, RN => 
                           rst, Q => registers_24_0_port, QN => n223);
   registers_reg_25_31_inst : DFFR_X1 port map( D => n3238, CK => n590, RN => 
                           rst, Q => registers_25_31_port, QN => net108258);
   registers_reg_25_30_inst : DFFR_X1 port map( D => n3237, CK => n569, RN => 
                           rst, Q => registers_25_30_port, QN => net108257);
   registers_reg_25_29_inst : DFFR_X1 port map( D => n3236, CK => n572, RN => 
                           rst, Q => registers_25_29_port, QN => net108256);
   registers_reg_25_28_inst : DFFR_X1 port map( D => n3235, CK => n575, RN => 
                           rst, Q => registers_25_28_port, QN => net108255);
   registers_reg_25_27_inst : DFFR_X1 port map( D => n3234, CK => n582, RN => 
                           rst, Q => registers_25_27_port, QN => net108254);
   registers_reg_25_26_inst : DFFR_X1 port map( D => n3233, CK => n547, RN => 
                           rst, Q => registers_25_26_port, QN => net108253);
   registers_reg_25_25_inst : DFFR_X1 port map( D => n3232, CK => n563, RN => 
                           rst, Q => registers_25_25_port, QN => net108252);
   registers_reg_25_24_inst : DFFR_X1 port map( D => n3231, CK => n585, RN => 
                           rst, Q => registers_25_24_port, QN => net108251);
   registers_reg_25_23_inst : DFFR_X1 port map( D => n3230, CK => n550, RN => 
                           rst, Q => registers_25_23_port, QN => net108250);
   registers_reg_25_22_inst : DFFR_X1 port map( D => n3229, CK => n566, RN => 
                           rst, Q => registers_25_22_port, QN => net108249);
   registers_reg_25_21_inst : DFFR_X1 port map( D => n3228, CK => n621, RN => 
                           rst, Q => registers_25_21_port, QN => net108248);
   registers_reg_25_20_inst : DFFR_X1 port map( D => n3227, CK => n553, RN => 
                           rst, Q => registers_25_20_port, QN => net108247);
   registers_reg_25_19_inst : DFFR_X1 port map( D => n3226, CK => n615, RN => 
                           rst, Q => registers_25_19_port, QN => net108246);
   registers_reg_25_18_inst : DFFR_X1 port map( D => n3225, CK => n623, RN => 
                           rst, Q => registers_25_18_port, QN => net108245);
   registers_reg_25_17_inst : DFFR_X1 port map( D => n3224, CK => n628, RN => 
                           rst, Q => registers_25_17_port, QN => net108244);
   registers_reg_25_16_inst : DFFR_X1 port map( D => n3223, CK => n630, RN => 
                           rst, Q => registers_25_16_port, QN => net108243);
   registers_reg_25_15_inst : DFFR_X1 port map( D => n3222, CK => n557, RN => 
                           rst, Q => registers_25_15_port, QN => net108242);
   registers_reg_25_14_inst : DFFR_X1 port map( D => n3221, CK => n597, RN => 
                           rst, Q => registers_25_14_port, QN => net108241);
   registers_reg_25_13_inst : DFFR_X1 port map( D => n3220, CK => n600, RN => 
                           rst, Q => registers_25_13_port, QN => net108240);
   registers_reg_25_12_inst : DFFR_X1 port map( D => n3219, CK => n603, RN => 
                           rst, Q => registers_25_12_port, QN => net108239);
   registers_reg_25_11_inst : DFFR_X1 port map( D => n3218, CK => n592, RN => 
                           rst, Q => registers_25_11_port, QN => net108238);
   registers_reg_25_10_inst : DFFR_X1 port map( D => n3217, CK => n609, RN => 
                           rst, Q => registers_25_10_port, QN => net108237);
   registers_reg_25_9_inst : DFFR_X1 port map( D => n3216, CK => n587, RN => 
                           rst, Q => registers_25_9_port, QN => net108236);
   registers_reg_25_8_inst : DFFR_X1 port map( D => n3215, CK => n560, RN => 
                           rst, Q => registers_25_8_port, QN => net108235);
   registers_reg_25_7_inst : DFFR_X1 port map( D => n3214, CK => n545, RN => 
                           rst, Q => registers_25_7_port, QN => net108234);
   registers_reg_25_6_inst : DFFR_X1 port map( D => n3213, CK => n594, RN => 
                           rst, Q => registers_25_6_port, QN => net108233);
   registers_reg_25_5_inst : DFFR_X1 port map( D => n3212, CK => n556, RN => 
                           rst, Q => registers_25_5_port, QN => net108232);
   registers_reg_25_4_inst : DFFR_X1 port map( D => n3211, CK => n618, RN => 
                           rst, Q => registers_25_4_port, QN => net108231);
   registers_reg_25_3_inst : DFFR_X1 port map( D => n3210, CK => n611, RN => 
                           rst, Q => registers_25_3_port, QN => net108230);
   registers_reg_25_2_inst : DFFR_X1 port map( D => n3209, CK => n606, RN => 
                           rst, Q => registers_25_2_port, QN => net108229);
   registers_reg_25_1_inst : DFFR_X1 port map( D => n3208, CK => n634, RN => 
                           rst, Q => registers_25_1_port, QN => net108228);
   registers_reg_25_0_inst : DFFR_X1 port map( D => n3207, CK => n578, RN => 
                           rst, Q => registers_25_0_port, QN => net108227);
   registers_reg_26_31_inst : DFFR_X1 port map( D => n3206, CK => n590, RN => 
                           rst, Q => registers_26_31_port, QN => n2);
   registers_reg_26_30_inst : DFFR_X1 port map( D => n3205, CK => n569, RN => 
                           rst, Q => registers_26_30_port, QN => n4);
   registers_reg_26_29_inst : DFFR_X1 port map( D => n3204, CK => n572, RN => 
                           rst, Q => registers_26_29_port, QN => n6);
   registers_reg_26_28_inst : DFFR_X1 port map( D => n3203, CK => n575, RN => 
                           rst, Q => registers_26_28_port, QN => n8);
   registers_reg_26_27_inst : DFFR_X1 port map( D => n3202, CK => n582, RN => 
                           rst, Q => registers_26_27_port, QN => n10);
   registers_reg_26_26_inst : DFFR_X1 port map( D => n3201, CK => n547, RN => 
                           rst, Q => registers_26_26_port, QN => n12);
   registers_reg_26_25_inst : DFFR_X1 port map( D => n3200, CK => n563, RN => 
                           rst, Q => registers_26_25_port, QN => n14);
   registers_reg_26_24_inst : DFFR_X1 port map( D => n3199, CK => n585, RN => 
                           rst, Q => registers_26_24_port, QN => n16);
   registers_reg_26_23_inst : DFFR_X1 port map( D => n3198, CK => n550, RN => 
                           rst, Q => registers_26_23_port, QN => n18_port);
   registers_reg_26_22_inst : DFFR_X1 port map( D => n3197, CK => n565, RN => 
                           rst, Q => registers_26_22_port, QN => n20);
   registers_reg_26_21_inst : DFFR_X1 port map( D => n3196, CK => n621, RN => 
                           rst, Q => registers_26_21_port, QN => n22);
   registers_reg_26_20_inst : DFFR_X1 port map( D => n3195, CK => n553, RN => 
                           rst, Q => registers_26_20_port, QN => n24);
   registers_reg_26_19_inst : DFFR_X1 port map( D => n3194, CK => n615, RN => 
                           rst, Q => registers_26_19_port, QN => n26);
   registers_reg_26_18_inst : DFFR_X1 port map( D => n3193, CK => n623, RN => 
                           rst, Q => registers_26_18_port, QN => n28);
   registers_reg_26_17_inst : DFFR_X1 port map( D => n3192, CK => n628, RN => 
                           rst, Q => registers_26_17_port, QN => n30);
   registers_reg_26_16_inst : DFFR_X1 port map( D => n3191, CK => n630, RN => 
                           rst, Q => registers_26_16_port, QN => n32);
   registers_reg_26_15_inst : DFFR_X1 port map( D => n3190, CK => n557, RN => 
                           rst, Q => registers_26_15_port, QN => n34);
   registers_reg_26_14_inst : DFFR_X1 port map( D => n3189, CK => n597, RN => 
                           rst, Q => registers_26_14_port, QN => n36);
   registers_reg_26_13_inst : DFFR_X1 port map( D => n3188, CK => n600, RN => 
                           rst, Q => registers_26_13_port, QN => n38);
   registers_reg_26_12_inst : DFFR_X1 port map( D => n3187, CK => n603, RN => 
                           rst, Q => registers_26_12_port, QN => n40);
   registers_reg_26_11_inst : DFFR_X1 port map( D => n3186, CK => n597, RN => 
                           rst, Q => registers_26_11_port, QN => n42);
   registers_reg_26_10_inst : DFFR_X1 port map( D => n3185, CK => n609, RN => 
                           rst, Q => registers_26_10_port, QN => n44);
   registers_reg_26_9_inst : DFFR_X1 port map( D => n3184, CK => n587, RN => 
                           rst, Q => registers_26_9_port, QN => n46);
   registers_reg_26_8_inst : DFFR_X1 port map( D => n3183, CK => n560, RN => 
                           rst, Q => registers_26_8_port, QN => n48);
   registers_reg_26_7_inst : DFFR_X1 port map( D => n3182, CK => n545, RN => 
                           rst, Q => registers_26_7_port, QN => n50);
   registers_reg_26_6_inst : DFFR_X1 port map( D => n3181, CK => n594, RN => 
                           rst, Q => registers_26_6_port, QN => n52);
   registers_reg_26_5_inst : DFFR_X1 port map( D => n3180, CK => n556, RN => 
                           rst, Q => registers_26_5_port, QN => n54);
   registers_reg_26_4_inst : DFFR_X1 port map( D => n3179, CK => n618, RN => 
                           rst, Q => registers_26_4_port, QN => n56);
   registers_reg_26_3_inst : DFFR_X1 port map( D => n3178, CK => n611, RN => 
                           rst, Q => registers_26_3_port, QN => n58);
   registers_reg_26_2_inst : DFFR_X1 port map( D => n3177, CK => n606, RN => 
                           rst, Q => registers_26_2_port, QN => n60);
   registers_reg_26_1_inst : DFFR_X1 port map( D => n3176, CK => n632, RN => 
                           rst, Q => registers_26_1_port, QN => n62);
   registers_reg_26_0_inst : DFFR_X1 port map( D => n3175, CK => n578, RN => 
                           rst, Q => registers_26_0_port, QN => n64);
   registers_reg_27_31_inst : DFFR_X1 port map( D => n3174, CK => n590, RN => 
                           rst, Q => registers_27_31_port, QN => n416);
   registers_reg_27_30_inst : DFFR_X1 port map( D => n3173, CK => n569, RN => 
                           rst, Q => registers_27_30_port, QN => n418);
   registers_reg_27_29_inst : DFFR_X1 port map( D => n3172, CK => n572, RN => 
                           rst, Q => registers_27_29_port, QN => n420);
   registers_reg_27_28_inst : DFFR_X1 port map( D => n3171, CK => n575, RN => 
                           rst, Q => registers_27_28_port, QN => n422);
   registers_reg_27_27_inst : DFFR_X1 port map( D => n3170, CK => n582, RN => 
                           rst, Q => registers_27_27_port, QN => n424);
   registers_reg_27_26_inst : DFFR_X1 port map( D => n3169, CK => n547, RN => 
                           rst, Q => registers_27_26_port, QN => n426);
   registers_reg_27_25_inst : DFFR_X1 port map( D => n3168, CK => n563, RN => 
                           rst, Q => registers_27_25_port, QN => n428);
   registers_reg_27_24_inst : DFFR_X1 port map( D => n3167, CK => n584, RN => 
                           rst, Q => registers_27_24_port, QN => n430);
   registers_reg_27_23_inst : DFFR_X1 port map( D => n3166, CK => n550, RN => 
                           rst, Q => registers_27_23_port, QN => n432);
   registers_reg_27_22_inst : DFFR_X1 port map( D => n3165, CK => n565, RN => 
                           rst, Q => registers_27_22_port, QN => n434);
   registers_reg_27_21_inst : DFFR_X1 port map( D => n3164, CK => n621, RN => 
                           rst, Q => registers_27_21_port, QN => n436);
   registers_reg_27_20_inst : DFFR_X1 port map( D => n3163, CK => n553, RN => 
                           rst, Q => registers_27_20_port, QN => n438);
   registers_reg_27_19_inst : DFFR_X1 port map( D => n3162, CK => n615, RN => 
                           rst, Q => registers_27_19_port, QN => n440);
   registers_reg_27_18_inst : DFFR_X1 port map( D => n3161, CK => n623, RN => 
                           rst, Q => registers_27_18_port, QN => n442);
   registers_reg_27_17_inst : DFFR_X1 port map( D => n3160, CK => n627, RN => 
                           rst, Q => registers_27_17_port, QN => n444);
   registers_reg_27_16_inst : DFFR_X1 port map( D => n3159, CK => n630, RN => 
                           rst, Q => registers_27_16_port, QN => n446);
   registers_reg_27_15_inst : DFFR_X1 port map( D => n3158, CK => n557, RN => 
                           rst, Q => registers_27_15_port, QN => n448);
   registers_reg_27_14_inst : DFFR_X1 port map( D => n3157, CK => n597, RN => 
                           rst, Q => registers_27_14_port, QN => n450);
   registers_reg_27_13_inst : DFFR_X1 port map( D => n3156, CK => n600, RN => 
                           rst, Q => registers_27_13_port, QN => n452);
   registers_reg_27_12_inst : DFFR_X1 port map( D => n3155, CK => n603, RN => 
                           rst, Q => registers_27_12_port, QN => n454);
   registers_reg_27_11_inst : DFFR_X1 port map( D => n3154, CK => n614, RN => 
                           rst, Q => registers_27_11_port, QN => n456);
   registers_reg_27_10_inst : DFFR_X1 port map( D => n3153, CK => n608, RN => 
                           rst, Q => registers_27_10_port, QN => n458);
   registers_reg_27_9_inst : DFFR_X1 port map( D => n3152, CK => n587, RN => 
                           rst, Q => registers_27_9_port, QN => n460);
   registers_reg_27_8_inst : DFFR_X1 port map( D => n3151, CK => n560, RN => 
                           rst, Q => registers_27_8_port, QN => n462);
   registers_reg_27_7_inst : DFFR_X1 port map( D => n3150, CK => n550, RN => 
                           rst, Q => registers_27_7_port, QN => n464);
   registers_reg_27_6_inst : DFFR_X1 port map( D => n3149, CK => n594, RN => 
                           rst, Q => registers_27_6_port, QN => n466);
   registers_reg_27_5_inst : DFFR_X1 port map( D => n3148, CK => n556, RN => 
                           rst, Q => registers_27_5_port, QN => n468);
   registers_reg_27_4_inst : DFFR_X1 port map( D => n3147, CK => n618, RN => 
                           rst, Q => registers_27_4_port, QN => n470);
   registers_reg_27_3_inst : DFFR_X1 port map( D => n3146, CK => n611, RN => 
                           rst, Q => registers_27_3_port, QN => n472);
   registers_reg_27_2_inst : DFFR_X1 port map( D => n3145, CK => n606, RN => 
                           rst, Q => registers_27_2_port, QN => n474);
   registers_reg_27_1_inst : DFFR_X1 port map( D => n3144, CK => n634, RN => 
                           rst, Q => registers_27_1_port, QN => n476);
   registers_reg_27_0_inst : DFFR_X1 port map( D => n3143, CK => n578, RN => 
                           rst, Q => registers_27_0_port, QN => n478);
   registers_reg_28_31_inst : DFFR_X1 port map( D => n3142, CK => n590, RN => 
                           rst, Q => registers_28_31_port, QN => net108226);
   registers_reg_28_30_inst : DFFR_X1 port map( D => n3141, CK => n569, RN => 
                           rst, Q => registers_28_30_port, QN => net108225);
   registers_reg_28_29_inst : DFFR_X1 port map( D => n3140, CK => n572, RN => 
                           rst, Q => registers_28_29_port, QN => net108224);
   registers_reg_28_28_inst : DFFR_X1 port map( D => n3139, CK => n575, RN => 
                           rst, Q => registers_28_28_port, QN => net108223);
   registers_reg_28_27_inst : DFFR_X1 port map( D => n3138, CK => n582, RN => 
                           rst, Q => registers_28_27_port, QN => net108222);
   registers_reg_28_26_inst : DFFR_X1 port map( D => n3137, CK => n547, RN => 
                           rst, Q => registers_28_26_port, QN => net108221);
   registers_reg_28_25_inst : DFFR_X1 port map( D => n3136, CK => n563, RN => 
                           rst, Q => registers_28_25_port, QN => net108220);
   registers_reg_28_24_inst : DFFR_X1 port map( D => n3135, CK => n584, RN => 
                           rst, Q => registers_28_24_port, QN => net108219);
   registers_reg_28_23_inst : DFFR_X1 port map( D => n3134, CK => n550, RN => 
                           rst, Q => registers_28_23_port, QN => net108218);
   registers_reg_28_22_inst : DFFR_X1 port map( D => n3133, CK => n565, RN => 
                           rst, Q => registers_28_22_port, QN => net108217);
   registers_reg_28_21_inst : DFFR_X1 port map( D => n3132, CK => n620, RN => 
                           rst, Q => registers_28_21_port, QN => net108216);
   registers_reg_28_20_inst : DFFR_X1 port map( D => n3131, CK => n553, RN => 
                           rst, Q => registers_28_20_port, QN => net108215);
   registers_reg_28_19_inst : DFFR_X1 port map( D => n3130, CK => n615, RN => 
                           rst, Q => registers_28_19_port, QN => net108214);
   registers_reg_28_18_inst : DFFR_X1 port map( D => n3129, CK => n623, RN => 
                           rst, Q => registers_28_18_port, QN => net108213);
   registers_reg_28_17_inst : DFFR_X1 port map( D => n3128, CK => n627, RN => 
                           rst, Q => registers_28_17_port, QN => net108212);
   registers_reg_28_16_inst : DFFR_X1 port map( D => n3127, CK => n630, RN => 
                           rst, Q => registers_28_16_port, QN => net108211);
   registers_reg_28_15_inst : DFFR_X1 port map( D => n3126, CK => n557, RN => 
                           rst, Q => registers_28_15_port, QN => net108210);
   registers_reg_28_14_inst : DFFR_X1 port map( D => n3125, CK => n597, RN => 
                           rst, Q => registers_28_14_port, QN => net108209);
   registers_reg_28_13_inst : DFFR_X1 port map( D => n3124, CK => n600, RN => 
                           rst, Q => registers_28_13_port, QN => net108208);
   registers_reg_28_12_inst : DFFR_X1 port map( D => n3123, CK => n602, RN => 
                           rst, Q => registers_28_12_port, QN => net108207);
   registers_reg_28_11_inst : DFFR_X1 port map( D => n3122, CK => n614, RN => 
                           rst, Q => registers_28_11_port, QN => net108206);
   registers_reg_28_10_inst : DFFR_X1 port map( D => n3121, CK => n608, RN => 
                           rst, Q => registers_28_10_port, QN => net108205);
   registers_reg_28_9_inst : DFFR_X1 port map( D => n3120, CK => n587, RN => 
                           rst, Q => registers_28_9_port, QN => net108204);
   registers_reg_28_8_inst : DFFR_X1 port map( D => n3119, CK => n560, RN => 
                           rst, Q => registers_28_8_port, QN => net108203);
   registers_reg_28_7_inst : DFFR_X1 port map( D => n3118, CK => n568, RN => 
                           rst, Q => registers_28_7_port, QN => net108202);
   registers_reg_28_6_inst : DFFR_X1 port map( D => n3117, CK => n594, RN => 
                           rst, Q => registers_28_6_port, QN => net108201);
   registers_reg_28_5_inst : DFFR_X1 port map( D => n3116, CK => n555, RN => 
                           rst, Q => registers_28_5_port, QN => net108200);
   registers_reg_28_4_inst : DFFR_X1 port map( D => n3115, CK => n618, RN => 
                           rst, Q => registers_28_4_port, QN => net108199);
   registers_reg_28_3_inst : DFFR_X1 port map( D => n3114, CK => n611, RN => 
                           rst, Q => registers_28_3_port, QN => net108198);
   registers_reg_28_2_inst : DFFR_X1 port map( D => n3113, CK => n606, RN => 
                           rst, Q => registers_28_2_port, QN => net108197);
   registers_reg_28_1_inst : DFFR_X1 port map( D => n3112, CK => n633, RN => 
                           rst, Q => registers_28_1_port, QN => net108196);
   registers_reg_28_0_inst : DFFR_X1 port map( D => n3111, CK => n578, RN => 
                           rst, Q => registers_28_0_port, QN => net108195);
   registers_reg_29_31_inst : DFFR_X1 port map( D => n3110, CK => n590, RN => 
                           rst, Q => registers_29_31_port, QN => n161);
   registers_reg_29_30_inst : DFFR_X1 port map( D => n3109, CK => n569, RN => 
                           rst, Q => registers_29_30_port, QN => n164);
   registers_reg_29_29_inst : DFFR_X1 port map( D => n3108, CK => n572, RN => 
                           rst, Q => registers_29_29_port, QN => n166);
   registers_reg_29_28_inst : DFFR_X1 port map( D => n3107, CK => n575, RN => 
                           rst, Q => registers_29_28_port, QN => n168);
   registers_reg_29_27_inst : DFFR_X1 port map( D => n3106, CK => n582, RN => 
                           rst, Q => registers_29_27_port, QN => n170);
   registers_reg_29_26_inst : DFFR_X1 port map( D => n3105, CK => n547, RN => 
                           rst, Q => registers_29_26_port, QN => n172);
   registers_reg_29_25_inst : DFFR_X1 port map( D => n3104, CK => n562, RN => 
                           rst, Q => registers_29_25_port, QN => n174);
   registers_reg_29_24_inst : DFFR_X1 port map( D => n3103, CK => n584, RN => 
                           rst, Q => registers_29_24_port, QN => n176);
   registers_reg_29_23_inst : DFFR_X1 port map( D => n3102, CK => n550, RN => 
                           rst, Q => registers_29_23_port, QN => n178);
   registers_reg_29_22_inst : DFFR_X1 port map( D => n3101, CK => n565, RN => 
                           rst, Q => registers_29_22_port, QN => n180);
   registers_reg_29_21_inst : DFFR_X1 port map( D => n3100, CK => n620, RN => 
                           rst, Q => registers_29_21_port, QN => n182);
   registers_reg_29_20_inst : DFFR_X1 port map( D => n3099, CK => n553, RN => 
                           rst, Q => registers_29_20_port, QN => n184);
   registers_reg_29_19_inst : DFFR_X1 port map( D => n3098, CK => n615, RN => 
                           rst, Q => registers_29_19_port, QN => n186);
   registers_reg_29_18_inst : DFFR_X1 port map( D => n3097, CK => n623, RN => 
                           rst, Q => registers_29_18_port, QN => n188);
   registers_reg_29_17_inst : DFFR_X1 port map( D => n3096, CK => n627, RN => 
                           rst, Q => registers_29_17_port, QN => n190);
   registers_reg_29_16_inst : DFFR_X1 port map( D => n3095, CK => n630, RN => 
                           rst, Q => registers_29_16_port, QN => n192);
   registers_reg_29_15_inst : DFFR_X1 port map( D => n3094, CK => n557, RN => 
                           rst, Q => registers_29_15_port, QN => n194);
   registers_reg_29_14_inst : DFFR_X1 port map( D => n3093, CK => n597, RN => 
                           rst, Q => registers_29_14_port, QN => n196);
   registers_reg_29_13_inst : DFFR_X1 port map( D => n3092, CK => n600, RN => 
                           rst, Q => registers_29_13_port, QN => n198);
   registers_reg_29_12_inst : DFFR_X1 port map( D => n3091, CK => n602, RN => 
                           rst, Q => registers_29_12_port, QN => n200);
   registers_reg_29_11_inst : DFFR_X1 port map( D => n3090, CK => n614, RN => 
                           rst, Q => registers_29_11_port, QN => n202);
   registers_reg_29_10_inst : DFFR_X1 port map( D => n3089, CK => n608, RN => 
                           rst, Q => registers_29_10_port, QN => n204);
   registers_reg_29_9_inst : DFFR_X1 port map( D => n3088, CK => n587, RN => 
                           rst, Q => registers_29_9_port, QN => n206);
   registers_reg_29_8_inst : DFFR_X1 port map( D => n3087, CK => n560, RN => 
                           rst, Q => registers_29_8_port, QN => n208);
   registers_reg_29_7_inst : DFFR_X1 port map( D => n3086, CK => n568, RN => 
                           rst, Q => registers_29_7_port, QN => n210);
   registers_reg_29_6_inst : DFFR_X1 port map( D => n3085, CK => n594, RN => 
                           rst, Q => registers_29_6_port, QN => n212);
   registers_reg_29_5_inst : DFFR_X1 port map( D => n3084, CK => n555, RN => 
                           rst, Q => registers_29_5_port, QN => n214);
   registers_reg_29_4_inst : DFFR_X1 port map( D => n3083, CK => n618, RN => 
                           rst, Q => registers_29_4_port, QN => n216);
   registers_reg_29_3_inst : DFFR_X1 port map( D => n3082, CK => n611, RN => 
                           rst, Q => registers_29_3_port, QN => n218);
   registers_reg_29_2_inst : DFFR_X1 port map( D => n3081, CK => n605, RN => 
                           rst, Q => registers_29_2_port, QN => n220);
   registers_reg_29_1_inst : DFFR_X1 port map( D => n3080, CK => n634, RN => 
                           rst, Q => registers_29_1_port, QN => n222);
   registers_reg_29_0_inst : DFFR_X1 port map( D => n3079, CK => n577, RN => 
                           rst, Q => registers_29_0_port, QN => n224);
   registers_reg_30_31_inst : DFFR_X1 port map( D => n3078, CK => n590, RN => 
                           rst, Q => registers_30_31_port, QN => net108194);
   registers_reg_30_30_inst : DFFR_X1 port map( D => n3077, CK => n569, RN => 
                           rst, Q => registers_30_30_port, QN => net108193);
   registers_reg_30_29_inst : DFFR_X1 port map( D => n3076, CK => n572, RN => 
                           rst, Q => registers_30_29_port, QN => net108192);
   registers_reg_30_28_inst : DFFR_X1 port map( D => n3075, CK => n574, RN => 
                           rst, Q => registers_30_28_port, QN => net108191);
   registers_reg_30_27_inst : DFFR_X1 port map( D => n3074, CK => n581, RN => 
                           rst, Q => registers_30_27_port, QN => net108190);
   registers_reg_30_26_inst : DFFR_X1 port map( D => n3073, CK => n547, RN => 
                           rst, Q => registers_30_26_port, QN => net108189);
   registers_reg_30_25_inst : DFFR_X1 port map( D => n3072, CK => n562, RN => 
                           rst, Q => registers_30_25_port, QN => net108188);
   registers_reg_30_24_inst : DFFR_X1 port map( D => n3071, CK => n584, RN => 
                           rst, Q => registers_30_24_port, QN => net108187);
   registers_reg_30_23_inst : DFFR_X1 port map( D => n3070, CK => n550, RN => 
                           rst, Q => registers_30_23_port, QN => net108186);
   registers_reg_30_22_inst : DFFR_X1 port map( D => n3069, CK => n565, RN => 
                           rst, Q => registers_30_22_port, QN => net108185);
   registers_reg_30_21_inst : DFFR_X1 port map( D => n3068, CK => n620, RN => 
                           rst, Q => registers_30_21_port, QN => net108184);
   registers_reg_30_20_inst : DFFR_X1 port map( D => n3067, CK => n553, RN => 
                           rst, Q => registers_30_20_port, QN => net108183);
   registers_reg_30_19_inst : DFFR_X1 port map( D => n3066, CK => n615, RN => 
                           rst, Q => registers_30_19_port, QN => net108182);
   registers_reg_30_18_inst : DFFR_X1 port map( D => n3065, CK => n623, RN => 
                           rst, Q => registers_30_18_port, QN => net108181);
   registers_reg_30_17_inst : DFFR_X1 port map( D => n3064, CK => n627, RN => 
                           rst, Q => registers_30_17_port, QN => net108180);
   registers_reg_30_16_inst : DFFR_X1 port map( D => n3063, CK => n630, RN => 
                           rst, Q => registers_30_16_port, QN => net108179);
   registers_reg_30_15_inst : DFFR_X1 port map( D => n3062, CK => n557, RN => 
                           rst, Q => registers_30_15_port, QN => net108178);
   registers_reg_30_14_inst : DFFR_X1 port map( D => n3061, CK => n597, RN => 
                           rst, Q => registers_30_14_port, QN => net108177);
   registers_reg_30_13_inst : DFFR_X1 port map( D => n3060, CK => n600, RN => 
                           rst, Q => registers_30_13_port, QN => net108176);
   registers_reg_30_12_inst : DFFR_X1 port map( D => n3059, CK => n602, RN => 
                           rst, Q => registers_30_12_port, QN => net108175);
   registers_reg_30_11_inst : DFFR_X1 port map( D => n3058, CK => n614, RN => 
                           rst, Q => registers_30_11_port, QN => net108174);
   registers_reg_30_10_inst : DFFR_X1 port map( D => n3057, CK => n608, RN => 
                           rst, Q => registers_30_10_port, QN => net108173);
   registers_reg_30_9_inst : DFFR_X1 port map( D => n3056, CK => n587, RN => 
                           rst, Q => registers_30_9_port, QN => net108172);
   registers_reg_30_8_inst : DFFR_X1 port map( D => n3055, CK => n560, RN => 
                           rst, Q => registers_30_8_port, QN => net108171);
   registers_reg_30_7_inst : DFFR_X1 port map( D => n3054, CK => n568, RN => 
                           rst, Q => registers_30_7_port, QN => net108170);
   registers_reg_30_6_inst : DFFR_X1 port map( D => n3053, CK => n594, RN => 
                           rst, Q => registers_30_6_port, QN => net108169);
   registers_reg_30_5_inst : DFFR_X1 port map( D => n3052, CK => n555, RN => 
                           rst, Q => registers_30_5_port, QN => net108168);
   registers_reg_30_4_inst : DFFR_X1 port map( D => n3051, CK => n617, RN => 
                           rst, Q => registers_30_4_port, QN => net108167);
   registers_reg_30_3_inst : DFFR_X1 port map( D => n3050, CK => n611, RN => 
                           rst, Q => registers_30_3_port, QN => net108166);
   registers_reg_30_2_inst : DFFR_X1 port map( D => n3049, CK => n605, RN => 
                           rst, Q => registers_30_2_port, QN => net108165);
   registers_reg_30_1_inst : DFFR_X1 port map( D => n3048, CK => n634, RN => 
                           rst, Q => registers_30_1_port, QN => net108164);
   registers_reg_30_0_inst : DFFR_X1 port map( D => n3047, CK => n577, RN => 
                           rst, Q => registers_30_0_port, QN => net108163);
   registers_reg_31_31_inst : DFFR_X1 port map( D => n3046, CK => n603, RN => 
                           rst, Q => net108162, QN => n289);
   d_out2_reg_31_inst : DFF_X1 port map( D => n3045, CK => n636, Q => 
                           d_out2_31_port, QN => net108161);
   registers_reg_31_30_inst : DFFR_X1 port map( D => n3044, CK => n603, RN => 
                           rst, Q => registers_31_30_port, QN => n322);
   d_out2_reg_30_inst : DFF_X1 port map( D => n3043, CK => n635, Q => 
                           d_out2_30_port, QN => n2949);
   registers_reg_31_29_inst : DFFR_X1 port map( D => n3042, CK => n603, RN => 
                           rst, Q => registers_31_29_port, QN => n323);
   d_out2_reg_29_inst : DFF_X1 port map( D => n3041, CK => n635, Q => 
                           d_out2_29_port, QN => n2948);
   registers_reg_31_28_inst : DFFR_X1 port map( D => n3040, CK => n577, RN => 
                           rst, Q => registers_31_28_port, QN => n324);
   d_out2_reg_28_inst : DFF_X1 port map( D => n3039, CK => n639, Q => 
                           d_out2_28_port, QN => n2947);
   registers_reg_31_27_inst : DFFR_X1 port map( D => n3038, CK => n603, RN => 
                           rst, Q => registers_31_27_port, QN => n325);
   d_out2_reg_27_inst : DFF_X1 port map( D => n3037, CK => n635, Q => 
                           d_out2_27_port, QN => n2946);
   registers_reg_31_26_inst : DFFR_X1 port map( D => n3036, CK => n603, RN => 
                           rst, Q => registers_31_26_port, QN => n326);
   d_out2_reg_26_inst : DFF_X1 port map( D => n3035, CK => n635, Q => 
                           d_out2_26_port, QN => n2945);
   registers_reg_31_25_inst : DFFR_X1 port map( D => n3034, CK => n603, RN => 
                           rst, Q => registers_31_25_port, QN => n327);
   d_out2_reg_25_inst : DFF_X1 port map( D => n3033, CK => n636, Q => 
                           d_out2_25_port, QN => n2944);
   registers_reg_31_24_inst : DFFR_X1 port map( D => n3032, CK => n603, RN => 
                           rst, Q => registers_31_24_port, QN => n328);
   d_out2_reg_24_inst : DFF_X1 port map( D => n3031, CK => n635, Q => 
                           d_out2_24_port, QN => n2943);
   registers_reg_31_23_inst : DFFR_X1 port map( D => n3030, CK => n604, RN => 
                           rst, Q => registers_31_23_port, QN => n329);
   d_out2_reg_23_inst : DFF_X1 port map( D => n3029, CK => n635, Q => 
                           d_out2_23_port, QN => n2942);
   registers_reg_31_22_inst : DFFR_X1 port map( D => n3028, CK => n604, RN => 
                           rst, Q => registers_31_22_port, QN => n330);
   d_out2_reg_22_inst : DFF_X1 port map( D => n3027, CK => n635, Q => 
                           d_out2_22_port, QN => n2941);
   registers_reg_31_21_inst : DFFR_X1 port map( D => n3026, CK => n604, RN => 
                           rst, Q => registers_31_21_port, QN => n331);
   d_out2_reg_21_inst : DFF_X1 port map( D => n3025, CK => n636, Q => 
                           d_out2_21_port, QN => n2940);
   registers_reg_31_20_inst : DFFR_X1 port map( D => n3024, CK => n603, RN => 
                           rst, Q => registers_31_20_port, QN => n332);
   d_out2_reg_20_inst : DFF_X1 port map( D => n3023, CK => n637, Q => 
                           d_out2_20_port, QN => n2939);
   registers_reg_31_19_inst : DFFR_X1 port map( D => n3022, CK => n604, RN => 
                           rst, Q => registers_31_19_port, QN => n333);
   d_out2_reg_19_inst : DFF_X1 port map( D => n3021, CK => n636, Q => 
                           d_out2_19_port, QN => n2938);
   registers_reg_31_18_inst : DFFR_X1 port map( D => n3020, CK => n604, RN => 
                           rst, Q => registers_31_18_port, QN => n334);
   d_out2_reg_18_inst : DFF_X1 port map( D => n3019, CK => n636, Q => 
                           d_out2_18_port, QN => n2937);
   registers_reg_31_17_inst : DFFR_X1 port map( D => n3018, CK => n604, RN => 
                           rst, Q => registers_31_17_port, QN => n335);
   d_out2_reg_17_inst : DFF_X1 port map( D => n3017, CK => n636, Q => 
                           d_out2_17_port, QN => n2936);
   registers_reg_31_16_inst : DFFR_X1 port map( D => n3016, CK => n604, RN => 
                           rst, Q => registers_31_16_port, QN => n336);
   d_out2_reg_16_inst : DFF_X1 port map( D => n3015, CK => n635, Q => 
                           d_out2_16_port, QN => n2935);
   registers_reg_31_15_inst : DFFR_X1 port map( D => n3014, CK => n604, RN => 
                           rst, Q => registers_31_15_port, QN => n337);
   d_out2_reg_15_inst : DFF_X1 port map( D => n3013, CK => n637, Q => 
                           d_out2_15_port, QN => n2934);
   registers_reg_31_14_inst : DFFR_X1 port map( D => n3012, CK => n604, RN => 
                           rst, Q => registers_31_14_port, QN => n338);
   d_out2_reg_14_inst : DFF_X1 port map( D => n3011, CK => n637, Q => 
                           d_out2_14_port, QN => n2933);
   registers_reg_31_13_inst : DFFR_X1 port map( D => n3010, CK => n604, RN => 
                           rst, Q => registers_31_13_port, QN => n339);
   d_out2_reg_13_inst : DFF_X1 port map( D => n3009, CK => n637, Q => 
                           d_out2_13_port, QN => n2932);
   registers_reg_31_12_inst : DFFR_X1 port map( D => n3008, CK => n604, RN => 
                           rst, Q => registers_31_12_port, QN => n340);
   d_out2_reg_12_inst : DFF_X1 port map( D => n3007, CK => n637, Q => 
                           d_out2_12_port, QN => n2931);
   registers_reg_31_11_inst : DFFR_X1 port map( D => n3006, CK => n605, RN => 
                           rst, Q => registers_31_11_port, QN => n341);
   d_out2_reg_11_inst : DFF_X1 port map( D => n3005, CK => n638, Q => 
                           d_out2_11_port, QN => n2930);
   registers_reg_31_10_inst : DFFR_X1 port map( D => n3004, CK => n605, RN => 
                           rst, Q => registers_31_10_port, QN => n342);
   d_out2_reg_10_inst : DFF_X1 port map( D => n3003, CK => n638, Q => 
                           d_out2_10_port, QN => n2929);
   registers_reg_31_9_inst : DFFR_X1 port map( D => n3002, CK => n605, RN => 
                           rst, Q => registers_31_9_port, QN => n343);
   d_out2_reg_9_inst : DFF_X1 port map( D => n3001, CK => n638, Q => 
                           d_out2_9_port, QN => n2928);
   registers_reg_31_8_inst : DFFR_X1 port map( D => n3000, CK => n605, RN => 
                           rst, Q => registers_31_8_port, QN => n344);
   d_out2_reg_8_inst : DFF_X1 port map( D => n2999, CK => n637, Q => 
                           d_out2_8_port, QN => n2927);
   registers_reg_31_7_inst : DFFR_X1 port map( D => n2998, CK => n605, RN => 
                           rst, Q => registers_31_7_port, QN => n345);
   d_out2_reg_7_inst : DFF_X1 port map( D => n2997, CK => n638, Q => 
                           d_out2_7_port, QN => n2926);
   registers_reg_31_6_inst : DFFR_X1 port map( D => n2996, CK => n605, RN => 
                           rst, Q => registers_31_6_port, QN => n346);
   d_out2_reg_6_inst : DFF_X1 port map( D => n2995, CK => n638, Q => 
                           d_out2_6_port, QN => n2925);
   registers_reg_31_5_inst : DFFR_X1 port map( D => n2994, CK => n605, RN => 
                           rst, Q => registers_31_5_port, QN => n347);
   d_out2_reg_5_inst : DFF_X1 port map( D => n2993, CK => n638, Q => 
                           d_out2_5_port, QN => n2924);
   registers_reg_31_4_inst : DFFR_X1 port map( D => n2992, CK => n605, RN => 
                           rst, Q => registers_31_4_port, QN => n348);
   d_out2_reg_4_inst : DFF_X1 port map( D => n2991, CK => n638, Q => 
                           d_out2_4_port, QN => n2923);
   registers_reg_31_3_inst : DFFR_X1 port map( D => n2990, CK => n605, RN => 
                           rst, Q => registers_31_3_port, QN => n349);
   d_out2_reg_3_inst : DFF_X1 port map( D => n2989, CK => n639, Q => 
                           d_out2_3_port, QN => n2922);
   registers_reg_31_2_inst : DFFR_X1 port map( D => n2988, CK => n608, RN => 
                           rst, Q => registers_31_2_port, QN => n350);
   d_out2_reg_2_inst : DFF_X1 port map( D => n2987, CK => n639, Q => 
                           d_out2_2_port, QN => n2921);
   registers_reg_31_1_inst : DFFR_X1 port map( D => n2986, CK => n634, RN => 
                           rst, Q => registers_31_1_port, QN => n351);
   d_out2_reg_1_inst : DFF_X1 port map( D => n2985, CK => n639, Q => 
                           d_out2_1_port, QN => n2920);
   registers_reg_31_0_inst : DFFR_X1 port map( D => n2984, CK => n577, RN => 
                           rst, Q => registers_31_0_port, QN => n352);
   d_out2_reg_0_inst : DFF_X1 port map( D => n2983, CK => n637, Q => 
                           d_out2_0_port, QN => n2919);
   d_out1_reg_31_inst : DFF_X1 port map( D => n2982, CK => n636, Q => 
                           d_out1_31_port, QN => net108160);
   d_out1_reg_30_inst : DFF_X1 port map( D => n2981, CK => n640, Q => 
                           d_out1_30_port, QN => net108159);
   d_out1_reg_29_inst : DFF_X1 port map( D => n2980, CK => n640, Q => 
                           d_out1_29_port, QN => net108158);
   d_out1_reg_28_inst : DFF_X1 port map( D => n2979, CK => n637, Q => 
                           d_out1_28_port, QN => net108157);
   d_out1_reg_27_inst : DFF_X1 port map( D => n2978, CK => n639, Q => 
                           d_out1_27_port, QN => net108156);
   d_out1_reg_26_inst : DFF_X1 port map( D => n2977, CK => n640, Q => 
                           d_out1_26_port, QN => net108155);
   d_out1_reg_25_inst : DFF_X1 port map( D => n2976, CK => n640, Q => 
                           d_out1_25_port, QN => net108154);
   d_out1_reg_24_inst : DFF_X1 port map( D => n2975, CK => n640, Q => 
                           d_out1_24_port, QN => net108153);
   d_out1_reg_23_inst : DFF_X1 port map( D => n2974, CK => n640, Q => 
                           d_out1_23_port, QN => net108152);
   d_out1_reg_22_inst : DFF_X1 port map( D => n2973, CK => n639, Q => 
                           d_out1_22_port, QN => net108151);
   d_out1_reg_21_inst : DFF_X1 port map( D => n2972, CK => n640, Q => 
                           d_out1_21_port, QN => net108150);
   d_out1_reg_20_inst : DFF_X1 port map( D => n2971, CK => n638, Q => 
                           d_out1_20_port, QN => net108149);
   d_out1_reg_19_inst : DFF_X1 port map( D => n2970, CK => n636, Q => 
                           d_out1_19_port, QN => net108148);
   d_out1_reg_18_inst : DFF_X1 port map( D => n2969, CK => n638, Q => 
                           d_out1_18_port, QN => net108147);
   d_out1_reg_17_inst : DFF_X1 port map( D => n2968, CK => n639, Q => 
                           d_out1_17_port, QN => net108146);
   d_out1_reg_16_inst : DFF_X1 port map( D => n2967, CK => n640, Q => 
                           d_out1_16_port, QN => net108145);
   d_out1_reg_15_inst : DFF_X1 port map( D => n2966, CK => n636, Q => 
                           d_out1_15_port, QN => net108144);
   d_out1_reg_14_inst : DFF_X1 port map( D => n2965, CK => n637, Q => 
                           d_out1_14_port, QN => net108143);
   d_out1_reg_13_inst : DFF_X1 port map( D => n2964, CK => n639, Q => 
                           d_out1_13_port, QN => net108142);
   d_out1_reg_12_inst : DFF_X1 port map( D => n2963, CK => n636, Q => 
                           d_out1_12_port, QN => net108141);
   d_out1_reg_11_inst : DFF_X1 port map( D => n2962, CK => n637, Q => 
                           d_out1_11_port, QN => net108140);
   d_out1_reg_10_inst : DFF_X1 port map( D => n2961, CK => n640, Q => 
                           d_out1_10_port, QN => net108139);
   d_out1_reg_9_inst : DFF_X1 port map( D => n2960, CK => n638, Q => 
                           d_out1_9_port, QN => net108138);
   d_out1_reg_8_inst : DFF_X1 port map( D => n2959, CK => n639, Q => 
                           d_out1_8_port, QN => net108137);
   d_out1_reg_7_inst : DFF_X1 port map( D => n2958, CK => n637, Q => 
                           d_out1_7_port, QN => net108136);
   d_out1_reg_6_inst : DFF_X1 port map( D => n2957, CK => n638, Q => 
                           d_out1_6_port, QN => net108135);
   d_out1_reg_5_inst : DFF_X1 port map( D => n2956, CK => n635, Q => 
                           d_out1_5_port, QN => net108134);
   d_out1_reg_4_inst : DFF_X1 port map( D => n2955, CK => n640, Q => 
                           d_out1_4_port, QN => net108133);
   d_out1_reg_3_inst : DFF_X1 port map( D => n2954, CK => n640, Q => 
                           d_out1_3_port, QN => net108132);
   d_out1_reg_2_inst : DFF_X1 port map( D => n2953, CK => n639, Q => 
                           d_out1_2_port, QN => net108131);
   d_out1_reg_1_inst : DFF_X1 port map( D => n2952, CK => n639, Q => 
                           d_out1_1_port, QN => net108130);
   d_out1_reg_0_inst : DFF_X1 port map( D => n2951, CK => n636, Q => 
                           d_out1_0_port, QN => net108129);
   U3 : NOR2_X4 port map( A1 => n2030, A2 => n1466, ZN => n1465);
   U4 : NOR2_X4 port map( A1 => n1397, A2 => link_en, ZN => n709);
   U5 : AND2_X2 port map( A1 => n658, A2 => n659, ZN => n657);
   U6 : AND2_X2 port map( A1 => n668, A2 => n669, ZN => n667);
   U7 : AND2_X2 port map( A1 => n2026, A2 => n2020, ZN => n1489);
   U8 : AND2_X2 port map( A1 => n2024, A2 => n2012, ZN => n1479);
   U9 : AND2_X2 port map( A1 => n1416, A2 => n1406, ZN => n760);
   U10 : AND2_X2 port map( A1 => n661, A2 => n659, ZN => n660);
   U11 : AND2_X2 port map( A1 => n669, A2 => n658, ZN => n670);
   U12 : AND2_X2 port map( A1 => n1408, A2 => n1407, ZN => n715);
   U13 : AND2_X2 port map( A1 => n2026, A2 => n2015, ZN => n1494);
   U14 : AND2_X2 port map( A1 => n1418, A2 => n1403, ZN => n745);
   U15 : NAND2_X2 port map( A1 => n1416, A2 => n1412, ZN => n753);
   U16 : NAND2_X2 port map( A1 => n2024, A2 => n2020, ZN => n1486);
   U17 : AND2_X2 port map( A1 => n663, A2 => n659, ZN => n662);
   U18 : AND2_X2 port map( A1 => n669, A2 => n661, ZN => n671);
   U19 : AND2_X2 port map( A1 => n674, A2 => n668, ZN => n673);
   U20 : AND2_X2 port map( A1 => n2020, A2 => n2014, ZN => n1454);
   U21 : AND3_X2 port map( A1 => n2013, A2 => n2019, A3 => n2026, ZN => n1459);
   U22 : NAND2_X2 port map( A1 => n1418, A2 => n1405, ZN => n748);
   U23 : NAND2_X2 port map( A1 => n2024, A2 => n2015, ZN => n1491);
   U24 : NAND2_X2 port map( A1 => n1416, A2 => n1408, ZN => n758);
   U25 : AND2_X2 port map( A1 => n669, A2 => n663, ZN => n672);
   U26 : AND2_X2 port map( A1 => n674, A2 => n661, ZN => n676);
   U27 : AND2_X2 port map( A1 => n679, A2 => n658, ZN => n680);
   U28 : AND3_X2 port map( A1 => n1406, A2 => n771, A3 => n1418, ZN => n726);
   U29 : NAND2_X2 port map( A1 => n1407, A2 => n1405, ZN => n731);
   U30 : NAND2_X2 port map( A1 => n2014, A2 => n2012, ZN => n1464);
   U31 : AND2_X2 port map( A1 => n1416, A2 => n1410, ZN => n755);
   U32 : AND3_X2 port map( A1 => n2023, A2 => n2019, A3 => n2026, ZN => n1460);
   U33 : NAND2_X2 port map( A1 => n2024, A2 => n2010, ZN => n1475);
   U34 : AND2_X2 port map( A1 => n674, A2 => n663, ZN => n677);
   U35 : AND2_X2 port map( A1 => n679, A2 => n661, ZN => n681);
   U36 : AND2_X2 port map( A1 => n686, A2 => n658, ZN => n687);
   U37 : AND2_X2 port map( A1 => n692, A2 => n668, ZN => n691);
   U38 : AND2_X2 port map( A1 => n1412, A2 => n1407, ZN => n721);
   U39 : AND2_X2 port map( A1 => n2015, A2 => n2014, ZN => n1448);
   U40 : NAND2_X2 port map( A1 => n1403, A2 => n1404, ZN => n720);
   U41 : NAND2_X2 port map( A1 => n2010, A2 => n2011, ZN => n1453);
   U42 : NAND2_X2 port map( A1 => n2026, A2 => n2012, ZN => n1481);
   U43 : NAND2_X2 port map( A1 => n2017, A2 => n2018, ZN => n1476);
   U44 : AND2_X2 port map( A1 => n1415, A2 => n1414, ZN => n750);
   U45 : AND2_X2 port map( A1 => n1418, A2 => n1408, ZN => n761);
   U46 : AND2_X2 port map( A1 => n1416, A2 => n1405, ZN => n746);
   U47 : NAND3_X2 port map( A1 => n2024, A2 => n2019, A3 => n2025, ZN => n1462)
                           ;
   U48 : AND2_X2 port map( A1 => n674, A2 => n658, ZN => n675);
   U49 : AND2_X2 port map( A1 => n679, A2 => n663, ZN => n682);
   U50 : AND2_X2 port map( A1 => n686, A2 => n661, ZN => n688);
   U51 : AND2_X2 port map( A1 => n697, A2 => n668, ZN => n696);
   U52 : NAND2_X2 port map( A1 => n1410, A2 => n1411, ZN => n743);
   U53 : AND2_X2 port map( A1 => n1406, A2 => n1404, ZN => n716);
   U54 : AND2_X2 port map( A1 => n1403, A2 => n1407, ZN => n722);
   U55 : AND2_X2 port map( A1 => n2010, A2 => n2014, ZN => n1455);
   U56 : AND2_X2 port map( A1 => n2013, A2 => n2011, ZN => n1449);
   U57 : AND3_X2 port map( A1 => n1415, A2 => n771, A3 => n1418, ZN => n727);
   U58 : NAND2_X2 port map( A1 => n2023, A2 => n2018, ZN => n1480);
   U59 : NAND3_X2 port map( A1 => n1416, A2 => n771, A3 => n1417, ZN => n729);
   U60 : NAND3_X2 port map( A1 => n2025, A2 => n2019, A3 => n2026, ZN => n1470)
                           ;
   U61 : AND2_X2 port map( A1 => n2024, A2 => n2017, ZN => n1488);
   U62 : AND2_X2 port map( A1 => n686, A2 => n663, ZN => n689);
   U63 : AND2_X2 port map( A1 => n692, A2 => n661, ZN => n694);
   U64 : AND2_X2 port map( A1 => n697, A2 => n658, ZN => n698);
   U65 : AND2_X2 port map( A1 => n702, A2 => n668, ZN => n701);
   U66 : NAND2_X2 port map( A1 => n1408, A2 => n1404, ZN => n724);
   U67 : NAND2_X2 port map( A1 => n2015, A2 => n2011, ZN => n1457);
   U68 : NAND2_X2 port map( A1 => n1406, A2 => n1407, ZN => n718);
   U69 : NAND2_X2 port map( A1 => n2013, A2 => n2014, ZN => n1451);
   U70 : NAND2_X2 port map( A1 => n2025, A2 => n2022, ZN => n1485);
   U71 : NAND2_X2 port map( A1 => n2026, A2 => n2017, ZN => n1490);
   U72 : NAND2_X2 port map( A1 => n1418, A2 => n1410, ZN => n757);
   U73 : AND2_X2 port map( A1 => n1417, A2 => n1411, ZN => n751);
   U74 : NAND3_X2 port map( A1 => n1415, A2 => n771, A3 => n1416, ZN => n730);
   U75 : NAND3_X2 port map( A1 => n2023, A2 => n2019, A3 => n2024, ZN => n1463)
                           ;
   U76 : AND2_X2 port map( A1 => n679, A2 => n668, ZN => n678);
   U77 : AND2_X2 port map( A1 => n692, A2 => n663, ZN => n695);
   U78 : AND2_X2 port map( A1 => n697, A2 => n661, ZN => n699);
   U79 : AND2_X2 port map( A1 => n702, A2 => n658, ZN => n703);
   U80 : INV_X2 port map( A => n732, ZN => n776);
   U81 : INV_X2 port map( A => n737, ZN => n770);
   U82 : INV_X2 port map( A => n733, ZN => n774);
   U83 : AND2_X2 port map( A1 => n2025, A2 => n2018, ZN => n1484);
   U84 : AND2_X2 port map( A1 => link_en, A2 => n707, ZN => n710);
   U85 : NAND2_X2 port map( A1 => n1416, A2 => n1403, ZN => n742);
   U86 : NAND2_X2 port map( A1 => n1410, A2 => n1407, ZN => n725);
   U87 : NAND2_X2 port map( A1 => n2017, A2 => n2014, ZN => n1458);
   U88 : NAND2_X2 port map( A1 => n1405, A2 => n1404, ZN => n719);
   U89 : NAND2_X2 port map( A1 => n2012, A2 => n2011, ZN => n1452);
   U90 : AND2_X2 port map( A1 => n1418, A2 => n1412, ZN => n756);
   U91 : AND2_X2 port map( A1 => n2023, A2 => n2022, ZN => n1483);
   U92 : AND2_X2 port map( A1 => n2024, A2 => n2013, ZN => n1493);
   U93 : AND2_X2 port map( A1 => n2026, A2 => n2010, ZN => n1478);
   U94 : NAND2_X2 port map( A1 => n1415, A2 => n1411, ZN => n747);
   U95 : NAND2_X2 port map( A1 => n1417, A2 => n1414, ZN => n752);
   U96 : NAND2_X2 port map( A1 => n2029, A2 => n2030, ZN => n1469);
   U97 : INV_X2 port map( A => n1397, ZN => n707);
   U98 : AND2_X2 port map( A1 => n686, A2 => n668, ZN => n685);
   U99 : AND2_X2 port map( A1 => n692, A2 => n658, ZN => n693);
   U100 : AND2_X2 port map( A1 => n697, A2 => n663, ZN => n700);
   U101 : AND2_X2 port map( A1 => n702, A2 => n661, ZN => n705);
   U102 : INV_X2 port map( A => n736, ZN => n771);
   U103 : NAND3_X2 port map( A1 => rst, A2 => en, A3 => rd1_en, ZN => n1466);
   U104 : BUF_X1 port map( A => N18, Z => n641);
   U105 : BUF_X1 port map( A => N18, Z => n646);
   U106 : BUF_X1 port map( A => N18, Z => n645);
   U107 : BUF_X1 port map( A => N18, Z => n648);
   U108 : BUF_X1 port map( A => N18, Z => n647);
   U109 : BUF_X1 port map( A => N18, Z => n642);
   U110 : BUF_X1 port map( A => N18, Z => n654);
   U111 : BUF_X1 port map( A => N18, Z => n644);
   U112 : BUF_X1 port map( A => N18, Z => n643);
   U113 : BUF_X1 port map( A => N18, Z => n655);
   U114 : BUF_X1 port map( A => N18, Z => n649);
   U115 : BUF_X1 port map( A => N18, Z => n653);
   U116 : BUF_X1 port map( A => N18, Z => n656);
   U117 : BUF_X1 port map( A => N18, Z => n650);
   U118 : BUF_X1 port map( A => N18, Z => n651);
   U119 : BUF_X1 port map( A => N18, Z => n652);
   U120 : CLKBUF_X1 port map( A => n656, Z => n545);
   U121 : CLKBUF_X1 port map( A => n656, Z => n546);
   U122 : CLKBUF_X1 port map( A => n656, Z => n547);
   U123 : CLKBUF_X1 port map( A => n656, Z => n548);
   U124 : CLKBUF_X1 port map( A => n656, Z => n549);
   U125 : CLKBUF_X1 port map( A => n656, Z => n550);
   U126 : CLKBUF_X1 port map( A => n655, Z => n551);
   U127 : CLKBUF_X1 port map( A => n655, Z => n552);
   U128 : CLKBUF_X1 port map( A => n655, Z => n553);
   U129 : CLKBUF_X1 port map( A => n655, Z => n554);
   U130 : CLKBUF_X1 port map( A => n655, Z => n555);
   U131 : CLKBUF_X1 port map( A => n655, Z => n556);
   U132 : CLKBUF_X1 port map( A => n654, Z => n557);
   U133 : CLKBUF_X1 port map( A => n654, Z => n558);
   U134 : CLKBUF_X1 port map( A => n654, Z => n559);
   U135 : CLKBUF_X1 port map( A => n654, Z => n560);
   U136 : CLKBUF_X1 port map( A => n654, Z => n561);
   U137 : CLKBUF_X1 port map( A => n654, Z => n562);
   U138 : CLKBUF_X1 port map( A => n653, Z => n563);
   U139 : CLKBUF_X1 port map( A => n653, Z => n564);
   U140 : CLKBUF_X1 port map( A => n653, Z => n565);
   U141 : CLKBUF_X1 port map( A => n653, Z => n566);
   U142 : CLKBUF_X1 port map( A => n653, Z => n567);
   U143 : CLKBUF_X1 port map( A => n653, Z => n568);
   U144 : CLKBUF_X1 port map( A => n652, Z => n569);
   U145 : CLKBUF_X1 port map( A => n652, Z => n570);
   U146 : CLKBUF_X1 port map( A => n652, Z => n571);
   U147 : CLKBUF_X1 port map( A => n652, Z => n572);
   U148 : CLKBUF_X1 port map( A => n652, Z => n573);
   U149 : CLKBUF_X1 port map( A => n652, Z => n574);
   U150 : CLKBUF_X1 port map( A => n651, Z => n575);
   U151 : CLKBUF_X1 port map( A => n651, Z => n576);
   U152 : CLKBUF_X1 port map( A => n651, Z => n577);
   U153 : CLKBUF_X1 port map( A => n651, Z => n578);
   U154 : CLKBUF_X1 port map( A => n651, Z => n579);
   U155 : CLKBUF_X1 port map( A => n651, Z => n580);
   U156 : CLKBUF_X1 port map( A => n650, Z => n581);
   U157 : CLKBUF_X1 port map( A => n650, Z => n582);
   U158 : CLKBUF_X1 port map( A => n650, Z => n583);
   U159 : CLKBUF_X1 port map( A => n650, Z => n584);
   U160 : CLKBUF_X1 port map( A => n650, Z => n585);
   U161 : CLKBUF_X1 port map( A => n650, Z => n586);
   U162 : CLKBUF_X1 port map( A => n649, Z => n587);
   U163 : CLKBUF_X1 port map( A => n649, Z => n588);
   U164 : CLKBUF_X1 port map( A => n649, Z => n589);
   U165 : CLKBUF_X1 port map( A => n649, Z => n590);
   U166 : CLKBUF_X1 port map( A => n649, Z => n591);
   U167 : CLKBUF_X1 port map( A => n649, Z => n592);
   U168 : CLKBUF_X1 port map( A => n648, Z => n593);
   U169 : CLKBUF_X1 port map( A => n648, Z => n594);
   U170 : CLKBUF_X1 port map( A => n648, Z => n595);
   U171 : CLKBUF_X1 port map( A => n648, Z => n596);
   U172 : CLKBUF_X1 port map( A => n648, Z => n597);
   U173 : CLKBUF_X1 port map( A => n648, Z => n598);
   U174 : CLKBUF_X1 port map( A => n647, Z => n599);
   U175 : CLKBUF_X1 port map( A => n647, Z => n600);
   U176 : CLKBUF_X1 port map( A => n647, Z => n601);
   U177 : CLKBUF_X1 port map( A => n647, Z => n602);
   U178 : CLKBUF_X1 port map( A => n647, Z => n603);
   U179 : CLKBUF_X1 port map( A => n647, Z => n604);
   U180 : CLKBUF_X1 port map( A => n646, Z => n605);
   U181 : CLKBUF_X1 port map( A => n646, Z => n606);
   U182 : CLKBUF_X1 port map( A => n646, Z => n607);
   U183 : CLKBUF_X1 port map( A => n646, Z => n608);
   U184 : CLKBUF_X1 port map( A => n646, Z => n609);
   U185 : CLKBUF_X1 port map( A => n646, Z => n610);
   U186 : CLKBUF_X1 port map( A => n645, Z => n611);
   U187 : CLKBUF_X1 port map( A => n645, Z => n612);
   U188 : CLKBUF_X1 port map( A => n645, Z => n613);
   U189 : CLKBUF_X1 port map( A => n645, Z => n614);
   U190 : CLKBUF_X1 port map( A => n645, Z => n615);
   U191 : CLKBUF_X1 port map( A => n645, Z => n616);
   U192 : CLKBUF_X1 port map( A => n644, Z => n617);
   U193 : CLKBUF_X1 port map( A => n644, Z => n618);
   U194 : CLKBUF_X1 port map( A => n644, Z => n619);
   U195 : CLKBUF_X1 port map( A => n644, Z => n620);
   U196 : CLKBUF_X1 port map( A => n644, Z => n621);
   U197 : CLKBUF_X1 port map( A => n644, Z => n622);
   U198 : CLKBUF_X1 port map( A => n643, Z => n623);
   U199 : CLKBUF_X1 port map( A => n643, Z => n624);
   U200 : CLKBUF_X1 port map( A => n643, Z => n625);
   U201 : CLKBUF_X1 port map( A => n643, Z => n626);
   U202 : CLKBUF_X1 port map( A => n643, Z => n627);
   U203 : CLKBUF_X1 port map( A => n643, Z => n628);
   U204 : CLKBUF_X1 port map( A => n642, Z => n629);
   U205 : CLKBUF_X1 port map( A => n642, Z => n630);
   U206 : CLKBUF_X1 port map( A => n642, Z => n631);
   U207 : CLKBUF_X1 port map( A => n642, Z => n632);
   U208 : CLKBUF_X1 port map( A => n642, Z => n633);
   U209 : CLKBUF_X1 port map( A => n642, Z => n634);
   U210 : CLKBUF_X1 port map( A => n641, Z => n635);
   U211 : CLKBUF_X1 port map( A => n641, Z => n636);
   U212 : CLKBUF_X1 port map( A => n641, Z => n637);
   U213 : CLKBUF_X1 port map( A => n641, Z => n638);
   U214 : CLKBUF_X1 port map( A => n641, Z => n639);
   U215 : CLKBUF_X1 port map( A => n641, Z => n640);
   U216 : MUX2_X1 port map( A => registers_1_31_port, B => d_in(31), S => n657,
                           Z => n4006);
   U217 : MUX2_X1 port map( A => registers_1_30_port, B => d_in(30), S => n657,
                           Z => n4005);
   U218 : MUX2_X1 port map( A => registers_1_29_port, B => d_in(29), S => n657,
                           Z => n4004);
   U219 : MUX2_X1 port map( A => registers_1_28_port, B => d_in(28), S => n657,
                           Z => n4003);
   U220 : MUX2_X1 port map( A => registers_1_27_port, B => d_in(27), S => n657,
                           Z => n4002);
   U221 : MUX2_X1 port map( A => registers_1_26_port, B => d_in(26), S => n657,
                           Z => n4001);
   U222 : MUX2_X1 port map( A => registers_1_25_port, B => d_in(25), S => n657,
                           Z => n4000);
   U223 : MUX2_X1 port map( A => registers_1_24_port, B => d_in(24), S => n657,
                           Z => n3999);
   U224 : MUX2_X1 port map( A => registers_1_23_port, B => d_in(23), S => n657,
                           Z => n3998);
   U225 : MUX2_X1 port map( A => registers_1_22_port, B => d_in(22), S => n657,
                           Z => n3997);
   U226 : MUX2_X1 port map( A => registers_1_21_port, B => d_in(21), S => n657,
                           Z => n3996);
   U227 : MUX2_X1 port map( A => registers_1_20_port, B => d_in(20), S => n657,
                           Z => n3995);
   U228 : MUX2_X1 port map( A => registers_1_19_port, B => d_in(19), S => n657,
                           Z => n3994);
   U229 : MUX2_X1 port map( A => registers_1_18_port, B => d_in(18), S => n657,
                           Z => n3993);
   U230 : MUX2_X1 port map( A => registers_1_17_port, B => d_in(17), S => n657,
                           Z => n3992);
   U231 : MUX2_X1 port map( A => registers_1_16_port, B => d_in(16), S => n657,
                           Z => n3991);
   U232 : MUX2_X1 port map( A => registers_1_15_port, B => d_in(15), S => n657,
                           Z => n3990);
   U233 : MUX2_X1 port map( A => registers_1_14_port, B => d_in(14), S => n657,
                           Z => n3989);
   U234 : MUX2_X1 port map( A => registers_1_13_port, B => d_in(13), S => n657,
                           Z => n3988);
   U235 : MUX2_X1 port map( A => registers_1_12_port, B => d_in(12), S => n657,
                           Z => n3987);
   U236 : MUX2_X1 port map( A => registers_1_11_port, B => d_in(11), S => n657,
                           Z => n3986);
   U237 : MUX2_X1 port map( A => registers_1_10_port, B => d_in(10), S => n657,
                           Z => n3985);
   U238 : MUX2_X1 port map( A => registers_1_9_port, B => d_in(9), S => n657, Z
                           => n3984);
   U239 : MUX2_X1 port map( A => registers_1_8_port, B => d_in(8), S => n657, Z
                           => n3983);
   U240 : MUX2_X1 port map( A => registers_1_7_port, B => d_in(7), S => n657, Z
                           => n3982);
   U241 : MUX2_X1 port map( A => registers_1_6_port, B => d_in(6), S => n657, Z
                           => n3981);
   U242 : MUX2_X1 port map( A => registers_1_5_port, B => d_in(5), S => n657, Z
                           => n3980);
   U243 : MUX2_X1 port map( A => registers_1_4_port, B => d_in(4), S => n657, Z
                           => n3979);
   U244 : MUX2_X1 port map( A => registers_1_3_port, B => d_in(3), S => n657, Z
                           => n3978);
   U245 : MUX2_X1 port map( A => registers_1_2_port, B => d_in(2), S => n657, Z
                           => n3977);
   U246 : MUX2_X1 port map( A => registers_1_1_port, B => d_in(1), S => n657, Z
                           => n3976);
   U247 : MUX2_X1 port map( A => registers_1_0_port, B => d_in(0), S => n657, Z
                           => n3975);
   U248 : MUX2_X1 port map( A => registers_2_31_port, B => d_in(31), S => n660,
                           Z => n3974);
   U249 : MUX2_X1 port map( A => registers_2_30_port, B => d_in(30), S => n660,
                           Z => n3973);
   U250 : MUX2_X1 port map( A => registers_2_29_port, B => d_in(29), S => n660,
                           Z => n3972);
   U251 : MUX2_X1 port map( A => registers_2_28_port, B => d_in(28), S => n660,
                           Z => n3971);
   U252 : MUX2_X1 port map( A => registers_2_27_port, B => d_in(27), S => n660,
                           Z => n3970);
   U253 : MUX2_X1 port map( A => registers_2_26_port, B => d_in(26), S => n660,
                           Z => n3969);
   U254 : MUX2_X1 port map( A => registers_2_25_port, B => d_in(25), S => n660,
                           Z => n3968);
   U255 : MUX2_X1 port map( A => registers_2_24_port, B => d_in(24), S => n660,
                           Z => n3967);
   U256 : MUX2_X1 port map( A => registers_2_23_port, B => d_in(23), S => n660,
                           Z => n3966);
   U257 : MUX2_X1 port map( A => registers_2_22_port, B => d_in(22), S => n660,
                           Z => n3965);
   U258 : MUX2_X1 port map( A => registers_2_21_port, B => d_in(21), S => n660,
                           Z => n3964);
   U259 : MUX2_X1 port map( A => registers_2_20_port, B => d_in(20), S => n660,
                           Z => n3963);
   U260 : MUX2_X1 port map( A => registers_2_19_port, B => d_in(19), S => n660,
                           Z => n3962);
   U261 : MUX2_X1 port map( A => registers_2_18_port, B => d_in(18), S => n660,
                           Z => n3961);
   U262 : MUX2_X1 port map( A => registers_2_17_port, B => d_in(17), S => n660,
                           Z => n3960);
   U263 : MUX2_X1 port map( A => registers_2_16_port, B => d_in(16), S => n660,
                           Z => n3959);
   U264 : MUX2_X1 port map( A => registers_2_15_port, B => d_in(15), S => n660,
                           Z => n3958);
   U265 : MUX2_X1 port map( A => registers_2_14_port, B => d_in(14), S => n660,
                           Z => n3957);
   U266 : MUX2_X1 port map( A => registers_2_13_port, B => d_in(13), S => n660,
                           Z => n3956);
   U267 : MUX2_X1 port map( A => registers_2_12_port, B => d_in(12), S => n660,
                           Z => n3955);
   U268 : MUX2_X1 port map( A => registers_2_11_port, B => d_in(11), S => n660,
                           Z => n3954);
   U269 : MUX2_X1 port map( A => registers_2_10_port, B => d_in(10), S => n660,
                           Z => n3953);
   U270 : MUX2_X1 port map( A => registers_2_9_port, B => d_in(9), S => n660, Z
                           => n3952);
   U271 : MUX2_X1 port map( A => registers_2_8_port, B => d_in(8), S => n660, Z
                           => n3951);
   U272 : MUX2_X1 port map( A => registers_2_7_port, B => d_in(7), S => n660, Z
                           => n3950);
   U273 : MUX2_X1 port map( A => registers_2_6_port, B => d_in(6), S => n660, Z
                           => n3949);
   U274 : MUX2_X1 port map( A => registers_2_5_port, B => d_in(5), S => n660, Z
                           => n3948);
   U275 : MUX2_X1 port map( A => registers_2_4_port, B => d_in(4), S => n660, Z
                           => n3947);
   U276 : MUX2_X1 port map( A => registers_2_3_port, B => d_in(3), S => n660, Z
                           => n3946);
   U277 : MUX2_X1 port map( A => registers_2_2_port, B => d_in(2), S => n660, Z
                           => n3945);
   U278 : MUX2_X1 port map( A => registers_2_1_port, B => d_in(1), S => n660, Z
                           => n3944);
   U279 : MUX2_X1 port map( A => registers_2_0_port, B => d_in(0), S => n660, Z
                           => n3943);
   U280 : MUX2_X1 port map( A => registers_3_31_port, B => d_in(31), S => n662,
                           Z => n3942);
   U281 : MUX2_X1 port map( A => registers_3_30_port, B => d_in(30), S => n662,
                           Z => n3941);
   U282 : MUX2_X1 port map( A => registers_3_29_port, B => d_in(29), S => n662,
                           Z => n3940);
   U283 : MUX2_X1 port map( A => registers_3_28_port, B => d_in(28), S => n662,
                           Z => n3939);
   U284 : MUX2_X1 port map( A => registers_3_27_port, B => d_in(27), S => n662,
                           Z => n3938);
   U285 : MUX2_X1 port map( A => registers_3_26_port, B => d_in(26), S => n662,
                           Z => n3937);
   U286 : MUX2_X1 port map( A => registers_3_25_port, B => d_in(25), S => n662,
                           Z => n3936);
   U287 : MUX2_X1 port map( A => registers_3_24_port, B => d_in(24), S => n662,
                           Z => n3935);
   U288 : MUX2_X1 port map( A => registers_3_23_port, B => d_in(23), S => n662,
                           Z => n3934);
   U289 : MUX2_X1 port map( A => registers_3_22_port, B => d_in(22), S => n662,
                           Z => n3933);
   U290 : MUX2_X1 port map( A => registers_3_21_port, B => d_in(21), S => n662,
                           Z => n3932);
   U291 : MUX2_X1 port map( A => registers_3_20_port, B => d_in(20), S => n662,
                           Z => n3931);
   U292 : MUX2_X1 port map( A => registers_3_19_port, B => d_in(19), S => n662,
                           Z => n3930);
   U293 : MUX2_X1 port map( A => registers_3_18_port, B => d_in(18), S => n662,
                           Z => n3929);
   U294 : MUX2_X1 port map( A => registers_3_17_port, B => d_in(17), S => n662,
                           Z => n3928);
   U295 : MUX2_X1 port map( A => registers_3_16_port, B => d_in(16), S => n662,
                           Z => n3927);
   U296 : MUX2_X1 port map( A => registers_3_15_port, B => d_in(15), S => n662,
                           Z => n3926);
   U297 : MUX2_X1 port map( A => registers_3_14_port, B => d_in(14), S => n662,
                           Z => n3925);
   U298 : MUX2_X1 port map( A => registers_3_13_port, B => d_in(13), S => n662,
                           Z => n3924);
   U299 : MUX2_X1 port map( A => registers_3_12_port, B => d_in(12), S => n662,
                           Z => n3923);
   U300 : MUX2_X1 port map( A => registers_3_11_port, B => d_in(11), S => n662,
                           Z => n3922);
   U301 : MUX2_X1 port map( A => registers_3_10_port, B => d_in(10), S => n662,
                           Z => n3921);
   U302 : MUX2_X1 port map( A => registers_3_9_port, B => d_in(9), S => n662, Z
                           => n3920);
   U303 : MUX2_X1 port map( A => registers_3_8_port, B => d_in(8), S => n662, Z
                           => n3919);
   U304 : MUX2_X1 port map( A => registers_3_7_port, B => d_in(7), S => n662, Z
                           => n3918);
   U305 : MUX2_X1 port map( A => registers_3_6_port, B => d_in(6), S => n662, Z
                           => n3917);
   U306 : MUX2_X1 port map( A => registers_3_5_port, B => d_in(5), S => n662, Z
                           => n3916);
   U307 : MUX2_X1 port map( A => registers_3_4_port, B => d_in(4), S => n662, Z
                           => n3915);
   U308 : MUX2_X1 port map( A => registers_3_3_port, B => d_in(3), S => n662, Z
                           => n3914);
   U309 : MUX2_X1 port map( A => registers_3_2_port, B => d_in(2), S => n662, Z
                           => n3913);
   U310 : MUX2_X1 port map( A => registers_3_1_port, B => d_in(1), S => n662, Z
                           => n3912);
   U311 : MUX2_X1 port map( A => registers_3_0_port, B => d_in(0), S => n662, Z
                           => n3911);
   U312 : AND3_X1 port map( A1 => n664, A2 => n665, A3 => n666, ZN => n659);
   U313 : MUX2_X1 port map( A => registers_4_31_port, B => d_in(31), S => n667,
                           Z => n3910);
   U314 : MUX2_X1 port map( A => registers_4_30_port, B => d_in(30), S => n667,
                           Z => n3909);
   U315 : MUX2_X1 port map( A => registers_4_29_port, B => d_in(29), S => n667,
                           Z => n3908);
   U316 : MUX2_X1 port map( A => registers_4_28_port, B => d_in(28), S => n667,
                           Z => n3907);
   U317 : MUX2_X1 port map( A => registers_4_27_port, B => d_in(27), S => n667,
                           Z => n3906);
   U318 : MUX2_X1 port map( A => registers_4_26_port, B => d_in(26), S => n667,
                           Z => n3905);
   U319 : MUX2_X1 port map( A => registers_4_25_port, B => d_in(25), S => n667,
                           Z => n3904);
   U320 : MUX2_X1 port map( A => registers_4_24_port, B => d_in(24), S => n667,
                           Z => n3903);
   U321 : MUX2_X1 port map( A => registers_4_23_port, B => d_in(23), S => n667,
                           Z => n3902);
   U322 : MUX2_X1 port map( A => registers_4_22_port, B => d_in(22), S => n667,
                           Z => n3901);
   U323 : MUX2_X1 port map( A => registers_4_21_port, B => d_in(21), S => n667,
                           Z => n3900);
   U324 : MUX2_X1 port map( A => registers_4_20_port, B => d_in(20), S => n667,
                           Z => n3899);
   U325 : MUX2_X1 port map( A => registers_4_19_port, B => d_in(19), S => n667,
                           Z => n3898);
   U326 : MUX2_X1 port map( A => registers_4_18_port, B => d_in(18), S => n667,
                           Z => n3897);
   U327 : MUX2_X1 port map( A => registers_4_17_port, B => d_in(17), S => n667,
                           Z => n3896);
   U328 : MUX2_X1 port map( A => registers_4_16_port, B => d_in(16), S => n667,
                           Z => n3895);
   U329 : MUX2_X1 port map( A => registers_4_15_port, B => d_in(15), S => n667,
                           Z => n3894);
   U330 : MUX2_X1 port map( A => registers_4_14_port, B => d_in(14), S => n667,
                           Z => n3893);
   U331 : MUX2_X1 port map( A => registers_4_13_port, B => d_in(13), S => n667,
                           Z => n3892);
   U332 : MUX2_X1 port map( A => registers_4_12_port, B => d_in(12), S => n667,
                           Z => n3891);
   U333 : MUX2_X1 port map( A => registers_4_11_port, B => d_in(11), S => n667,
                           Z => n3890);
   U334 : MUX2_X1 port map( A => registers_4_10_port, B => d_in(10), S => n667,
                           Z => n3889);
   U335 : MUX2_X1 port map( A => registers_4_9_port, B => d_in(9), S => n667, Z
                           => n3888);
   U336 : MUX2_X1 port map( A => registers_4_8_port, B => d_in(8), S => n667, Z
                           => n3887);
   U337 : MUX2_X1 port map( A => registers_4_7_port, B => d_in(7), S => n667, Z
                           => n3886);
   U338 : MUX2_X1 port map( A => registers_4_6_port, B => d_in(6), S => n667, Z
                           => n3885);
   U339 : MUX2_X1 port map( A => registers_4_5_port, B => d_in(5), S => n667, Z
                           => n3884);
   U340 : MUX2_X1 port map( A => registers_4_4_port, B => d_in(4), S => n667, Z
                           => n3883);
   U341 : MUX2_X1 port map( A => registers_4_3_port, B => d_in(3), S => n667, Z
                           => n3882);
   U342 : MUX2_X1 port map( A => registers_4_2_port, B => d_in(2), S => n667, Z
                           => n3881);
   U343 : MUX2_X1 port map( A => registers_4_1_port, B => d_in(1), S => n667, Z
                           => n3880);
   U344 : MUX2_X1 port map( A => registers_4_0_port, B => d_in(0), S => n667, Z
                           => n3879);
   U345 : MUX2_X1 port map( A => registers_5_31_port, B => d_in(31), S => n670,
                           Z => n3878);
   U346 : MUX2_X1 port map( A => registers_5_30_port, B => d_in(30), S => n670,
                           Z => n3877);
   U347 : MUX2_X1 port map( A => registers_5_29_port, B => d_in(29), S => n670,
                           Z => n3876);
   U348 : MUX2_X1 port map( A => registers_5_28_port, B => d_in(28), S => n670,
                           Z => n3875);
   U349 : MUX2_X1 port map( A => registers_5_27_port, B => d_in(27), S => n670,
                           Z => n3874);
   U350 : MUX2_X1 port map( A => registers_5_26_port, B => d_in(26), S => n670,
                           Z => n3873);
   U351 : MUX2_X1 port map( A => registers_5_25_port, B => d_in(25), S => n670,
                           Z => n3872);
   U352 : MUX2_X1 port map( A => registers_5_24_port, B => d_in(24), S => n670,
                           Z => n3871);
   U353 : MUX2_X1 port map( A => registers_5_23_port, B => d_in(23), S => n670,
                           Z => n3870);
   U354 : MUX2_X1 port map( A => registers_5_22_port, B => d_in(22), S => n670,
                           Z => n3869);
   U355 : MUX2_X1 port map( A => registers_5_21_port, B => d_in(21), S => n670,
                           Z => n3868);
   U356 : MUX2_X1 port map( A => registers_5_20_port, B => d_in(20), S => n670,
                           Z => n3867);
   U357 : MUX2_X1 port map( A => registers_5_19_port, B => d_in(19), S => n670,
                           Z => n3866);
   U358 : MUX2_X1 port map( A => registers_5_18_port, B => d_in(18), S => n670,
                           Z => n3865);
   U359 : MUX2_X1 port map( A => registers_5_17_port, B => d_in(17), S => n670,
                           Z => n3864);
   U360 : MUX2_X1 port map( A => registers_5_16_port, B => d_in(16), S => n670,
                           Z => n3863);
   U361 : MUX2_X1 port map( A => registers_5_15_port, B => d_in(15), S => n670,
                           Z => n3862);
   U362 : MUX2_X1 port map( A => registers_5_14_port, B => d_in(14), S => n670,
                           Z => n3861);
   U363 : MUX2_X1 port map( A => registers_5_13_port, B => d_in(13), S => n670,
                           Z => n3860);
   U364 : MUX2_X1 port map( A => registers_5_12_port, B => d_in(12), S => n670,
                           Z => n3859);
   U365 : MUX2_X1 port map( A => registers_5_11_port, B => d_in(11), S => n670,
                           Z => n3858);
   U366 : MUX2_X1 port map( A => registers_5_10_port, B => d_in(10), S => n670,
                           Z => n3857);
   U367 : MUX2_X1 port map( A => registers_5_9_port, B => d_in(9), S => n670, Z
                           => n3856);
   U368 : MUX2_X1 port map( A => registers_5_8_port, B => d_in(8), S => n670, Z
                           => n3855);
   U369 : MUX2_X1 port map( A => registers_5_7_port, B => d_in(7), S => n670, Z
                           => n3854);
   U370 : MUX2_X1 port map( A => registers_5_6_port, B => d_in(6), S => n670, Z
                           => n3853);
   U371 : MUX2_X1 port map( A => registers_5_5_port, B => d_in(5), S => n670, Z
                           => n3852);
   U372 : MUX2_X1 port map( A => registers_5_4_port, B => d_in(4), S => n670, Z
                           => n3851);
   U373 : MUX2_X1 port map( A => registers_5_3_port, B => d_in(3), S => n670, Z
                           => n3850);
   U374 : MUX2_X1 port map( A => registers_5_2_port, B => d_in(2), S => n670, Z
                           => n3849);
   U375 : MUX2_X1 port map( A => registers_5_1_port, B => d_in(1), S => n670, Z
                           => n3848);
   U376 : MUX2_X1 port map( A => registers_5_0_port, B => d_in(0), S => n670, Z
                           => n3847);
   U377 : MUX2_X1 port map( A => registers_6_31_port, B => d_in(31), S => n671,
                           Z => n3846);
   U378 : MUX2_X1 port map( A => registers_6_30_port, B => d_in(30), S => n671,
                           Z => n3845);
   U379 : MUX2_X1 port map( A => registers_6_29_port, B => d_in(29), S => n671,
                           Z => n3844);
   U380 : MUX2_X1 port map( A => registers_6_28_port, B => d_in(28), S => n671,
                           Z => n3843);
   U381 : MUX2_X1 port map( A => registers_6_27_port, B => d_in(27), S => n671,
                           Z => n3842);
   U382 : MUX2_X1 port map( A => registers_6_26_port, B => d_in(26), S => n671,
                           Z => n3841);
   U383 : MUX2_X1 port map( A => registers_6_25_port, B => d_in(25), S => n671,
                           Z => n3840);
   U384 : MUX2_X1 port map( A => registers_6_24_port, B => d_in(24), S => n671,
                           Z => n3839);
   U385 : MUX2_X1 port map( A => registers_6_23_port, B => d_in(23), S => n671,
                           Z => n3838);
   U386 : MUX2_X1 port map( A => registers_6_22_port, B => d_in(22), S => n671,
                           Z => n3837);
   U387 : MUX2_X1 port map( A => registers_6_21_port, B => d_in(21), S => n671,
                           Z => n3836);
   U388 : MUX2_X1 port map( A => registers_6_20_port, B => d_in(20), S => n671,
                           Z => n3835);
   U389 : MUX2_X1 port map( A => registers_6_19_port, B => d_in(19), S => n671,
                           Z => n3834);
   U390 : MUX2_X1 port map( A => registers_6_18_port, B => d_in(18), S => n671,
                           Z => n3833);
   U391 : MUX2_X1 port map( A => registers_6_17_port, B => d_in(17), S => n671,
                           Z => n3832);
   U392 : MUX2_X1 port map( A => registers_6_16_port, B => d_in(16), S => n671,
                           Z => n3831);
   U393 : MUX2_X1 port map( A => registers_6_15_port, B => d_in(15), S => n671,
                           Z => n3830);
   U394 : MUX2_X1 port map( A => registers_6_14_port, B => d_in(14), S => n671,
                           Z => n3829);
   U395 : MUX2_X1 port map( A => registers_6_13_port, B => d_in(13), S => n671,
                           Z => n3828);
   U396 : MUX2_X1 port map( A => registers_6_12_port, B => d_in(12), S => n671,
                           Z => n3827);
   U397 : MUX2_X1 port map( A => registers_6_11_port, B => d_in(11), S => n671,
                           Z => n3826);
   U398 : MUX2_X1 port map( A => registers_6_10_port, B => d_in(10), S => n671,
                           Z => n3825);
   U399 : MUX2_X1 port map( A => registers_6_9_port, B => d_in(9), S => n671, Z
                           => n3824);
   U400 : MUX2_X1 port map( A => registers_6_8_port, B => d_in(8), S => n671, Z
                           => n3823);
   U401 : MUX2_X1 port map( A => registers_6_7_port, B => d_in(7), S => n671, Z
                           => n3822);
   U402 : MUX2_X1 port map( A => registers_6_6_port, B => d_in(6), S => n671, Z
                           => n3821);
   U403 : MUX2_X1 port map( A => registers_6_5_port, B => d_in(5), S => n671, Z
                           => n3820);
   U404 : MUX2_X1 port map( A => registers_6_4_port, B => d_in(4), S => n671, Z
                           => n3819);
   U405 : MUX2_X1 port map( A => registers_6_3_port, B => d_in(3), S => n671, Z
                           => n3818);
   U406 : MUX2_X1 port map( A => registers_6_2_port, B => d_in(2), S => n671, Z
                           => n3817);
   U407 : MUX2_X1 port map( A => registers_6_1_port, B => d_in(1), S => n671, Z
                           => n3816);
   U408 : MUX2_X1 port map( A => registers_6_0_port, B => d_in(0), S => n671, Z
                           => n3815);
   U409 : MUX2_X1 port map( A => registers_7_31_port, B => d_in(31), S => n672,
                           Z => n3814);
   U410 : MUX2_X1 port map( A => registers_7_30_port, B => d_in(30), S => n672,
                           Z => n3813);
   U411 : MUX2_X1 port map( A => registers_7_29_port, B => d_in(29), S => n672,
                           Z => n3812);
   U412 : MUX2_X1 port map( A => registers_7_28_port, B => d_in(28), S => n672,
                           Z => n3811);
   U413 : MUX2_X1 port map( A => registers_7_27_port, B => d_in(27), S => n672,
                           Z => n3810);
   U414 : MUX2_X1 port map( A => registers_7_26_port, B => d_in(26), S => n672,
                           Z => n3809);
   U415 : MUX2_X1 port map( A => registers_7_25_port, B => d_in(25), S => n672,
                           Z => n3808);
   U416 : MUX2_X1 port map( A => registers_7_24_port, B => d_in(24), S => n672,
                           Z => n3807);
   U417 : MUX2_X1 port map( A => registers_7_23_port, B => d_in(23), S => n672,
                           Z => n3806);
   U418 : MUX2_X1 port map( A => registers_7_22_port, B => d_in(22), S => n672,
                           Z => n3805);
   U419 : MUX2_X1 port map( A => registers_7_21_port, B => d_in(21), S => n672,
                           Z => n3804);
   U420 : MUX2_X1 port map( A => registers_7_20_port, B => d_in(20), S => n672,
                           Z => n3803);
   U421 : MUX2_X1 port map( A => registers_7_19_port, B => d_in(19), S => n672,
                           Z => n3802);
   U422 : MUX2_X1 port map( A => registers_7_18_port, B => d_in(18), S => n672,
                           Z => n3801);
   U423 : MUX2_X1 port map( A => registers_7_17_port, B => d_in(17), S => n672,
                           Z => n3800);
   U424 : MUX2_X1 port map( A => registers_7_16_port, B => d_in(16), S => n672,
                           Z => n3799);
   U425 : MUX2_X1 port map( A => registers_7_15_port, B => d_in(15), S => n672,
                           Z => n3798);
   U426 : MUX2_X1 port map( A => registers_7_14_port, B => d_in(14), S => n672,
                           Z => n3797);
   U427 : MUX2_X1 port map( A => registers_7_13_port, B => d_in(13), S => n672,
                           Z => n3796);
   U428 : MUX2_X1 port map( A => registers_7_12_port, B => d_in(12), S => n672,
                           Z => n3795);
   U429 : MUX2_X1 port map( A => registers_7_11_port, B => d_in(11), S => n672,
                           Z => n3794);
   U430 : MUX2_X1 port map( A => registers_7_10_port, B => d_in(10), S => n672,
                           Z => n3793);
   U431 : MUX2_X1 port map( A => registers_7_9_port, B => d_in(9), S => n672, Z
                           => n3792);
   U432 : MUX2_X1 port map( A => registers_7_8_port, B => d_in(8), S => n672, Z
                           => n3791);
   U433 : MUX2_X1 port map( A => registers_7_7_port, B => d_in(7), S => n672, Z
                           => n3790);
   U434 : MUX2_X1 port map( A => registers_7_6_port, B => d_in(6), S => n672, Z
                           => n3789);
   U435 : MUX2_X1 port map( A => registers_7_5_port, B => d_in(5), S => n672, Z
                           => n3788);
   U436 : MUX2_X1 port map( A => registers_7_4_port, B => d_in(4), S => n672, Z
                           => n3787);
   U437 : MUX2_X1 port map( A => registers_7_3_port, B => d_in(3), S => n672, Z
                           => n3786);
   U438 : MUX2_X1 port map( A => registers_7_2_port, B => d_in(2), S => n672, Z
                           => n3785);
   U439 : MUX2_X1 port map( A => registers_7_1_port, B => d_in(1), S => n672, Z
                           => n3784);
   U440 : MUX2_X1 port map( A => registers_7_0_port, B => d_in(0), S => n672, Z
                           => n3783);
   U441 : AND3_X1 port map( A1 => n666, A2 => n665, A3 => wr_addr(2), ZN => 
                           n669);
   U442 : MUX2_X1 port map( A => registers_8_31_port, B => d_in(31), S => n673,
                           Z => n3782);
   U443 : MUX2_X1 port map( A => registers_8_30_port, B => d_in(30), S => n673,
                           Z => n3781);
   U444 : MUX2_X1 port map( A => registers_8_29_port, B => d_in(29), S => n673,
                           Z => n3780);
   U445 : MUX2_X1 port map( A => registers_8_28_port, B => d_in(28), S => n673,
                           Z => n3779);
   U446 : MUX2_X1 port map( A => registers_8_27_port, B => d_in(27), S => n673,
                           Z => n3778);
   U447 : MUX2_X1 port map( A => registers_8_26_port, B => d_in(26), S => n673,
                           Z => n3777);
   U448 : MUX2_X1 port map( A => registers_8_25_port, B => d_in(25), S => n673,
                           Z => n3776);
   U449 : MUX2_X1 port map( A => registers_8_24_port, B => d_in(24), S => n673,
                           Z => n3775);
   U450 : MUX2_X1 port map( A => registers_8_23_port, B => d_in(23), S => n673,
                           Z => n3774);
   U451 : MUX2_X1 port map( A => registers_8_22_port, B => d_in(22), S => n673,
                           Z => n3773);
   U452 : MUX2_X1 port map( A => registers_8_21_port, B => d_in(21), S => n673,
                           Z => n3772);
   U453 : MUX2_X1 port map( A => registers_8_20_port, B => d_in(20), S => n673,
                           Z => n3771);
   U454 : MUX2_X1 port map( A => registers_8_19_port, B => d_in(19), S => n673,
                           Z => n3770);
   U455 : MUX2_X1 port map( A => registers_8_18_port, B => d_in(18), S => n673,
                           Z => n3769);
   U456 : MUX2_X1 port map( A => registers_8_17_port, B => d_in(17), S => n673,
                           Z => n3768);
   U457 : MUX2_X1 port map( A => registers_8_16_port, B => d_in(16), S => n673,
                           Z => n3767);
   U458 : MUX2_X1 port map( A => registers_8_15_port, B => d_in(15), S => n673,
                           Z => n3766);
   U459 : MUX2_X1 port map( A => registers_8_14_port, B => d_in(14), S => n673,
                           Z => n3765);
   U460 : MUX2_X1 port map( A => registers_8_13_port, B => d_in(13), S => n673,
                           Z => n3764);
   U461 : MUX2_X1 port map( A => registers_8_12_port, B => d_in(12), S => n673,
                           Z => n3763);
   U462 : MUX2_X1 port map( A => registers_8_11_port, B => d_in(11), S => n673,
                           Z => n3762);
   U463 : MUX2_X1 port map( A => registers_8_10_port, B => d_in(10), S => n673,
                           Z => n3761);
   U464 : MUX2_X1 port map( A => registers_8_9_port, B => d_in(9), S => n673, Z
                           => n3760);
   U465 : MUX2_X1 port map( A => registers_8_8_port, B => d_in(8), S => n673, Z
                           => n3759);
   U466 : MUX2_X1 port map( A => registers_8_7_port, B => d_in(7), S => n673, Z
                           => n3758);
   U467 : MUX2_X1 port map( A => registers_8_6_port, B => d_in(6), S => n673, Z
                           => n3757);
   U468 : MUX2_X1 port map( A => registers_8_5_port, B => d_in(5), S => n673, Z
                           => n3756);
   U469 : MUX2_X1 port map( A => registers_8_4_port, B => d_in(4), S => n673, Z
                           => n3755);
   U470 : MUX2_X1 port map( A => registers_8_3_port, B => d_in(3), S => n673, Z
                           => n3754);
   U471 : MUX2_X1 port map( A => registers_8_2_port, B => d_in(2), S => n673, Z
                           => n3753);
   U472 : MUX2_X1 port map( A => registers_8_1_port, B => d_in(1), S => n673, Z
                           => n3752);
   U473 : MUX2_X1 port map( A => registers_8_0_port, B => d_in(0), S => n673, Z
                           => n3751);
   U474 : MUX2_X1 port map( A => registers_9_31_port, B => d_in(31), S => n675,
                           Z => n3750);
   U475 : MUX2_X1 port map( A => registers_9_30_port, B => d_in(30), S => n675,
                           Z => n3749);
   U476 : MUX2_X1 port map( A => registers_9_29_port, B => d_in(29), S => n675,
                           Z => n3748);
   U477 : MUX2_X1 port map( A => registers_9_28_port, B => d_in(28), S => n675,
                           Z => n3747);
   U478 : MUX2_X1 port map( A => registers_9_27_port, B => d_in(27), S => n675,
                           Z => n3746);
   U479 : MUX2_X1 port map( A => registers_9_26_port, B => d_in(26), S => n675,
                           Z => n3745);
   U480 : MUX2_X1 port map( A => registers_9_25_port, B => d_in(25), S => n675,
                           Z => n3744);
   U481 : MUX2_X1 port map( A => registers_9_24_port, B => d_in(24), S => n675,
                           Z => n3743);
   U482 : MUX2_X1 port map( A => registers_9_23_port, B => d_in(23), S => n675,
                           Z => n3742);
   U483 : MUX2_X1 port map( A => registers_9_22_port, B => d_in(22), S => n675,
                           Z => n3741);
   U484 : MUX2_X1 port map( A => registers_9_21_port, B => d_in(21), S => n675,
                           Z => n3740);
   U485 : MUX2_X1 port map( A => registers_9_20_port, B => d_in(20), S => n675,
                           Z => n3739);
   U486 : MUX2_X1 port map( A => registers_9_19_port, B => d_in(19), S => n675,
                           Z => n3738);
   U487 : MUX2_X1 port map( A => registers_9_18_port, B => d_in(18), S => n675,
                           Z => n3737);
   U488 : MUX2_X1 port map( A => registers_9_17_port, B => d_in(17), S => n675,
                           Z => n3736);
   U489 : MUX2_X1 port map( A => registers_9_16_port, B => d_in(16), S => n675,
                           Z => n3735);
   U490 : MUX2_X1 port map( A => registers_9_15_port, B => d_in(15), S => n675,
                           Z => n3734);
   U491 : MUX2_X1 port map( A => registers_9_14_port, B => d_in(14), S => n675,
                           Z => n3733);
   U492 : MUX2_X1 port map( A => registers_9_13_port, B => d_in(13), S => n675,
                           Z => n3732);
   U493 : MUX2_X1 port map( A => registers_9_12_port, B => d_in(12), S => n675,
                           Z => n3731);
   U494 : MUX2_X1 port map( A => registers_9_11_port, B => d_in(11), S => n675,
                           Z => n3730);
   U495 : MUX2_X1 port map( A => registers_9_10_port, B => d_in(10), S => n675,
                           Z => n3729);
   U496 : MUX2_X1 port map( A => registers_9_9_port, B => d_in(9), S => n675, Z
                           => n3728);
   U497 : MUX2_X1 port map( A => registers_9_8_port, B => d_in(8), S => n675, Z
                           => n3727);
   U498 : MUX2_X1 port map( A => registers_9_7_port, B => d_in(7), S => n675, Z
                           => n3726);
   U499 : MUX2_X1 port map( A => registers_9_6_port, B => d_in(6), S => n675, Z
                           => n3725);
   U500 : MUX2_X1 port map( A => registers_9_5_port, B => d_in(5), S => n675, Z
                           => n3724);
   U501 : MUX2_X1 port map( A => registers_9_4_port, B => d_in(4), S => n675, Z
                           => n3723);
   U502 : MUX2_X1 port map( A => registers_9_3_port, B => d_in(3), S => n675, Z
                           => n3722);
   U503 : MUX2_X1 port map( A => registers_9_2_port, B => d_in(2), S => n675, Z
                           => n3721);
   U504 : MUX2_X1 port map( A => registers_9_1_port, B => d_in(1), S => n675, Z
                           => n3720);
   U505 : MUX2_X1 port map( A => registers_9_0_port, B => d_in(0), S => n675, Z
                           => n3719);
   U506 : MUX2_X1 port map( A => registers_10_31_port, B => d_in(31), S => n676
                           , Z => n3718);
   U507 : MUX2_X1 port map( A => registers_10_30_port, B => d_in(30), S => n676
                           , Z => n3717);
   U508 : MUX2_X1 port map( A => registers_10_29_port, B => d_in(29), S => n676
                           , Z => n3716);
   U509 : MUX2_X1 port map( A => registers_10_28_port, B => d_in(28), S => n676
                           , Z => n3715);
   U510 : MUX2_X1 port map( A => registers_10_27_port, B => d_in(27), S => n676
                           , Z => n3714);
   U511 : MUX2_X1 port map( A => registers_10_26_port, B => d_in(26), S => n676
                           , Z => n3713);
   U512 : MUX2_X1 port map( A => registers_10_25_port, B => d_in(25), S => n676
                           , Z => n3712);
   U513 : MUX2_X1 port map( A => registers_10_24_port, B => d_in(24), S => n676
                           , Z => n3711);
   U514 : MUX2_X1 port map( A => registers_10_23_port, B => d_in(23), S => n676
                           , Z => n3710);
   U515 : MUX2_X1 port map( A => registers_10_22_port, B => d_in(22), S => n676
                           , Z => n3709);
   U516 : MUX2_X1 port map( A => registers_10_21_port, B => d_in(21), S => n676
                           , Z => n3708);
   U517 : MUX2_X1 port map( A => registers_10_20_port, B => d_in(20), S => n676
                           , Z => n3707);
   U518 : MUX2_X1 port map( A => registers_10_19_port, B => d_in(19), S => n676
                           , Z => n3706);
   U519 : MUX2_X1 port map( A => registers_10_18_port, B => d_in(18), S => n676
                           , Z => n3705);
   U520 : MUX2_X1 port map( A => registers_10_17_port, B => d_in(17), S => n676
                           , Z => n3704);
   U521 : MUX2_X1 port map( A => registers_10_16_port, B => d_in(16), S => n676
                           , Z => n3703);
   U522 : MUX2_X1 port map( A => registers_10_15_port, B => d_in(15), S => n676
                           , Z => n3702);
   U523 : MUX2_X1 port map( A => registers_10_14_port, B => d_in(14), S => n676
                           , Z => n3701);
   U524 : MUX2_X1 port map( A => registers_10_13_port, B => d_in(13), S => n676
                           , Z => n3700);
   U525 : MUX2_X1 port map( A => registers_10_12_port, B => d_in(12), S => n676
                           , Z => n3699);
   U526 : MUX2_X1 port map( A => registers_10_11_port, B => d_in(11), S => n676
                           , Z => n3698);
   U527 : MUX2_X1 port map( A => registers_10_10_port, B => d_in(10), S => n676
                           , Z => n3697);
   U528 : MUX2_X1 port map( A => registers_10_9_port, B => d_in(9), S => n676, 
                           Z => n3696);
   U529 : MUX2_X1 port map( A => registers_10_8_port, B => d_in(8), S => n676, 
                           Z => n3695);
   U530 : MUX2_X1 port map( A => registers_10_7_port, B => d_in(7), S => n676, 
                           Z => n3694);
   U531 : MUX2_X1 port map( A => registers_10_6_port, B => d_in(6), S => n676, 
                           Z => n3693);
   U532 : MUX2_X1 port map( A => registers_10_5_port, B => d_in(5), S => n676, 
                           Z => n3692);
   U533 : MUX2_X1 port map( A => registers_10_4_port, B => d_in(4), S => n676, 
                           Z => n3691);
   U534 : MUX2_X1 port map( A => registers_10_3_port, B => d_in(3), S => n676, 
                           Z => n3690);
   U535 : MUX2_X1 port map( A => registers_10_2_port, B => d_in(2), S => n676, 
                           Z => n3689);
   U536 : MUX2_X1 port map( A => registers_10_1_port, B => d_in(1), S => n676, 
                           Z => n3688);
   U537 : MUX2_X1 port map( A => registers_10_0_port, B => d_in(0), S => n676, 
                           Z => n3687);
   U538 : MUX2_X1 port map( A => registers_11_31_port, B => d_in(31), S => n677
                           , Z => n3686);
   U539 : MUX2_X1 port map( A => registers_11_30_port, B => d_in(30), S => n677
                           , Z => n3685);
   U540 : MUX2_X1 port map( A => registers_11_29_port, B => d_in(29), S => n677
                           , Z => n3684);
   U541 : MUX2_X1 port map( A => registers_11_28_port, B => d_in(28), S => n677
                           , Z => n3683);
   U542 : MUX2_X1 port map( A => registers_11_27_port, B => d_in(27), S => n677
                           , Z => n3682);
   U543 : MUX2_X1 port map( A => registers_11_26_port, B => d_in(26), S => n677
                           , Z => n3681);
   U544 : MUX2_X1 port map( A => registers_11_25_port, B => d_in(25), S => n677
                           , Z => n3680);
   U545 : MUX2_X1 port map( A => registers_11_24_port, B => d_in(24), S => n677
                           , Z => n3679);
   U546 : MUX2_X1 port map( A => registers_11_23_port, B => d_in(23), S => n677
                           , Z => n3678);
   U547 : MUX2_X1 port map( A => registers_11_22_port, B => d_in(22), S => n677
                           , Z => n3677);
   U548 : MUX2_X1 port map( A => registers_11_21_port, B => d_in(21), S => n677
                           , Z => n3676);
   U549 : MUX2_X1 port map( A => registers_11_20_port, B => d_in(20), S => n677
                           , Z => n3675);
   U550 : MUX2_X1 port map( A => registers_11_19_port, B => d_in(19), S => n677
                           , Z => n3674);
   U551 : MUX2_X1 port map( A => registers_11_18_port, B => d_in(18), S => n677
                           , Z => n3673);
   U552 : MUX2_X1 port map( A => registers_11_17_port, B => d_in(17), S => n677
                           , Z => n3672);
   U553 : MUX2_X1 port map( A => registers_11_16_port, B => d_in(16), S => n677
                           , Z => n3671);
   U554 : MUX2_X1 port map( A => registers_11_15_port, B => d_in(15), S => n677
                           , Z => n3670);
   U555 : MUX2_X1 port map( A => registers_11_14_port, B => d_in(14), S => n677
                           , Z => n3669);
   U556 : MUX2_X1 port map( A => registers_11_13_port, B => d_in(13), S => n677
                           , Z => n3668);
   U557 : MUX2_X1 port map( A => registers_11_12_port, B => d_in(12), S => n677
                           , Z => n3667);
   U558 : MUX2_X1 port map( A => registers_11_11_port, B => d_in(11), S => n677
                           , Z => n3666);
   U559 : MUX2_X1 port map( A => registers_11_10_port, B => d_in(10), S => n677
                           , Z => n3665);
   U560 : MUX2_X1 port map( A => registers_11_9_port, B => d_in(9), S => n677, 
                           Z => n3664);
   U561 : MUX2_X1 port map( A => registers_11_8_port, B => d_in(8), S => n677, 
                           Z => n3663);
   U562 : MUX2_X1 port map( A => registers_11_7_port, B => d_in(7), S => n677, 
                           Z => n3662);
   U563 : MUX2_X1 port map( A => registers_11_6_port, B => d_in(6), S => n677, 
                           Z => n3661);
   U564 : MUX2_X1 port map( A => registers_11_5_port, B => d_in(5), S => n677, 
                           Z => n3660);
   U565 : MUX2_X1 port map( A => registers_11_4_port, B => d_in(4), S => n677, 
                           Z => n3659);
   U566 : MUX2_X1 port map( A => registers_11_3_port, B => d_in(3), S => n677, 
                           Z => n3658);
   U567 : MUX2_X1 port map( A => registers_11_2_port, B => d_in(2), S => n677, 
                           Z => n3657);
   U568 : MUX2_X1 port map( A => registers_11_1_port, B => d_in(1), S => n677, 
                           Z => n3656);
   U569 : MUX2_X1 port map( A => registers_11_0_port, B => d_in(0), S => n677, 
                           Z => n3655);
   U570 : AND3_X1 port map( A1 => n666, A2 => n664, A3 => wr_addr(3), ZN => 
                           n674);
   U571 : MUX2_X1 port map( A => registers_12_31_port, B => d_in(31), S => n678
                           , Z => n3654);
   U572 : MUX2_X1 port map( A => registers_12_30_port, B => d_in(30), S => n678
                           , Z => n3653);
   U573 : MUX2_X1 port map( A => registers_12_29_port, B => d_in(29), S => n678
                           , Z => n3652);
   U574 : MUX2_X1 port map( A => registers_12_28_port, B => d_in(28), S => n678
                           , Z => n3651);
   U575 : MUX2_X1 port map( A => registers_12_27_port, B => d_in(27), S => n678
                           , Z => n3650);
   U576 : MUX2_X1 port map( A => registers_12_26_port, B => d_in(26), S => n678
                           , Z => n3649);
   U577 : MUX2_X1 port map( A => registers_12_25_port, B => d_in(25), S => n678
                           , Z => n3648);
   U578 : MUX2_X1 port map( A => registers_12_24_port, B => d_in(24), S => n678
                           , Z => n3647);
   U579 : MUX2_X1 port map( A => registers_12_23_port, B => d_in(23), S => n678
                           , Z => n3646);
   U580 : MUX2_X1 port map( A => registers_12_22_port, B => d_in(22), S => n678
                           , Z => n3645);
   U581 : MUX2_X1 port map( A => registers_12_21_port, B => d_in(21), S => n678
                           , Z => n3644);
   U582 : MUX2_X1 port map( A => registers_12_20_port, B => d_in(20), S => n678
                           , Z => n3643);
   U583 : MUX2_X1 port map( A => registers_12_19_port, B => d_in(19), S => n678
                           , Z => n3642);
   U584 : MUX2_X1 port map( A => registers_12_18_port, B => d_in(18), S => n678
                           , Z => n3641);
   U585 : MUX2_X1 port map( A => registers_12_17_port, B => d_in(17), S => n678
                           , Z => n3640);
   U586 : MUX2_X1 port map( A => registers_12_16_port, B => d_in(16), S => n678
                           , Z => n3639);
   U587 : MUX2_X1 port map( A => registers_12_15_port, B => d_in(15), S => n678
                           , Z => n3638);
   U588 : MUX2_X1 port map( A => registers_12_14_port, B => d_in(14), S => n678
                           , Z => n3637);
   U589 : MUX2_X1 port map( A => registers_12_13_port, B => d_in(13), S => n678
                           , Z => n3636);
   U590 : MUX2_X1 port map( A => registers_12_12_port, B => d_in(12), S => n678
                           , Z => n3635);
   U591 : MUX2_X1 port map( A => registers_12_11_port, B => d_in(11), S => n678
                           , Z => n3634);
   U592 : MUX2_X1 port map( A => registers_12_10_port, B => d_in(10), S => n678
                           , Z => n3633);
   U593 : MUX2_X1 port map( A => registers_12_9_port, B => d_in(9), S => n678, 
                           Z => n3632);
   U594 : MUX2_X1 port map( A => registers_12_8_port, B => d_in(8), S => n678, 
                           Z => n3631);
   U595 : MUX2_X1 port map( A => registers_12_7_port, B => d_in(7), S => n678, 
                           Z => n3630);
   U596 : MUX2_X1 port map( A => registers_12_6_port, B => d_in(6), S => n678, 
                           Z => n3629);
   U597 : MUX2_X1 port map( A => registers_12_5_port, B => d_in(5), S => n678, 
                           Z => n3628);
   U598 : MUX2_X1 port map( A => registers_12_4_port, B => d_in(4), S => n678, 
                           Z => n3627);
   U599 : MUX2_X1 port map( A => registers_12_3_port, B => d_in(3), S => n678, 
                           Z => n3626);
   U600 : MUX2_X1 port map( A => registers_12_2_port, B => d_in(2), S => n678, 
                           Z => n3625);
   U601 : MUX2_X1 port map( A => registers_12_1_port, B => d_in(1), S => n678, 
                           Z => n3624);
   U602 : MUX2_X1 port map( A => registers_12_0_port, B => d_in(0), S => n678, 
                           Z => n3623);
   U603 : MUX2_X1 port map( A => registers_13_31_port, B => d_in(31), S => n680
                           , Z => n3622);
   U604 : MUX2_X1 port map( A => registers_13_30_port, B => d_in(30), S => n680
                           , Z => n3621);
   U605 : MUX2_X1 port map( A => registers_13_29_port, B => d_in(29), S => n680
                           , Z => n3620);
   U606 : MUX2_X1 port map( A => registers_13_28_port, B => d_in(28), S => n680
                           , Z => n3619);
   U607 : MUX2_X1 port map( A => registers_13_27_port, B => d_in(27), S => n680
                           , Z => n3618);
   U608 : MUX2_X1 port map( A => registers_13_26_port, B => d_in(26), S => n680
                           , Z => n3617);
   U609 : MUX2_X1 port map( A => registers_13_25_port, B => d_in(25), S => n680
                           , Z => n3616);
   U610 : MUX2_X1 port map( A => registers_13_24_port, B => d_in(24), S => n680
                           , Z => n3615);
   U611 : MUX2_X1 port map( A => registers_13_23_port, B => d_in(23), S => n680
                           , Z => n3614);
   U612 : MUX2_X1 port map( A => registers_13_22_port, B => d_in(22), S => n680
                           , Z => n3613);
   U613 : MUX2_X1 port map( A => registers_13_21_port, B => d_in(21), S => n680
                           , Z => n3612);
   U614 : MUX2_X1 port map( A => registers_13_20_port, B => d_in(20), S => n680
                           , Z => n3611);
   U615 : MUX2_X1 port map( A => registers_13_19_port, B => d_in(19), S => n680
                           , Z => n3610);
   U616 : MUX2_X1 port map( A => registers_13_18_port, B => d_in(18), S => n680
                           , Z => n3609);
   U617 : MUX2_X1 port map( A => registers_13_17_port, B => d_in(17), S => n680
                           , Z => n3608);
   U618 : MUX2_X1 port map( A => registers_13_16_port, B => d_in(16), S => n680
                           , Z => n3607);
   U619 : MUX2_X1 port map( A => registers_13_15_port, B => d_in(15), S => n680
                           , Z => n3606);
   U620 : MUX2_X1 port map( A => registers_13_14_port, B => d_in(14), S => n680
                           , Z => n3605);
   U621 : MUX2_X1 port map( A => registers_13_13_port, B => d_in(13), S => n680
                           , Z => n3604);
   U622 : MUX2_X1 port map( A => registers_13_12_port, B => d_in(12), S => n680
                           , Z => n3603);
   U623 : MUX2_X1 port map( A => registers_13_11_port, B => d_in(11), S => n680
                           , Z => n3602);
   U624 : MUX2_X1 port map( A => registers_13_10_port, B => d_in(10), S => n680
                           , Z => n3601);
   U625 : MUX2_X1 port map( A => registers_13_9_port, B => d_in(9), S => n680, 
                           Z => n3600);
   U626 : MUX2_X1 port map( A => registers_13_8_port, B => d_in(8), S => n680, 
                           Z => n3599);
   U627 : MUX2_X1 port map( A => registers_13_7_port, B => d_in(7), S => n680, 
                           Z => n3598);
   U628 : MUX2_X1 port map( A => registers_13_6_port, B => d_in(6), S => n680, 
                           Z => n3597);
   U629 : MUX2_X1 port map( A => registers_13_5_port, B => d_in(5), S => n680, 
                           Z => n3596);
   U630 : MUX2_X1 port map( A => registers_13_4_port, B => d_in(4), S => n680, 
                           Z => n3595);
   U631 : MUX2_X1 port map( A => registers_13_3_port, B => d_in(3), S => n680, 
                           Z => n3594);
   U632 : MUX2_X1 port map( A => registers_13_2_port, B => d_in(2), S => n680, 
                           Z => n3593);
   U633 : MUX2_X1 port map( A => registers_13_1_port, B => d_in(1), S => n680, 
                           Z => n3592);
   U634 : MUX2_X1 port map( A => registers_13_0_port, B => d_in(0), S => n680, 
                           Z => n3591);
   U635 : MUX2_X1 port map( A => registers_14_31_port, B => d_in(31), S => n681
                           , Z => n3590);
   U636 : MUX2_X1 port map( A => registers_14_30_port, B => d_in(30), S => n681
                           , Z => n3589);
   U637 : MUX2_X1 port map( A => registers_14_29_port, B => d_in(29), S => n681
                           , Z => n3588);
   U638 : MUX2_X1 port map( A => registers_14_28_port, B => d_in(28), S => n681
                           , Z => n3587);
   U639 : MUX2_X1 port map( A => registers_14_27_port, B => d_in(27), S => n681
                           , Z => n3586);
   U640 : MUX2_X1 port map( A => registers_14_26_port, B => d_in(26), S => n681
                           , Z => n3585);
   U641 : MUX2_X1 port map( A => registers_14_25_port, B => d_in(25), S => n681
                           , Z => n3584);
   U642 : MUX2_X1 port map( A => registers_14_24_port, B => d_in(24), S => n681
                           , Z => n3583);
   U643 : MUX2_X1 port map( A => registers_14_23_port, B => d_in(23), S => n681
                           , Z => n3582);
   U644 : MUX2_X1 port map( A => registers_14_22_port, B => d_in(22), S => n681
                           , Z => n3581);
   U645 : MUX2_X1 port map( A => registers_14_21_port, B => d_in(21), S => n681
                           , Z => n3580);
   U646 : MUX2_X1 port map( A => registers_14_20_port, B => d_in(20), S => n681
                           , Z => n3579);
   U647 : MUX2_X1 port map( A => registers_14_19_port, B => d_in(19), S => n681
                           , Z => n3578);
   U648 : MUX2_X1 port map( A => registers_14_18_port, B => d_in(18), S => n681
                           , Z => n3577);
   U649 : MUX2_X1 port map( A => registers_14_17_port, B => d_in(17), S => n681
                           , Z => n3576);
   U650 : MUX2_X1 port map( A => registers_14_16_port, B => d_in(16), S => n681
                           , Z => n3575);
   U651 : MUX2_X1 port map( A => registers_14_15_port, B => d_in(15), S => n681
                           , Z => n3574);
   U652 : MUX2_X1 port map( A => registers_14_14_port, B => d_in(14), S => n681
                           , Z => n3573);
   U653 : MUX2_X1 port map( A => registers_14_13_port, B => d_in(13), S => n681
                           , Z => n3572);
   U654 : MUX2_X1 port map( A => registers_14_12_port, B => d_in(12), S => n681
                           , Z => n3571);
   U655 : MUX2_X1 port map( A => registers_14_11_port, B => d_in(11), S => n681
                           , Z => n3570);
   U656 : MUX2_X1 port map( A => registers_14_10_port, B => d_in(10), S => n681
                           , Z => n3569);
   U657 : MUX2_X1 port map( A => registers_14_9_port, B => d_in(9), S => n681, 
                           Z => n3568);
   U658 : MUX2_X1 port map( A => registers_14_8_port, B => d_in(8), S => n681, 
                           Z => n3567);
   U659 : MUX2_X1 port map( A => registers_14_7_port, B => d_in(7), S => n681, 
                           Z => n3566);
   U660 : MUX2_X1 port map( A => registers_14_6_port, B => d_in(6), S => n681, 
                           Z => n3565);
   U661 : MUX2_X1 port map( A => registers_14_5_port, B => d_in(5), S => n681, 
                           Z => n3564);
   U662 : MUX2_X1 port map( A => registers_14_4_port, B => d_in(4), S => n681, 
                           Z => n3563);
   U663 : MUX2_X1 port map( A => registers_14_3_port, B => d_in(3), S => n681, 
                           Z => n3562);
   U664 : MUX2_X1 port map( A => registers_14_2_port, B => d_in(2), S => n681, 
                           Z => n3561);
   U665 : MUX2_X1 port map( A => registers_14_1_port, B => d_in(1), S => n681, 
                           Z => n3560);
   U666 : MUX2_X1 port map( A => registers_14_0_port, B => d_in(0), S => n681, 
                           Z => n3559);
   U667 : MUX2_X1 port map( A => registers_15_31_port, B => d_in(31), S => n682
                           , Z => n3558);
   U668 : MUX2_X1 port map( A => registers_15_30_port, B => d_in(30), S => n682
                           , Z => n3557);
   U669 : MUX2_X1 port map( A => registers_15_29_port, B => d_in(29), S => n682
                           , Z => n3556);
   U670 : MUX2_X1 port map( A => registers_15_28_port, B => d_in(28), S => n682
                           , Z => n3555);
   U671 : MUX2_X1 port map( A => registers_15_27_port, B => d_in(27), S => n682
                           , Z => n3554);
   U672 : MUX2_X1 port map( A => registers_15_26_port, B => d_in(26), S => n682
                           , Z => n3553);
   U673 : MUX2_X1 port map( A => registers_15_25_port, B => d_in(25), S => n682
                           , Z => n3552);
   U674 : MUX2_X1 port map( A => registers_15_24_port, B => d_in(24), S => n682
                           , Z => n3551);
   U675 : MUX2_X1 port map( A => registers_15_23_port, B => d_in(23), S => n682
                           , Z => n3550);
   U676 : MUX2_X1 port map( A => registers_15_22_port, B => d_in(22), S => n682
                           , Z => n3549);
   U677 : MUX2_X1 port map( A => registers_15_21_port, B => d_in(21), S => n682
                           , Z => n3548);
   U678 : MUX2_X1 port map( A => registers_15_20_port, B => d_in(20), S => n682
                           , Z => n3547);
   U679 : MUX2_X1 port map( A => registers_15_19_port, B => d_in(19), S => n682
                           , Z => n3546);
   U680 : MUX2_X1 port map( A => registers_15_18_port, B => d_in(18), S => n682
                           , Z => n3545);
   U681 : MUX2_X1 port map( A => registers_15_17_port, B => d_in(17), S => n682
                           , Z => n3544);
   U682 : MUX2_X1 port map( A => registers_15_16_port, B => d_in(16), S => n682
                           , Z => n3543);
   U683 : MUX2_X1 port map( A => registers_15_15_port, B => d_in(15), S => n682
                           , Z => n3542);
   U684 : MUX2_X1 port map( A => registers_15_14_port, B => d_in(14), S => n682
                           , Z => n3541);
   U685 : MUX2_X1 port map( A => registers_15_13_port, B => d_in(13), S => n682
                           , Z => n3540);
   U686 : MUX2_X1 port map( A => registers_15_12_port, B => d_in(12), S => n682
                           , Z => n3539);
   U687 : MUX2_X1 port map( A => registers_15_11_port, B => d_in(11), S => n682
                           , Z => n3538);
   U688 : MUX2_X1 port map( A => registers_15_10_port, B => d_in(10), S => n682
                           , Z => n3537);
   U689 : MUX2_X1 port map( A => registers_15_9_port, B => d_in(9), S => n682, 
                           Z => n3536);
   U690 : MUX2_X1 port map( A => registers_15_8_port, B => d_in(8), S => n682, 
                           Z => n3535);
   U691 : MUX2_X1 port map( A => registers_15_7_port, B => d_in(7), S => n682, 
                           Z => n3534);
   U692 : MUX2_X1 port map( A => registers_15_6_port, B => d_in(6), S => n682, 
                           Z => n3533);
   U693 : MUX2_X1 port map( A => registers_15_5_port, B => d_in(5), S => n682, 
                           Z => n3532);
   U694 : MUX2_X1 port map( A => registers_15_4_port, B => d_in(4), S => n682, 
                           Z => n3531);
   U695 : MUX2_X1 port map( A => registers_15_3_port, B => d_in(3), S => n682, 
                           Z => n3530);
   U696 : MUX2_X1 port map( A => registers_15_2_port, B => d_in(2), S => n682, 
                           Z => n3529);
   U697 : MUX2_X1 port map( A => registers_15_1_port, B => d_in(1), S => n682, 
                           Z => n3528);
   U698 : MUX2_X1 port map( A => registers_15_0_port, B => d_in(0), S => n682, 
                           Z => n3527);
   U699 : AND3_X1 port map( A1 => wr_addr(2), A2 => n666, A3 => wr_addr(3), ZN 
                           => n679);
   U700 : NOR3_X1 port map( A1 => n683, A2 => wr_addr(4), A3 => n684, ZN => 
                           n666);
   U701 : INV_X1 port map( A => en, ZN => n683);
   U702 : MUX2_X1 port map( A => registers_16_31_port, B => d_in(31), S => n685
                           , Z => n3526);
   U703 : MUX2_X1 port map( A => registers_16_30_port, B => d_in(30), S => n685
                           , Z => n3525);
   U704 : MUX2_X1 port map( A => registers_16_29_port, B => d_in(29), S => n685
                           , Z => n3524);
   U705 : MUX2_X1 port map( A => registers_16_28_port, B => d_in(28), S => n685
                           , Z => n3523);
   U706 : MUX2_X1 port map( A => registers_16_27_port, B => d_in(27), S => n685
                           , Z => n3522);
   U707 : MUX2_X1 port map( A => registers_16_26_port, B => d_in(26), S => n685
                           , Z => n3521);
   U708 : MUX2_X1 port map( A => registers_16_25_port, B => d_in(25), S => n685
                           , Z => n3520);
   U709 : MUX2_X1 port map( A => registers_16_24_port, B => d_in(24), S => n685
                           , Z => n3519);
   U710 : MUX2_X1 port map( A => registers_16_23_port, B => d_in(23), S => n685
                           , Z => n3518);
   U711 : MUX2_X1 port map( A => registers_16_22_port, B => d_in(22), S => n685
                           , Z => n3517);
   U712 : MUX2_X1 port map( A => registers_16_21_port, B => d_in(21), S => n685
                           , Z => n3516);
   U713 : MUX2_X1 port map( A => registers_16_20_port, B => d_in(20), S => n685
                           , Z => n3515);
   U714 : MUX2_X1 port map( A => registers_16_19_port, B => d_in(19), S => n685
                           , Z => n3514);
   U715 : MUX2_X1 port map( A => registers_16_18_port, B => d_in(18), S => n685
                           , Z => n3513);
   U716 : MUX2_X1 port map( A => registers_16_17_port, B => d_in(17), S => n685
                           , Z => n3512);
   U717 : MUX2_X1 port map( A => registers_16_16_port, B => d_in(16), S => n685
                           , Z => n3511);
   U718 : MUX2_X1 port map( A => registers_16_15_port, B => d_in(15), S => n685
                           , Z => n3510);
   U719 : MUX2_X1 port map( A => registers_16_14_port, B => d_in(14), S => n685
                           , Z => n3509);
   U720 : MUX2_X1 port map( A => registers_16_13_port, B => d_in(13), S => n685
                           , Z => n3508);
   U721 : MUX2_X1 port map( A => registers_16_12_port, B => d_in(12), S => n685
                           , Z => n3507);
   U722 : MUX2_X1 port map( A => registers_16_11_port, B => d_in(11), S => n685
                           , Z => n3506);
   U723 : MUX2_X1 port map( A => registers_16_10_port, B => d_in(10), S => n685
                           , Z => n3505);
   U724 : MUX2_X1 port map( A => registers_16_9_port, B => d_in(9), S => n685, 
                           Z => n3504);
   U725 : MUX2_X1 port map( A => registers_16_8_port, B => d_in(8), S => n685, 
                           Z => n3503);
   U726 : MUX2_X1 port map( A => registers_16_7_port, B => d_in(7), S => n685, 
                           Z => n3502);
   U727 : MUX2_X1 port map( A => registers_16_6_port, B => d_in(6), S => n685, 
                           Z => n3501);
   U728 : MUX2_X1 port map( A => registers_16_5_port, B => d_in(5), S => n685, 
                           Z => n3500);
   U729 : MUX2_X1 port map( A => registers_16_4_port, B => d_in(4), S => n685, 
                           Z => n3499);
   U730 : MUX2_X1 port map( A => registers_16_3_port, B => d_in(3), S => n685, 
                           Z => n3498);
   U731 : MUX2_X1 port map( A => registers_16_2_port, B => d_in(2), S => n685, 
                           Z => n3497);
   U732 : MUX2_X1 port map( A => registers_16_1_port, B => d_in(1), S => n685, 
                           Z => n3496);
   U733 : MUX2_X1 port map( A => registers_16_0_port, B => d_in(0), S => n685, 
                           Z => n3495);
   U734 : MUX2_X1 port map( A => registers_17_31_port, B => d_in(31), S => n687
                           , Z => n3494);
   U735 : MUX2_X1 port map( A => registers_17_30_port, B => d_in(30), S => n687
                           , Z => n3493);
   U736 : MUX2_X1 port map( A => registers_17_29_port, B => d_in(29), S => n687
                           , Z => n3492);
   U737 : MUX2_X1 port map( A => registers_17_28_port, B => d_in(28), S => n687
                           , Z => n3491);
   U738 : MUX2_X1 port map( A => registers_17_27_port, B => d_in(27), S => n687
                           , Z => n3490);
   U739 : MUX2_X1 port map( A => registers_17_26_port, B => d_in(26), S => n687
                           , Z => n3489);
   U740 : MUX2_X1 port map( A => registers_17_25_port, B => d_in(25), S => n687
                           , Z => n3488);
   U741 : MUX2_X1 port map( A => registers_17_24_port, B => d_in(24), S => n687
                           , Z => n3487);
   U742 : MUX2_X1 port map( A => registers_17_23_port, B => d_in(23), S => n687
                           , Z => n3486);
   U743 : MUX2_X1 port map( A => registers_17_22_port, B => d_in(22), S => n687
                           , Z => n3485);
   U744 : MUX2_X1 port map( A => registers_17_21_port, B => d_in(21), S => n687
                           , Z => n3484);
   U745 : MUX2_X1 port map( A => registers_17_20_port, B => d_in(20), S => n687
                           , Z => n3483);
   U746 : MUX2_X1 port map( A => registers_17_19_port, B => d_in(19), S => n687
                           , Z => n3482);
   U747 : MUX2_X1 port map( A => registers_17_18_port, B => d_in(18), S => n687
                           , Z => n3481);
   U748 : MUX2_X1 port map( A => registers_17_17_port, B => d_in(17), S => n687
                           , Z => n3480);
   U749 : MUX2_X1 port map( A => registers_17_16_port, B => d_in(16), S => n687
                           , Z => n3479);
   U750 : MUX2_X1 port map( A => registers_17_15_port, B => d_in(15), S => n687
                           , Z => n3478);
   U751 : MUX2_X1 port map( A => registers_17_14_port, B => d_in(14), S => n687
                           , Z => n3477);
   U752 : MUX2_X1 port map( A => registers_17_13_port, B => d_in(13), S => n687
                           , Z => n3476);
   U753 : MUX2_X1 port map( A => registers_17_12_port, B => d_in(12), S => n687
                           , Z => n3475);
   U754 : MUX2_X1 port map( A => registers_17_11_port, B => d_in(11), S => n687
                           , Z => n3474);
   U755 : MUX2_X1 port map( A => registers_17_10_port, B => d_in(10), S => n687
                           , Z => n3473);
   U756 : MUX2_X1 port map( A => registers_17_9_port, B => d_in(9), S => n687, 
                           Z => n3472);
   U757 : MUX2_X1 port map( A => registers_17_8_port, B => d_in(8), S => n687, 
                           Z => n3471);
   U758 : MUX2_X1 port map( A => registers_17_7_port, B => d_in(7), S => n687, 
                           Z => n3470);
   U759 : MUX2_X1 port map( A => registers_17_6_port, B => d_in(6), S => n687, 
                           Z => n3469);
   U760 : MUX2_X1 port map( A => registers_17_5_port, B => d_in(5), S => n687, 
                           Z => n3468);
   U761 : MUX2_X1 port map( A => registers_17_4_port, B => d_in(4), S => n687, 
                           Z => n3467);
   U762 : MUX2_X1 port map( A => registers_17_3_port, B => d_in(3), S => n687, 
                           Z => n3466);
   U763 : MUX2_X1 port map( A => registers_17_2_port, B => d_in(2), S => n687, 
                           Z => n3465);
   U764 : MUX2_X1 port map( A => registers_17_1_port, B => d_in(1), S => n687, 
                           Z => n3464);
   U765 : MUX2_X1 port map( A => registers_17_0_port, B => d_in(0), S => n687, 
                           Z => n3463);
   U766 : MUX2_X1 port map( A => registers_18_31_port, B => d_in(31), S => n688
                           , Z => n3462);
   U767 : MUX2_X1 port map( A => registers_18_30_port, B => d_in(30), S => n688
                           , Z => n3461);
   U768 : MUX2_X1 port map( A => registers_18_29_port, B => d_in(29), S => n688
                           , Z => n3460);
   U769 : MUX2_X1 port map( A => registers_18_28_port, B => d_in(28), S => n688
                           , Z => n3459);
   U770 : MUX2_X1 port map( A => registers_18_27_port, B => d_in(27), S => n688
                           , Z => n3458);
   U771 : MUX2_X1 port map( A => registers_18_26_port, B => d_in(26), S => n688
                           , Z => n3457);
   U772 : MUX2_X1 port map( A => registers_18_25_port, B => d_in(25), S => n688
                           , Z => n3456);
   U773 : MUX2_X1 port map( A => registers_18_24_port, B => d_in(24), S => n688
                           , Z => n3455);
   U774 : MUX2_X1 port map( A => registers_18_23_port, B => d_in(23), S => n688
                           , Z => n3454);
   U775 : MUX2_X1 port map( A => registers_18_22_port, B => d_in(22), S => n688
                           , Z => n3453);
   U776 : MUX2_X1 port map( A => registers_18_21_port, B => d_in(21), S => n688
                           , Z => n3452);
   U777 : MUX2_X1 port map( A => registers_18_20_port, B => d_in(20), S => n688
                           , Z => n3451);
   U778 : MUX2_X1 port map( A => registers_18_19_port, B => d_in(19), S => n688
                           , Z => n3450);
   U779 : MUX2_X1 port map( A => registers_18_18_port, B => d_in(18), S => n688
                           , Z => n3449);
   U780 : MUX2_X1 port map( A => registers_18_17_port, B => d_in(17), S => n688
                           , Z => n3448);
   U781 : MUX2_X1 port map( A => registers_18_16_port, B => d_in(16), S => n688
                           , Z => n3447);
   U782 : MUX2_X1 port map( A => registers_18_15_port, B => d_in(15), S => n688
                           , Z => n3446);
   U783 : MUX2_X1 port map( A => registers_18_14_port, B => d_in(14), S => n688
                           , Z => n3445);
   U784 : MUX2_X1 port map( A => registers_18_13_port, B => d_in(13), S => n688
                           , Z => n3444);
   U785 : MUX2_X1 port map( A => registers_18_12_port, B => d_in(12), S => n688
                           , Z => n3443);
   U786 : MUX2_X1 port map( A => registers_18_11_port, B => d_in(11), S => n688
                           , Z => n3442);
   U787 : MUX2_X1 port map( A => registers_18_10_port, B => d_in(10), S => n688
                           , Z => n3441);
   U788 : MUX2_X1 port map( A => registers_18_9_port, B => d_in(9), S => n688, 
                           Z => n3440);
   U789 : MUX2_X1 port map( A => registers_18_8_port, B => d_in(8), S => n688, 
                           Z => n3439);
   U790 : MUX2_X1 port map( A => registers_18_7_port, B => d_in(7), S => n688, 
                           Z => n3438);
   U791 : MUX2_X1 port map( A => registers_18_6_port, B => d_in(6), S => n688, 
                           Z => n3437);
   U792 : MUX2_X1 port map( A => registers_18_5_port, B => d_in(5), S => n688, 
                           Z => n3436);
   U793 : MUX2_X1 port map( A => registers_18_4_port, B => d_in(4), S => n688, 
                           Z => n3435);
   U794 : MUX2_X1 port map( A => registers_18_3_port, B => d_in(3), S => n688, 
                           Z => n3434);
   U795 : MUX2_X1 port map( A => registers_18_2_port, B => d_in(2), S => n688, 
                           Z => n3433);
   U796 : MUX2_X1 port map( A => registers_18_1_port, B => d_in(1), S => n688, 
                           Z => n3432);
   U797 : MUX2_X1 port map( A => registers_18_0_port, B => d_in(0), S => n688, 
                           Z => n3431);
   U798 : MUX2_X1 port map( A => registers_19_31_port, B => d_in(31), S => n689
                           , Z => n3430);
   U799 : MUX2_X1 port map( A => registers_19_30_port, B => d_in(30), S => n689
                           , Z => n3429);
   U800 : MUX2_X1 port map( A => registers_19_29_port, B => d_in(29), S => n689
                           , Z => n3428);
   U801 : MUX2_X1 port map( A => registers_19_28_port, B => d_in(28), S => n689
                           , Z => n3427);
   U802 : MUX2_X1 port map( A => registers_19_27_port, B => d_in(27), S => n689
                           , Z => n3426);
   U803 : MUX2_X1 port map( A => registers_19_26_port, B => d_in(26), S => n689
                           , Z => n3425);
   U804 : MUX2_X1 port map( A => registers_19_25_port, B => d_in(25), S => n689
                           , Z => n3424);
   U805 : MUX2_X1 port map( A => registers_19_24_port, B => d_in(24), S => n689
                           , Z => n3423);
   U806 : MUX2_X1 port map( A => registers_19_23_port, B => d_in(23), S => n689
                           , Z => n3422);
   U807 : MUX2_X1 port map( A => registers_19_22_port, B => d_in(22), S => n689
                           , Z => n3421);
   U808 : MUX2_X1 port map( A => registers_19_21_port, B => d_in(21), S => n689
                           , Z => n3420);
   U809 : MUX2_X1 port map( A => registers_19_20_port, B => d_in(20), S => n689
                           , Z => n3419);
   U810 : MUX2_X1 port map( A => registers_19_19_port, B => d_in(19), S => n689
                           , Z => n3418);
   U811 : MUX2_X1 port map( A => registers_19_18_port, B => d_in(18), S => n689
                           , Z => n3417);
   U812 : MUX2_X1 port map( A => registers_19_17_port, B => d_in(17), S => n689
                           , Z => n3416);
   U813 : MUX2_X1 port map( A => registers_19_16_port, B => d_in(16), S => n689
                           , Z => n3415);
   U814 : MUX2_X1 port map( A => registers_19_15_port, B => d_in(15), S => n689
                           , Z => n3414);
   U815 : MUX2_X1 port map( A => registers_19_14_port, B => d_in(14), S => n689
                           , Z => n3413);
   U816 : MUX2_X1 port map( A => registers_19_13_port, B => d_in(13), S => n689
                           , Z => n3412);
   U817 : MUX2_X1 port map( A => registers_19_12_port, B => d_in(12), S => n689
                           , Z => n3411);
   U818 : MUX2_X1 port map( A => registers_19_11_port, B => d_in(11), S => n689
                           , Z => n3410);
   U819 : MUX2_X1 port map( A => registers_19_10_port, B => d_in(10), S => n689
                           , Z => n3409);
   U820 : MUX2_X1 port map( A => registers_19_9_port, B => d_in(9), S => n689, 
                           Z => n3408);
   U821 : MUX2_X1 port map( A => registers_19_8_port, B => d_in(8), S => n689, 
                           Z => n3407);
   U822 : MUX2_X1 port map( A => registers_19_7_port, B => d_in(7), S => n689, 
                           Z => n3406);
   U823 : MUX2_X1 port map( A => registers_19_6_port, B => d_in(6), S => n689, 
                           Z => n3405);
   U824 : MUX2_X1 port map( A => registers_19_5_port, B => d_in(5), S => n689, 
                           Z => n3404);
   U825 : MUX2_X1 port map( A => registers_19_4_port, B => d_in(4), S => n689, 
                           Z => n3403);
   U826 : MUX2_X1 port map( A => registers_19_3_port, B => d_in(3), S => n689, 
                           Z => n3402);
   U827 : MUX2_X1 port map( A => registers_19_2_port, B => d_in(2), S => n689, 
                           Z => n3401);
   U828 : MUX2_X1 port map( A => registers_19_1_port, B => d_in(1), S => n689, 
                           Z => n3400);
   U829 : MUX2_X1 port map( A => registers_19_0_port, B => d_in(0), S => n689, 
                           Z => n3399);
   U830 : AND3_X1 port map( A1 => n664, A2 => n665, A3 => n690, ZN => n686);
   U831 : MUX2_X1 port map( A => registers_20_31_port, B => d_in(31), S => n691
                           , Z => n3398);
   U832 : MUX2_X1 port map( A => registers_20_30_port, B => d_in(30), S => n691
                           , Z => n3397);
   U833 : MUX2_X1 port map( A => registers_20_29_port, B => d_in(29), S => n691
                           , Z => n3396);
   U834 : MUX2_X1 port map( A => registers_20_28_port, B => d_in(28), S => n691
                           , Z => n3395);
   U835 : MUX2_X1 port map( A => registers_20_27_port, B => d_in(27), S => n691
                           , Z => n3394);
   U836 : MUX2_X1 port map( A => registers_20_26_port, B => d_in(26), S => n691
                           , Z => n3393);
   U837 : MUX2_X1 port map( A => registers_20_25_port, B => d_in(25), S => n691
                           , Z => n3392);
   U838 : MUX2_X1 port map( A => registers_20_24_port, B => d_in(24), S => n691
                           , Z => n3391);
   U839 : MUX2_X1 port map( A => registers_20_23_port, B => d_in(23), S => n691
                           , Z => n3390);
   U840 : MUX2_X1 port map( A => registers_20_22_port, B => d_in(22), S => n691
                           , Z => n3389);
   U841 : MUX2_X1 port map( A => registers_20_21_port, B => d_in(21), S => n691
                           , Z => n3388);
   U842 : MUX2_X1 port map( A => registers_20_20_port, B => d_in(20), S => n691
                           , Z => n3387);
   U843 : MUX2_X1 port map( A => registers_20_19_port, B => d_in(19), S => n691
                           , Z => n3386);
   U844 : MUX2_X1 port map( A => registers_20_18_port, B => d_in(18), S => n691
                           , Z => n3385);
   U845 : MUX2_X1 port map( A => registers_20_17_port, B => d_in(17), S => n691
                           , Z => n3384);
   U846 : MUX2_X1 port map( A => registers_20_16_port, B => d_in(16), S => n691
                           , Z => n3383);
   U847 : MUX2_X1 port map( A => registers_20_15_port, B => d_in(15), S => n691
                           , Z => n3382);
   U848 : MUX2_X1 port map( A => registers_20_14_port, B => d_in(14), S => n691
                           , Z => n3381);
   U849 : MUX2_X1 port map( A => registers_20_13_port, B => d_in(13), S => n691
                           , Z => n3380);
   U850 : MUX2_X1 port map( A => registers_20_12_port, B => d_in(12), S => n691
                           , Z => n3379);
   U851 : MUX2_X1 port map( A => registers_20_11_port, B => d_in(11), S => n691
                           , Z => n3378);
   U852 : MUX2_X1 port map( A => registers_20_10_port, B => d_in(10), S => n691
                           , Z => n3377);
   U853 : MUX2_X1 port map( A => registers_20_9_port, B => d_in(9), S => n691, 
                           Z => n3376);
   U854 : MUX2_X1 port map( A => registers_20_8_port, B => d_in(8), S => n691, 
                           Z => n3375);
   U855 : MUX2_X1 port map( A => registers_20_7_port, B => d_in(7), S => n691, 
                           Z => n3374);
   U856 : MUX2_X1 port map( A => registers_20_6_port, B => d_in(6), S => n691, 
                           Z => n3373);
   U857 : MUX2_X1 port map( A => registers_20_5_port, B => d_in(5), S => n691, 
                           Z => n3372);
   U858 : MUX2_X1 port map( A => registers_20_4_port, B => d_in(4), S => n691, 
                           Z => n3371);
   U859 : MUX2_X1 port map( A => registers_20_3_port, B => d_in(3), S => n691, 
                           Z => n3370);
   U860 : MUX2_X1 port map( A => registers_20_2_port, B => d_in(2), S => n691, 
                           Z => n3369);
   U861 : MUX2_X1 port map( A => registers_20_1_port, B => d_in(1), S => n691, 
                           Z => n3368);
   U862 : MUX2_X1 port map( A => registers_20_0_port, B => d_in(0), S => n691, 
                           Z => n3367);
   U863 : MUX2_X1 port map( A => registers_21_31_port, B => d_in(31), S => n693
                           , Z => n3366);
   U864 : MUX2_X1 port map( A => registers_21_30_port, B => d_in(30), S => n693
                           , Z => n3365);
   U865 : MUX2_X1 port map( A => registers_21_29_port, B => d_in(29), S => n693
                           , Z => n3364);
   U866 : MUX2_X1 port map( A => registers_21_28_port, B => d_in(28), S => n693
                           , Z => n3363);
   U867 : MUX2_X1 port map( A => registers_21_27_port, B => d_in(27), S => n693
                           , Z => n3362);
   U868 : MUX2_X1 port map( A => registers_21_26_port, B => d_in(26), S => n693
                           , Z => n3361);
   U869 : MUX2_X1 port map( A => registers_21_25_port, B => d_in(25), S => n693
                           , Z => n3360);
   U870 : MUX2_X1 port map( A => registers_21_24_port, B => d_in(24), S => n693
                           , Z => n3359);
   U871 : MUX2_X1 port map( A => registers_21_23_port, B => d_in(23), S => n693
                           , Z => n3358);
   U872 : MUX2_X1 port map( A => registers_21_22_port, B => d_in(22), S => n693
                           , Z => n3357);
   U873 : MUX2_X1 port map( A => registers_21_21_port, B => d_in(21), S => n693
                           , Z => n3356);
   U874 : MUX2_X1 port map( A => registers_21_20_port, B => d_in(20), S => n693
                           , Z => n3355);
   U875 : MUX2_X1 port map( A => registers_21_19_port, B => d_in(19), S => n693
                           , Z => n3354);
   U876 : MUX2_X1 port map( A => registers_21_18_port, B => d_in(18), S => n693
                           , Z => n3353);
   U877 : MUX2_X1 port map( A => registers_21_17_port, B => d_in(17), S => n693
                           , Z => n3352);
   U878 : MUX2_X1 port map( A => registers_21_16_port, B => d_in(16), S => n693
                           , Z => n3351);
   U879 : MUX2_X1 port map( A => registers_21_15_port, B => d_in(15), S => n693
                           , Z => n3350);
   U880 : MUX2_X1 port map( A => registers_21_14_port, B => d_in(14), S => n693
                           , Z => n3349);
   U881 : MUX2_X1 port map( A => registers_21_13_port, B => d_in(13), S => n693
                           , Z => n3348);
   U882 : MUX2_X1 port map( A => registers_21_12_port, B => d_in(12), S => n693
                           , Z => n3347);
   U883 : MUX2_X1 port map( A => registers_21_11_port, B => d_in(11), S => n693
                           , Z => n3346);
   U884 : MUX2_X1 port map( A => registers_21_10_port, B => d_in(10), S => n693
                           , Z => n3345);
   U885 : MUX2_X1 port map( A => registers_21_9_port, B => d_in(9), S => n693, 
                           Z => n3344);
   U886 : MUX2_X1 port map( A => registers_21_8_port, B => d_in(8), S => n693, 
                           Z => n3343);
   U887 : MUX2_X1 port map( A => registers_21_7_port, B => d_in(7), S => n693, 
                           Z => n3342);
   U888 : MUX2_X1 port map( A => registers_21_6_port, B => d_in(6), S => n693, 
                           Z => n3341);
   U889 : MUX2_X1 port map( A => registers_21_5_port, B => d_in(5), S => n693, 
                           Z => n3340);
   U890 : MUX2_X1 port map( A => registers_21_4_port, B => d_in(4), S => n693, 
                           Z => n3339);
   U891 : MUX2_X1 port map( A => registers_21_3_port, B => d_in(3), S => n693, 
                           Z => n3338);
   U892 : MUX2_X1 port map( A => registers_21_2_port, B => d_in(2), S => n693, 
                           Z => n3337);
   U893 : MUX2_X1 port map( A => registers_21_1_port, B => d_in(1), S => n693, 
                           Z => n3336);
   U894 : MUX2_X1 port map( A => registers_21_0_port, B => d_in(0), S => n693, 
                           Z => n3335);
   U895 : MUX2_X1 port map( A => registers_22_31_port, B => d_in(31), S => n694
                           , Z => n3334);
   U896 : MUX2_X1 port map( A => registers_22_30_port, B => d_in(30), S => n694
                           , Z => n3333);
   U897 : MUX2_X1 port map( A => registers_22_29_port, B => d_in(29), S => n694
                           , Z => n3332);
   U898 : MUX2_X1 port map( A => registers_22_28_port, B => d_in(28), S => n694
                           , Z => n3331);
   U899 : MUX2_X1 port map( A => registers_22_27_port, B => d_in(27), S => n694
                           , Z => n3330);
   U900 : MUX2_X1 port map( A => registers_22_26_port, B => d_in(26), S => n694
                           , Z => n3329);
   U901 : MUX2_X1 port map( A => registers_22_25_port, B => d_in(25), S => n694
                           , Z => n3328);
   U902 : MUX2_X1 port map( A => registers_22_24_port, B => d_in(24), S => n694
                           , Z => n3327);
   U903 : MUX2_X1 port map( A => registers_22_23_port, B => d_in(23), S => n694
                           , Z => n3326);
   U904 : MUX2_X1 port map( A => registers_22_22_port, B => d_in(22), S => n694
                           , Z => n3325);
   U905 : MUX2_X1 port map( A => registers_22_21_port, B => d_in(21), S => n694
                           , Z => n3324);
   U906 : MUX2_X1 port map( A => registers_22_20_port, B => d_in(20), S => n694
                           , Z => n3323);
   U907 : MUX2_X1 port map( A => registers_22_19_port, B => d_in(19), S => n694
                           , Z => n3322);
   U908 : MUX2_X1 port map( A => registers_22_18_port, B => d_in(18), S => n694
                           , Z => n3321);
   U909 : MUX2_X1 port map( A => registers_22_17_port, B => d_in(17), S => n694
                           , Z => n3320);
   U910 : MUX2_X1 port map( A => registers_22_16_port, B => d_in(16), S => n694
                           , Z => n3319);
   U911 : MUX2_X1 port map( A => registers_22_15_port, B => d_in(15), S => n694
                           , Z => n3318);
   U912 : MUX2_X1 port map( A => registers_22_14_port, B => d_in(14), S => n694
                           , Z => n3317);
   U913 : MUX2_X1 port map( A => registers_22_13_port, B => d_in(13), S => n694
                           , Z => n3316);
   U914 : MUX2_X1 port map( A => registers_22_12_port, B => d_in(12), S => n694
                           , Z => n3315);
   U915 : MUX2_X1 port map( A => registers_22_11_port, B => d_in(11), S => n694
                           , Z => n3314);
   U916 : MUX2_X1 port map( A => registers_22_10_port, B => d_in(10), S => n694
                           , Z => n3313);
   U917 : MUX2_X1 port map( A => registers_22_9_port, B => d_in(9), S => n694, 
                           Z => n3312);
   U918 : MUX2_X1 port map( A => registers_22_8_port, B => d_in(8), S => n694, 
                           Z => n3311);
   U919 : MUX2_X1 port map( A => registers_22_7_port, B => d_in(7), S => n694, 
                           Z => n3310);
   U920 : MUX2_X1 port map( A => registers_22_6_port, B => d_in(6), S => n694, 
                           Z => n3309);
   U921 : MUX2_X1 port map( A => registers_22_5_port, B => d_in(5), S => n694, 
                           Z => n3308);
   U922 : MUX2_X1 port map( A => registers_22_4_port, B => d_in(4), S => n694, 
                           Z => n3307);
   U923 : MUX2_X1 port map( A => registers_22_3_port, B => d_in(3), S => n694, 
                           Z => n3306);
   U924 : MUX2_X1 port map( A => registers_22_2_port, B => d_in(2), S => n694, 
                           Z => n3305);
   U925 : MUX2_X1 port map( A => registers_22_1_port, B => d_in(1), S => n694, 
                           Z => n3304);
   U926 : MUX2_X1 port map( A => registers_22_0_port, B => d_in(0), S => n694, 
                           Z => n3303);
   U927 : MUX2_X1 port map( A => registers_23_31_port, B => d_in(31), S => n695
                           , Z => n3302);
   U928 : MUX2_X1 port map( A => registers_23_30_port, B => d_in(30), S => n695
                           , Z => n3301);
   U929 : MUX2_X1 port map( A => registers_23_29_port, B => d_in(29), S => n695
                           , Z => n3300);
   U930 : MUX2_X1 port map( A => registers_23_28_port, B => d_in(28), S => n695
                           , Z => n3299);
   U931 : MUX2_X1 port map( A => registers_23_27_port, B => d_in(27), S => n695
                           , Z => n3298);
   U932 : MUX2_X1 port map( A => registers_23_26_port, B => d_in(26), S => n695
                           , Z => n3297);
   U933 : MUX2_X1 port map( A => registers_23_25_port, B => d_in(25), S => n695
                           , Z => n3296);
   U934 : MUX2_X1 port map( A => registers_23_24_port, B => d_in(24), S => n695
                           , Z => n3295);
   U935 : MUX2_X1 port map( A => registers_23_23_port, B => d_in(23), S => n695
                           , Z => n3294);
   U936 : MUX2_X1 port map( A => registers_23_22_port, B => d_in(22), S => n695
                           , Z => n3293);
   U937 : MUX2_X1 port map( A => registers_23_21_port, B => d_in(21), S => n695
                           , Z => n3292);
   U938 : MUX2_X1 port map( A => registers_23_20_port, B => d_in(20), S => n695
                           , Z => n3291);
   U939 : MUX2_X1 port map( A => registers_23_19_port, B => d_in(19), S => n695
                           , Z => n3290);
   U940 : MUX2_X1 port map( A => registers_23_18_port, B => d_in(18), S => n695
                           , Z => n3289);
   U941 : MUX2_X1 port map( A => registers_23_17_port, B => d_in(17), S => n695
                           , Z => n3288);
   U942 : MUX2_X1 port map( A => registers_23_16_port, B => d_in(16), S => n695
                           , Z => n3287);
   U943 : MUX2_X1 port map( A => registers_23_15_port, B => d_in(15), S => n695
                           , Z => n3286);
   U944 : MUX2_X1 port map( A => registers_23_14_port, B => d_in(14), S => n695
                           , Z => n3285);
   U945 : MUX2_X1 port map( A => registers_23_13_port, B => d_in(13), S => n695
                           , Z => n3284);
   U946 : MUX2_X1 port map( A => registers_23_12_port, B => d_in(12), S => n695
                           , Z => n3283);
   U947 : MUX2_X1 port map( A => registers_23_11_port, B => d_in(11), S => n695
                           , Z => n3282);
   U948 : MUX2_X1 port map( A => registers_23_10_port, B => d_in(10), S => n695
                           , Z => n3281);
   U949 : MUX2_X1 port map( A => registers_23_9_port, B => d_in(9), S => n695, 
                           Z => n3280);
   U950 : MUX2_X1 port map( A => registers_23_8_port, B => d_in(8), S => n695, 
                           Z => n3279);
   U951 : MUX2_X1 port map( A => registers_23_7_port, B => d_in(7), S => n695, 
                           Z => n3278);
   U952 : MUX2_X1 port map( A => registers_23_6_port, B => d_in(6), S => n695, 
                           Z => n3277);
   U953 : MUX2_X1 port map( A => registers_23_5_port, B => d_in(5), S => n695, 
                           Z => n3276);
   U954 : MUX2_X1 port map( A => registers_23_4_port, B => d_in(4), S => n695, 
                           Z => n3275);
   U955 : MUX2_X1 port map( A => registers_23_3_port, B => d_in(3), S => n695, 
                           Z => n3274);
   U956 : MUX2_X1 port map( A => registers_23_2_port, B => d_in(2), S => n695, 
                           Z => n3273);
   U957 : MUX2_X1 port map( A => registers_23_1_port, B => d_in(1), S => n695, 
                           Z => n3272);
   U958 : MUX2_X1 port map( A => registers_23_0_port, B => d_in(0), S => n695, 
                           Z => n3271);
   U959 : AND3_X1 port map( A1 => wr_addr(2), A2 => n665, A3 => n690, ZN => 
                           n692);
   U960 : INV_X1 port map( A => wr_addr(3), ZN => n665);
   U961 : MUX2_X1 port map( A => registers_24_31_port, B => d_in(31), S => n696
                           , Z => n3270);
   U962 : MUX2_X1 port map( A => registers_24_30_port, B => d_in(30), S => n696
                           , Z => n3269);
   U963 : MUX2_X1 port map( A => registers_24_29_port, B => d_in(29), S => n696
                           , Z => n3268);
   U964 : MUX2_X1 port map( A => registers_24_28_port, B => d_in(28), S => n696
                           , Z => n3267);
   U965 : MUX2_X1 port map( A => registers_24_27_port, B => d_in(27), S => n696
                           , Z => n3266);
   U966 : MUX2_X1 port map( A => registers_24_26_port, B => d_in(26), S => n696
                           , Z => n3265);
   U967 : MUX2_X1 port map( A => registers_24_25_port, B => d_in(25), S => n696
                           , Z => n3264);
   U968 : MUX2_X1 port map( A => registers_24_24_port, B => d_in(24), S => n696
                           , Z => n3263);
   U969 : MUX2_X1 port map( A => registers_24_23_port, B => d_in(23), S => n696
                           , Z => n3262);
   U970 : MUX2_X1 port map( A => registers_24_22_port, B => d_in(22), S => n696
                           , Z => n3261);
   U971 : MUX2_X1 port map( A => registers_24_21_port, B => d_in(21), S => n696
                           , Z => n3260);
   U972 : MUX2_X1 port map( A => registers_24_20_port, B => d_in(20), S => n696
                           , Z => n3259);
   U973 : MUX2_X1 port map( A => registers_24_19_port, B => d_in(19), S => n696
                           , Z => n3258);
   U974 : MUX2_X1 port map( A => registers_24_18_port, B => d_in(18), S => n696
                           , Z => n3257);
   U975 : MUX2_X1 port map( A => registers_24_17_port, B => d_in(17), S => n696
                           , Z => n3256);
   U976 : MUX2_X1 port map( A => registers_24_16_port, B => d_in(16), S => n696
                           , Z => n3255);
   U977 : MUX2_X1 port map( A => registers_24_15_port, B => d_in(15), S => n696
                           , Z => n3254);
   U978 : MUX2_X1 port map( A => registers_24_14_port, B => d_in(14), S => n696
                           , Z => n3253);
   U979 : MUX2_X1 port map( A => registers_24_13_port, B => d_in(13), S => n696
                           , Z => n3252);
   U980 : MUX2_X1 port map( A => registers_24_12_port, B => d_in(12), S => n696
                           , Z => n3251);
   U981 : MUX2_X1 port map( A => registers_24_11_port, B => d_in(11), S => n696
                           , Z => n3250);
   U982 : MUX2_X1 port map( A => registers_24_10_port, B => d_in(10), S => n696
                           , Z => n3249);
   U983 : MUX2_X1 port map( A => registers_24_9_port, B => d_in(9), S => n696, 
                           Z => n3248);
   U984 : MUX2_X1 port map( A => registers_24_8_port, B => d_in(8), S => n696, 
                           Z => n3247);
   U985 : MUX2_X1 port map( A => registers_24_7_port, B => d_in(7), S => n696, 
                           Z => n3246);
   U986 : MUX2_X1 port map( A => registers_24_6_port, B => d_in(6), S => n696, 
                           Z => n3245);
   U987 : MUX2_X1 port map( A => registers_24_5_port, B => d_in(5), S => n696, 
                           Z => n3244);
   U988 : MUX2_X1 port map( A => registers_24_4_port, B => d_in(4), S => n696, 
                           Z => n3243);
   U989 : MUX2_X1 port map( A => registers_24_3_port, B => d_in(3), S => n696, 
                           Z => n3242);
   U990 : MUX2_X1 port map( A => registers_24_2_port, B => d_in(2), S => n696, 
                           Z => n3241);
   U991 : MUX2_X1 port map( A => registers_24_1_port, B => d_in(1), S => n696, 
                           Z => n3240);
   U992 : MUX2_X1 port map( A => registers_24_0_port, B => d_in(0), S => n696, 
                           Z => n3239);
   U993 : MUX2_X1 port map( A => registers_25_31_port, B => d_in(31), S => n698
                           , Z => n3238);
   U994 : MUX2_X1 port map( A => registers_25_30_port, B => d_in(30), S => n698
                           , Z => n3237);
   U995 : MUX2_X1 port map( A => registers_25_29_port, B => d_in(29), S => n698
                           , Z => n3236);
   U996 : MUX2_X1 port map( A => registers_25_28_port, B => d_in(28), S => n698
                           , Z => n3235);
   U997 : MUX2_X1 port map( A => registers_25_27_port, B => d_in(27), S => n698
                           , Z => n3234);
   U998 : MUX2_X1 port map( A => registers_25_26_port, B => d_in(26), S => n698
                           , Z => n3233);
   U999 : MUX2_X1 port map( A => registers_25_25_port, B => d_in(25), S => n698
                           , Z => n3232);
   U1000 : MUX2_X1 port map( A => registers_25_24_port, B => d_in(24), S => 
                           n698, Z => n3231);
   U1001 : MUX2_X1 port map( A => registers_25_23_port, B => d_in(23), S => 
                           n698, Z => n3230);
   U1002 : MUX2_X1 port map( A => registers_25_22_port, B => d_in(22), S => 
                           n698, Z => n3229);
   U1003 : MUX2_X1 port map( A => registers_25_21_port, B => d_in(21), S => 
                           n698, Z => n3228);
   U1004 : MUX2_X1 port map( A => registers_25_20_port, B => d_in(20), S => 
                           n698, Z => n3227);
   U1005 : MUX2_X1 port map( A => registers_25_19_port, B => d_in(19), S => 
                           n698, Z => n3226);
   U1006 : MUX2_X1 port map( A => registers_25_18_port, B => d_in(18), S => 
                           n698, Z => n3225);
   U1007 : MUX2_X1 port map( A => registers_25_17_port, B => d_in(17), S => 
                           n698, Z => n3224);
   U1008 : MUX2_X1 port map( A => registers_25_16_port, B => d_in(16), S => 
                           n698, Z => n3223);
   U1009 : MUX2_X1 port map( A => registers_25_15_port, B => d_in(15), S => 
                           n698, Z => n3222);
   U1010 : MUX2_X1 port map( A => registers_25_14_port, B => d_in(14), S => 
                           n698, Z => n3221);
   U1011 : MUX2_X1 port map( A => registers_25_13_port, B => d_in(13), S => 
                           n698, Z => n3220);
   U1012 : MUX2_X1 port map( A => registers_25_12_port, B => d_in(12), S => 
                           n698, Z => n3219);
   U1013 : MUX2_X1 port map( A => registers_25_11_port, B => d_in(11), S => 
                           n698, Z => n3218);
   U1014 : MUX2_X1 port map( A => registers_25_10_port, B => d_in(10), S => 
                           n698, Z => n3217);
   U1015 : MUX2_X1 port map( A => registers_25_9_port, B => d_in(9), S => n698,
                           Z => n3216);
   U1016 : MUX2_X1 port map( A => registers_25_8_port, B => d_in(8), S => n698,
                           Z => n3215);
   U1017 : MUX2_X1 port map( A => registers_25_7_port, B => d_in(7), S => n698,
                           Z => n3214);
   U1018 : MUX2_X1 port map( A => registers_25_6_port, B => d_in(6), S => n698,
                           Z => n3213);
   U1019 : MUX2_X1 port map( A => registers_25_5_port, B => d_in(5), S => n698,
                           Z => n3212);
   U1020 : MUX2_X1 port map( A => registers_25_4_port, B => d_in(4), S => n698,
                           Z => n3211);
   U1021 : MUX2_X1 port map( A => registers_25_3_port, B => d_in(3), S => n698,
                           Z => n3210);
   U1022 : MUX2_X1 port map( A => registers_25_2_port, B => d_in(2), S => n698,
                           Z => n3209);
   U1023 : MUX2_X1 port map( A => registers_25_1_port, B => d_in(1), S => n698,
                           Z => n3208);
   U1024 : MUX2_X1 port map( A => registers_25_0_port, B => d_in(0), S => n698,
                           Z => n3207);
   U1025 : MUX2_X1 port map( A => registers_26_31_port, B => d_in(31), S => 
                           n699, Z => n3206);
   U1026 : MUX2_X1 port map( A => registers_26_30_port, B => d_in(30), S => 
                           n699, Z => n3205);
   U1027 : MUX2_X1 port map( A => registers_26_29_port, B => d_in(29), S => 
                           n699, Z => n3204);
   U1028 : MUX2_X1 port map( A => registers_26_28_port, B => d_in(28), S => 
                           n699, Z => n3203);
   U1029 : MUX2_X1 port map( A => registers_26_27_port, B => d_in(27), S => 
                           n699, Z => n3202);
   U1030 : MUX2_X1 port map( A => registers_26_26_port, B => d_in(26), S => 
                           n699, Z => n3201);
   U1031 : MUX2_X1 port map( A => registers_26_25_port, B => d_in(25), S => 
                           n699, Z => n3200);
   U1032 : MUX2_X1 port map( A => registers_26_24_port, B => d_in(24), S => 
                           n699, Z => n3199);
   U1033 : MUX2_X1 port map( A => registers_26_23_port, B => d_in(23), S => 
                           n699, Z => n3198);
   U1034 : MUX2_X1 port map( A => registers_26_22_port, B => d_in(22), S => 
                           n699, Z => n3197);
   U1035 : MUX2_X1 port map( A => registers_26_21_port, B => d_in(21), S => 
                           n699, Z => n3196);
   U1036 : MUX2_X1 port map( A => registers_26_20_port, B => d_in(20), S => 
                           n699, Z => n3195);
   U1037 : MUX2_X1 port map( A => registers_26_19_port, B => d_in(19), S => 
                           n699, Z => n3194);
   U1038 : MUX2_X1 port map( A => registers_26_18_port, B => d_in(18), S => 
                           n699, Z => n3193);
   U1039 : MUX2_X1 port map( A => registers_26_17_port, B => d_in(17), S => 
                           n699, Z => n3192);
   U1040 : MUX2_X1 port map( A => registers_26_16_port, B => d_in(16), S => 
                           n699, Z => n3191);
   U1041 : MUX2_X1 port map( A => registers_26_15_port, B => d_in(15), S => 
                           n699, Z => n3190);
   U1042 : MUX2_X1 port map( A => registers_26_14_port, B => d_in(14), S => 
                           n699, Z => n3189);
   U1043 : MUX2_X1 port map( A => registers_26_13_port, B => d_in(13), S => 
                           n699, Z => n3188);
   U1044 : MUX2_X1 port map( A => registers_26_12_port, B => d_in(12), S => 
                           n699, Z => n3187);
   U1045 : MUX2_X1 port map( A => registers_26_11_port, B => d_in(11), S => 
                           n699, Z => n3186);
   U1046 : MUX2_X1 port map( A => registers_26_10_port, B => d_in(10), S => 
                           n699, Z => n3185);
   U1047 : MUX2_X1 port map( A => registers_26_9_port, B => d_in(9), S => n699,
                           Z => n3184);
   U1048 : MUX2_X1 port map( A => registers_26_8_port, B => d_in(8), S => n699,
                           Z => n3183);
   U1049 : MUX2_X1 port map( A => registers_26_7_port, B => d_in(7), S => n699,
                           Z => n3182);
   U1050 : MUX2_X1 port map( A => registers_26_6_port, B => d_in(6), S => n699,
                           Z => n3181);
   U1051 : MUX2_X1 port map( A => registers_26_5_port, B => d_in(5), S => n699,
                           Z => n3180);
   U1052 : MUX2_X1 port map( A => registers_26_4_port, B => d_in(4), S => n699,
                           Z => n3179);
   U1053 : MUX2_X1 port map( A => registers_26_3_port, B => d_in(3), S => n699,
                           Z => n3178);
   U1054 : MUX2_X1 port map( A => registers_26_2_port, B => d_in(2), S => n699,
                           Z => n3177);
   U1055 : MUX2_X1 port map( A => registers_26_1_port, B => d_in(1), S => n699,
                           Z => n3176);
   U1056 : MUX2_X1 port map( A => registers_26_0_port, B => d_in(0), S => n699,
                           Z => n3175);
   U1057 : MUX2_X1 port map( A => registers_27_31_port, B => d_in(31), S => 
                           n700, Z => n3174);
   U1058 : MUX2_X1 port map( A => registers_27_30_port, B => d_in(30), S => 
                           n700, Z => n3173);
   U1059 : MUX2_X1 port map( A => registers_27_29_port, B => d_in(29), S => 
                           n700, Z => n3172);
   U1060 : MUX2_X1 port map( A => registers_27_28_port, B => d_in(28), S => 
                           n700, Z => n3171);
   U1061 : MUX2_X1 port map( A => registers_27_27_port, B => d_in(27), S => 
                           n700, Z => n3170);
   U1062 : MUX2_X1 port map( A => registers_27_26_port, B => d_in(26), S => 
                           n700, Z => n3169);
   U1063 : MUX2_X1 port map( A => registers_27_25_port, B => d_in(25), S => 
                           n700, Z => n3168);
   U1064 : MUX2_X1 port map( A => registers_27_24_port, B => d_in(24), S => 
                           n700, Z => n3167);
   U1065 : MUX2_X1 port map( A => registers_27_23_port, B => d_in(23), S => 
                           n700, Z => n3166);
   U1066 : MUX2_X1 port map( A => registers_27_22_port, B => d_in(22), S => 
                           n700, Z => n3165);
   U1067 : MUX2_X1 port map( A => registers_27_21_port, B => d_in(21), S => 
                           n700, Z => n3164);
   U1068 : MUX2_X1 port map( A => registers_27_20_port, B => d_in(20), S => 
                           n700, Z => n3163);
   U1069 : MUX2_X1 port map( A => registers_27_19_port, B => d_in(19), S => 
                           n700, Z => n3162);
   U1070 : MUX2_X1 port map( A => registers_27_18_port, B => d_in(18), S => 
                           n700, Z => n3161);
   U1071 : MUX2_X1 port map( A => registers_27_17_port, B => d_in(17), S => 
                           n700, Z => n3160);
   U1072 : MUX2_X1 port map( A => registers_27_16_port, B => d_in(16), S => 
                           n700, Z => n3159);
   U1073 : MUX2_X1 port map( A => registers_27_15_port, B => d_in(15), S => 
                           n700, Z => n3158);
   U1074 : MUX2_X1 port map( A => registers_27_14_port, B => d_in(14), S => 
                           n700, Z => n3157);
   U1075 : MUX2_X1 port map( A => registers_27_13_port, B => d_in(13), S => 
                           n700, Z => n3156);
   U1076 : MUX2_X1 port map( A => registers_27_12_port, B => d_in(12), S => 
                           n700, Z => n3155);
   U1077 : MUX2_X1 port map( A => registers_27_11_port, B => d_in(11), S => 
                           n700, Z => n3154);
   U1078 : MUX2_X1 port map( A => registers_27_10_port, B => d_in(10), S => 
                           n700, Z => n3153);
   U1079 : MUX2_X1 port map( A => registers_27_9_port, B => d_in(9), S => n700,
                           Z => n3152);
   U1080 : MUX2_X1 port map( A => registers_27_8_port, B => d_in(8), S => n700,
                           Z => n3151);
   U1081 : MUX2_X1 port map( A => registers_27_7_port, B => d_in(7), S => n700,
                           Z => n3150);
   U1082 : MUX2_X1 port map( A => registers_27_6_port, B => d_in(6), S => n700,
                           Z => n3149);
   U1083 : MUX2_X1 port map( A => registers_27_5_port, B => d_in(5), S => n700,
                           Z => n3148);
   U1084 : MUX2_X1 port map( A => registers_27_4_port, B => d_in(4), S => n700,
                           Z => n3147);
   U1085 : MUX2_X1 port map( A => registers_27_3_port, B => d_in(3), S => n700,
                           Z => n3146);
   U1086 : MUX2_X1 port map( A => registers_27_2_port, B => d_in(2), S => n700,
                           Z => n3145);
   U1087 : MUX2_X1 port map( A => registers_27_1_port, B => d_in(1), S => n700,
                           Z => n3144);
   U1088 : MUX2_X1 port map( A => registers_27_0_port, B => d_in(0), S => n700,
                           Z => n3143);
   U1089 : AND3_X1 port map( A1 => wr_addr(3), A2 => n664, A3 => n690, ZN => 
                           n697);
   U1090 : INV_X1 port map( A => wr_addr(2), ZN => n664);
   U1091 : MUX2_X1 port map( A => registers_28_31_port, B => d_in(31), S => 
                           n701, Z => n3142);
   U1092 : MUX2_X1 port map( A => registers_28_30_port, B => d_in(30), S => 
                           n701, Z => n3141);
   U1093 : MUX2_X1 port map( A => registers_28_29_port, B => d_in(29), S => 
                           n701, Z => n3140);
   U1094 : MUX2_X1 port map( A => registers_28_28_port, B => d_in(28), S => 
                           n701, Z => n3139);
   U1095 : MUX2_X1 port map( A => registers_28_27_port, B => d_in(27), S => 
                           n701, Z => n3138);
   U1096 : MUX2_X1 port map( A => registers_28_26_port, B => d_in(26), S => 
                           n701, Z => n3137);
   U1097 : MUX2_X1 port map( A => registers_28_25_port, B => d_in(25), S => 
                           n701, Z => n3136);
   U1098 : MUX2_X1 port map( A => registers_28_24_port, B => d_in(24), S => 
                           n701, Z => n3135);
   U1099 : MUX2_X1 port map( A => registers_28_23_port, B => d_in(23), S => 
                           n701, Z => n3134);
   U1100 : MUX2_X1 port map( A => registers_28_22_port, B => d_in(22), S => 
                           n701, Z => n3133);
   U1101 : MUX2_X1 port map( A => registers_28_21_port, B => d_in(21), S => 
                           n701, Z => n3132);
   U1102 : MUX2_X1 port map( A => registers_28_20_port, B => d_in(20), S => 
                           n701, Z => n3131);
   U1103 : MUX2_X1 port map( A => registers_28_19_port, B => d_in(19), S => 
                           n701, Z => n3130);
   U1104 : MUX2_X1 port map( A => registers_28_18_port, B => d_in(18), S => 
                           n701, Z => n3129);
   U1105 : MUX2_X1 port map( A => registers_28_17_port, B => d_in(17), S => 
                           n701, Z => n3128);
   U1106 : MUX2_X1 port map( A => registers_28_16_port, B => d_in(16), S => 
                           n701, Z => n3127);
   U1107 : MUX2_X1 port map( A => registers_28_15_port, B => d_in(15), S => 
                           n701, Z => n3126);
   U1108 : MUX2_X1 port map( A => registers_28_14_port, B => d_in(14), S => 
                           n701, Z => n3125);
   U1109 : MUX2_X1 port map( A => registers_28_13_port, B => d_in(13), S => 
                           n701, Z => n3124);
   U1110 : MUX2_X1 port map( A => registers_28_12_port, B => d_in(12), S => 
                           n701, Z => n3123);
   U1111 : MUX2_X1 port map( A => registers_28_11_port, B => d_in(11), S => 
                           n701, Z => n3122);
   U1112 : MUX2_X1 port map( A => registers_28_10_port, B => d_in(10), S => 
                           n701, Z => n3121);
   U1113 : MUX2_X1 port map( A => registers_28_9_port, B => d_in(9), S => n701,
                           Z => n3120);
   U1114 : MUX2_X1 port map( A => registers_28_8_port, B => d_in(8), S => n701,
                           Z => n3119);
   U1115 : MUX2_X1 port map( A => registers_28_7_port, B => d_in(7), S => n701,
                           Z => n3118);
   U1116 : MUX2_X1 port map( A => registers_28_6_port, B => d_in(6), S => n701,
                           Z => n3117);
   U1117 : MUX2_X1 port map( A => registers_28_5_port, B => d_in(5), S => n701,
                           Z => n3116);
   U1118 : MUX2_X1 port map( A => registers_28_4_port, B => d_in(4), S => n701,
                           Z => n3115);
   U1119 : MUX2_X1 port map( A => registers_28_3_port, B => d_in(3), S => n701,
                           Z => n3114);
   U1120 : MUX2_X1 port map( A => registers_28_2_port, B => d_in(2), S => n701,
                           Z => n3113);
   U1121 : MUX2_X1 port map( A => registers_28_1_port, B => d_in(1), S => n701,
                           Z => n3112);
   U1122 : MUX2_X1 port map( A => registers_28_0_port, B => d_in(0), S => n701,
                           Z => n3111);
   U1123 : NOR2_X1 port map( A1 => wr_addr(0), A2 => wr_addr(1), ZN => n668);
   U1124 : MUX2_X1 port map( A => registers_29_31_port, B => d_in(31), S => 
                           n703, Z => n3110);
   U1125 : MUX2_X1 port map( A => registers_29_30_port, B => d_in(30), S => 
                           n703, Z => n3109);
   U1126 : MUX2_X1 port map( A => registers_29_29_port, B => d_in(29), S => 
                           n703, Z => n3108);
   U1127 : MUX2_X1 port map( A => registers_29_28_port, B => d_in(28), S => 
                           n703, Z => n3107);
   U1128 : MUX2_X1 port map( A => registers_29_27_port, B => d_in(27), S => 
                           n703, Z => n3106);
   U1129 : MUX2_X1 port map( A => registers_29_26_port, B => d_in(26), S => 
                           n703, Z => n3105);
   U1130 : MUX2_X1 port map( A => registers_29_25_port, B => d_in(25), S => 
                           n703, Z => n3104);
   U1131 : MUX2_X1 port map( A => registers_29_24_port, B => d_in(24), S => 
                           n703, Z => n3103);
   U1132 : MUX2_X1 port map( A => registers_29_23_port, B => d_in(23), S => 
                           n703, Z => n3102);
   U1133 : MUX2_X1 port map( A => registers_29_22_port, B => d_in(22), S => 
                           n703, Z => n3101);
   U1134 : MUX2_X1 port map( A => registers_29_21_port, B => d_in(21), S => 
                           n703, Z => n3100);
   U1135 : MUX2_X1 port map( A => registers_29_20_port, B => d_in(20), S => 
                           n703, Z => n3099);
   U1136 : MUX2_X1 port map( A => registers_29_19_port, B => d_in(19), S => 
                           n703, Z => n3098);
   U1137 : MUX2_X1 port map( A => registers_29_18_port, B => d_in(18), S => 
                           n703, Z => n3097);
   U1138 : MUX2_X1 port map( A => registers_29_17_port, B => d_in(17), S => 
                           n703, Z => n3096);
   U1139 : MUX2_X1 port map( A => registers_29_16_port, B => d_in(16), S => 
                           n703, Z => n3095);
   U1140 : MUX2_X1 port map( A => registers_29_15_port, B => d_in(15), S => 
                           n703, Z => n3094);
   U1141 : MUX2_X1 port map( A => registers_29_14_port, B => d_in(14), S => 
                           n703, Z => n3093);
   U1142 : MUX2_X1 port map( A => registers_29_13_port, B => d_in(13), S => 
                           n703, Z => n3092);
   U1143 : MUX2_X1 port map( A => registers_29_12_port, B => d_in(12), S => 
                           n703, Z => n3091);
   U1144 : MUX2_X1 port map( A => registers_29_11_port, B => d_in(11), S => 
                           n703, Z => n3090);
   U1145 : MUX2_X1 port map( A => registers_29_10_port, B => d_in(10), S => 
                           n703, Z => n3089);
   U1146 : MUX2_X1 port map( A => registers_29_9_port, B => d_in(9), S => n703,
                           Z => n3088);
   U1147 : MUX2_X1 port map( A => registers_29_8_port, B => d_in(8), S => n703,
                           Z => n3087);
   U1148 : MUX2_X1 port map( A => registers_29_7_port, B => d_in(7), S => n703,
                           Z => n3086);
   U1149 : MUX2_X1 port map( A => registers_29_6_port, B => d_in(6), S => n703,
                           Z => n3085);
   U1150 : MUX2_X1 port map( A => registers_29_5_port, B => d_in(5), S => n703,
                           Z => n3084);
   U1151 : MUX2_X1 port map( A => registers_29_4_port, B => d_in(4), S => n703,
                           Z => n3083);
   U1152 : MUX2_X1 port map( A => registers_29_3_port, B => d_in(3), S => n703,
                           Z => n3082);
   U1153 : MUX2_X1 port map( A => registers_29_2_port, B => d_in(2), S => n703,
                           Z => n3081);
   U1154 : MUX2_X1 port map( A => registers_29_1_port, B => d_in(1), S => n703,
                           Z => n3080);
   U1155 : MUX2_X1 port map( A => registers_29_0_port, B => d_in(0), S => n703,
                           Z => n3079);
   U1156 : NOR2_X1 port map( A1 => n704, A2 => wr_addr(1), ZN => n658);
   U1157 : MUX2_X1 port map( A => registers_30_31_port, B => d_in(31), S => 
                           n705, Z => n3078);
   U1158 : MUX2_X1 port map( A => registers_30_30_port, B => d_in(30), S => 
                           n705, Z => n3077);
   U1159 : MUX2_X1 port map( A => registers_30_29_port, B => d_in(29), S => 
                           n705, Z => n3076);
   U1160 : MUX2_X1 port map( A => registers_30_28_port, B => d_in(28), S => 
                           n705, Z => n3075);
   U1161 : MUX2_X1 port map( A => registers_30_27_port, B => d_in(27), S => 
                           n705, Z => n3074);
   U1162 : MUX2_X1 port map( A => registers_30_26_port, B => d_in(26), S => 
                           n705, Z => n3073);
   U1163 : MUX2_X1 port map( A => registers_30_25_port, B => d_in(25), S => 
                           n705, Z => n3072);
   U1164 : MUX2_X1 port map( A => registers_30_24_port, B => d_in(24), S => 
                           n705, Z => n3071);
   U1165 : MUX2_X1 port map( A => registers_30_23_port, B => d_in(23), S => 
                           n705, Z => n3070);
   U1166 : MUX2_X1 port map( A => registers_30_22_port, B => d_in(22), S => 
                           n705, Z => n3069);
   U1167 : MUX2_X1 port map( A => registers_30_21_port, B => d_in(21), S => 
                           n705, Z => n3068);
   U1168 : MUX2_X1 port map( A => registers_30_20_port, B => d_in(20), S => 
                           n705, Z => n3067);
   U1169 : MUX2_X1 port map( A => registers_30_19_port, B => d_in(19), S => 
                           n705, Z => n3066);
   U1170 : MUX2_X1 port map( A => registers_30_18_port, B => d_in(18), S => 
                           n705, Z => n3065);
   U1171 : MUX2_X1 port map( A => registers_30_17_port, B => d_in(17), S => 
                           n705, Z => n3064);
   U1172 : MUX2_X1 port map( A => registers_30_16_port, B => d_in(16), S => 
                           n705, Z => n3063);
   U1173 : MUX2_X1 port map( A => registers_30_15_port, B => d_in(15), S => 
                           n705, Z => n3062);
   U1174 : MUX2_X1 port map( A => registers_30_14_port, B => d_in(14), S => 
                           n705, Z => n3061);
   U1175 : MUX2_X1 port map( A => registers_30_13_port, B => d_in(13), S => 
                           n705, Z => n3060);
   U1176 : MUX2_X1 port map( A => registers_30_12_port, B => d_in(12), S => 
                           n705, Z => n3059);
   U1177 : MUX2_X1 port map( A => registers_30_11_port, B => d_in(11), S => 
                           n705, Z => n3058);
   U1178 : MUX2_X1 port map( A => registers_30_10_port, B => d_in(10), S => 
                           n705, Z => n3057);
   U1179 : MUX2_X1 port map( A => registers_30_9_port, B => d_in(9), S => n705,
                           Z => n3056);
   U1180 : MUX2_X1 port map( A => registers_30_8_port, B => d_in(8), S => n705,
                           Z => n3055);
   U1181 : MUX2_X1 port map( A => registers_30_7_port, B => d_in(7), S => n705,
                           Z => n3054);
   U1182 : MUX2_X1 port map( A => registers_30_6_port, B => d_in(6), S => n705,
                           Z => n3053);
   U1183 : MUX2_X1 port map( A => registers_30_5_port, B => d_in(5), S => n705,
                           Z => n3052);
   U1184 : MUX2_X1 port map( A => registers_30_4_port, B => d_in(4), S => n705,
                           Z => n3051);
   U1185 : MUX2_X1 port map( A => registers_30_3_port, B => d_in(3), S => n705,
                           Z => n3050);
   U1186 : MUX2_X1 port map( A => registers_30_2_port, B => d_in(2), S => n705,
                           Z => n3049);
   U1187 : MUX2_X1 port map( A => registers_30_1_port, B => d_in(1), S => n705,
                           Z => n3048);
   U1188 : MUX2_X1 port map( A => registers_30_0_port, B => d_in(0), S => n705,
                           Z => n3047);
   U1189 : NOR2_X1 port map( A1 => n706, A2 => wr_addr(0), ZN => n661);
   U1190 : OAI21_X1 port map( B1 => n707, B2 => n289, A => n708, ZN => n3046);
   U1191 : AOI22_X1 port map( A1 => n709, A2 => d_in(31), B1 => d_link(31), B2 
                           => n710, ZN => n708);
   U1192 : NAND4_X1 port map( A1 => n711, A2 => n712, A3 => n713, A4 => n714, 
                           ZN => n3045);
   U1193 : AOI221_X1 port map( B1 => n715, B2 => registers_12_31_port, C1 => 
                           n716, C2 => registers_9_31_port, A => n717, ZN => 
                           n714);
   U1194 : OAI222_X1 port map( A1 => n415, A2 => n718, B1 => n1, B2 => n719, C1
                           => n225, C2 => n720, ZN => n717);
   U1195 : AOI221_X1 port map( B1 => n721, B2 => registers_4_31_port, C1 => 
                           n722, C2 => registers_20_31_port, A => n723, ZN => 
                           n713);
   U1196 : OAI22_X1 port map( A1 => n65, A2 => n724, B1 => n290, B2 => n725, ZN
                           => n723);
   U1197 : AOI221_X1 port map( B1 => n726, B2 => registers_15_31_port, C1 => 
                           n727, C2 => registers_30_31_port, A => n728, ZN => 
                           n712);
   U1198 : OAI222_X1 port map( A1 => n416, A2 => n729, B1 => n2, B2 => n730, C1
                           => n226, C2 => n731, ZN => n728);
   U1199 : AOI221_X1 port map( B1 => n732, B2 => d_in(31), C1 => n733, C2 => 
                           d_out2_31_port, A => n734, ZN => n711);
   U1200 : OAI22_X1 port map( A1 => n735, A2 => n736, B1 => n289, B2 => n737, 
                           ZN => n734);
   U1201 : NOR4_X1 port map( A1 => n738, A2 => n739, A3 => n740, A4 => n741, ZN
                           => n735);
   U1202 : OAI221_X1 port map( B1 => n159, B2 => n742, C1 => n541, C2 => n743, 
                           A => n744, ZN => n741);
   U1203 : AOI22_X1 port map( A1 => n745, A2 => registers_22_31_port, B1 => 
                           n746, B2 => registers_19_31_port, ZN => n744);
   U1204 : OAI221_X1 port map( B1 => n160, B2 => n747, C1 => n542, C2 => n748, 
                           A => n749, ZN => n740);
   U1205 : AOI22_X1 port map( A1 => n750, A2 => registers_28_31_port, B1 => 
                           n751, B2 => registers_25_31_port, ZN => n749);
   U1206 : OAI221_X1 port map( B1 => n161, B2 => n752, C1 => n543, C2 => n753, 
                           A => n754, ZN => n739);
   U1207 : AOI22_X1 port map( A1 => n755, A2 => registers_3_31_port, B1 => n756
                           , B2 => registers_6_31_port, ZN => n754);
   U1208 : OAI221_X1 port map( B1 => n162, B2 => n757, C1 => n544, C2 => n758, 
                           A => n759, ZN => n738);
   U1209 : AOI22_X1 port map( A1 => n760, A2 => registers_11_31_port, B1 => 
                           n761, B2 => registers_14_31_port, ZN => n759);
   U1210 : OAI21_X1 port map( B1 => n707, B2 => n322, A => n762, ZN => n3044);
   U1211 : AOI22_X1 port map( A1 => n709, A2 => d_in(30), B1 => d_link(30), B2 
                           => n710, ZN => n762);
   U1212 : NAND4_X1 port map( A1 => n763, A2 => n764, A3 => n765, A4 => n766, 
                           ZN => n3043);
   U1213 : AOI221_X1 port map( B1 => n715, B2 => registers_12_30_port, C1 => 
                           n716, C2 => registers_9_30_port, A => n767, ZN => 
                           n766);
   U1214 : OAI222_X1 port map( A1 => n417, A2 => n718, B1 => n3, B2 => n719, C1
                           => n227, C2 => n720, ZN => n767);
   U1215 : AOI221_X1 port map( B1 => n721, B2 => registers_4_30_port, C1 => 
                           n722, C2 => registers_20_30_port, A => n768, ZN => 
                           n765);
   U1216 : OAI22_X1 port map( A1 => n66, A2 => n724, B1 => n291, B2 => n725, ZN
                           => n768);
   U1217 : AOI221_X1 port map( B1 => n726, B2 => registers_15_30_port, C1 => 
                           n727, C2 => registers_30_30_port, A => n769, ZN => 
                           n764);
   U1218 : OAI222_X1 port map( A1 => n418, A2 => n729, B1 => n4, B2 => n730, C1
                           => n228, C2 => n731, ZN => n769);
   U1219 : AOI221_X1 port map( B1 => registers_31_30_port, B2 => n770, C1 => 
                           n771, C2 => n772, A => n773, ZN => n763);
   U1220 : OAI22_X1 port map( A1 => n2949, A2 => n774, B1 => n775, B2 => n776, 
                           ZN => n773);
   U1221 : INV_X1 port map( A => d_in(30), ZN => n775);
   U1222 : NAND4_X1 port map( A1 => n777, A2 => n778, A3 => n779, A4 => n780, 
                           ZN => n772);
   U1223 : AOI221_X1 port map( B1 => n760, B2 => registers_11_30_port, C1 => 
                           n761, C2 => registers_14_30_port, A => n781, ZN => 
                           n780);
   U1224 : OAI22_X1 port map( A1 => n354, A2 => n758, B1 => n98, B2 => n757, ZN
                           => n781);
   U1225 : INV_X1 port map( A => n782, ZN => n779);
   U1226 : OAI221_X1 port map( B1 => n752, B2 => n164, C1 => n753, C2 => n480, 
                           A => n783, ZN => n782);
   U1227 : AOI22_X1 port map( A1 => registers_6_30_port, A2 => n756, B1 => 
                           registers_3_30_port, B2 => n755, ZN => n783);
   U1228 : INV_X1 port map( A => n784, ZN => n778);
   U1229 : OAI221_X1 port map( B1 => n747, B2 => n163, C1 => n748, C2 => n479, 
                           A => n785, ZN => n784);
   U1230 : AOI22_X1 port map( A1 => registers_25_30_port, A2 => n751, B1 => 
                           registers_28_30_port, B2 => n750, ZN => n785);
   U1231 : AOI221_X1 port map( B1 => n745, B2 => registers_22_30_port, C1 => 
                           n746, C2 => registers_19_30_port, A => n786, ZN => 
                           n777);
   U1232 : OAI22_X1 port map( A1 => n353, A2 => n743, B1 => n97, B2 => n742, ZN
                           => n786);
   U1233 : OAI21_X1 port map( B1 => n707, B2 => n323, A => n787, ZN => n3042);
   U1234 : AOI22_X1 port map( A1 => n709, A2 => d_in(29), B1 => d_link(29), B2 
                           => n710, ZN => n787);
   U1235 : NAND4_X1 port map( A1 => n788, A2 => n789, A3 => n790, A4 => n791, 
                           ZN => n3041);
   U1236 : AOI221_X1 port map( B1 => n715, B2 => registers_12_29_port, C1 => 
                           n716, C2 => registers_9_29_port, A => n792, ZN => 
                           n791);
   U1237 : OAI222_X1 port map( A1 => n419, A2 => n718, B1 => n5, B2 => n719, C1
                           => n229, C2 => n720, ZN => n792);
   U1238 : AOI221_X1 port map( B1 => n721, B2 => registers_4_29_port, C1 => 
                           n722, C2 => registers_20_29_port, A => n793, ZN => 
                           n790);
   U1239 : OAI22_X1 port map( A1 => n67, A2 => n724, B1 => n292, B2 => n725, ZN
                           => n793);
   U1240 : AOI221_X1 port map( B1 => n726, B2 => registers_15_29_port, C1 => 
                           n727, C2 => registers_30_29_port, A => n794, ZN => 
                           n789);
   U1241 : OAI222_X1 port map( A1 => n420, A2 => n729, B1 => n6, B2 => n730, C1
                           => n230, C2 => n731, ZN => n794);
   U1242 : AOI221_X1 port map( B1 => registers_31_29_port, B2 => n770, C1 => 
                           n771, C2 => n795, A => n796, ZN => n788);
   U1243 : OAI22_X1 port map( A1 => n2948, A2 => n774, B1 => n797, B2 => n776, 
                           ZN => n796);
   U1244 : INV_X1 port map( A => d_in(29), ZN => n797);
   U1245 : NAND4_X1 port map( A1 => n798, A2 => n799, A3 => n800, A4 => n801, 
                           ZN => n795);
   U1246 : AOI221_X1 port map( B1 => n760, B2 => registers_11_29_port, C1 => 
                           n761, C2 => registers_14_29_port, A => n802, ZN => 
                           n801);
   U1247 : OAI22_X1 port map( A1 => n356, A2 => n758, B1 => n100, B2 => n757, 
                           ZN => n802);
   U1248 : INV_X1 port map( A => n803, ZN => n800);
   U1249 : OAI221_X1 port map( B1 => n752, B2 => n166, C1 => n753, C2 => n482, 
                           A => n804, ZN => n803);
   U1250 : AOI22_X1 port map( A1 => registers_6_29_port, A2 => n756, B1 => 
                           registers_3_29_port, B2 => n755, ZN => n804);
   U1251 : INV_X1 port map( A => n805, ZN => n799);
   U1252 : OAI221_X1 port map( B1 => n747, B2 => n165, C1 => n748, C2 => n481, 
                           A => n806, ZN => n805);
   U1253 : AOI22_X1 port map( A1 => registers_25_29_port, A2 => n751, B1 => 
                           registers_28_29_port, B2 => n750, ZN => n806);
   U1254 : AOI221_X1 port map( B1 => n745, B2 => registers_22_29_port, C1 => 
                           n746, C2 => registers_19_29_port, A => n807, ZN => 
                           n798);
   U1255 : OAI22_X1 port map( A1 => n355, A2 => n743, B1 => n99, B2 => n742, ZN
                           => n807);
   U1256 : OAI21_X1 port map( B1 => n707, B2 => n324, A => n808, ZN => n3040);
   U1257 : AOI22_X1 port map( A1 => n709, A2 => d_in(28), B1 => d_link(28), B2 
                           => n710, ZN => n808);
   U1258 : NAND4_X1 port map( A1 => n809, A2 => n810, A3 => n811, A4 => n812, 
                           ZN => n3039);
   U1259 : AOI221_X1 port map( B1 => n715, B2 => registers_12_28_port, C1 => 
                           n716, C2 => registers_9_28_port, A => n813, ZN => 
                           n812);
   U1260 : OAI222_X1 port map( A1 => n421, A2 => n718, B1 => n7, B2 => n719, C1
                           => n231, C2 => n720, ZN => n813);
   U1261 : AOI221_X1 port map( B1 => n721, B2 => registers_4_28_port, C1 => 
                           n722, C2 => registers_20_28_port, A => n814, ZN => 
                           n811);
   U1262 : OAI22_X1 port map( A1 => n68, A2 => n724, B1 => n293, B2 => n725, ZN
                           => n814);
   U1263 : AOI221_X1 port map( B1 => n726, B2 => registers_15_28_port, C1 => 
                           n727, C2 => registers_30_28_port, A => n815, ZN => 
                           n810);
   U1264 : OAI222_X1 port map( A1 => n422, A2 => n729, B1 => n8, B2 => n730, C1
                           => n232, C2 => n731, ZN => n815);
   U1265 : AOI221_X1 port map( B1 => registers_31_28_port, B2 => n770, C1 => 
                           n771, C2 => n816, A => n817, ZN => n809);
   U1266 : OAI22_X1 port map( A1 => n2947, A2 => n774, B1 => n818, B2 => n776, 
                           ZN => n817);
   U1267 : INV_X1 port map( A => d_in(28), ZN => n818);
   U1268 : NAND4_X1 port map( A1 => n819, A2 => n820, A3 => n821, A4 => n822, 
                           ZN => n816);
   U1269 : AOI221_X1 port map( B1 => n760, B2 => registers_11_28_port, C1 => 
                           n761, C2 => registers_14_28_port, A => n823, ZN => 
                           n822);
   U1270 : OAI22_X1 port map( A1 => n358, A2 => n758, B1 => n102, B2 => n757, 
                           ZN => n823);
   U1271 : INV_X1 port map( A => n824, ZN => n821);
   U1272 : OAI221_X1 port map( B1 => n752, B2 => n168, C1 => n753, C2 => n484, 
                           A => n825, ZN => n824);
   U1273 : AOI22_X1 port map( A1 => registers_6_28_port, A2 => n756, B1 => 
                           registers_3_28_port, B2 => n755, ZN => n825);
   U1274 : INV_X1 port map( A => n826, ZN => n820);
   U1275 : OAI221_X1 port map( B1 => n747, B2 => n167, C1 => n748, C2 => n483, 
                           A => n827, ZN => n826);
   U1276 : AOI22_X1 port map( A1 => registers_25_28_port, A2 => n751, B1 => 
                           registers_28_28_port, B2 => n750, ZN => n827);
   U1277 : AOI221_X1 port map( B1 => n745, B2 => registers_22_28_port, C1 => 
                           n746, C2 => registers_19_28_port, A => n828, ZN => 
                           n819);
   U1278 : OAI22_X1 port map( A1 => n357, A2 => n743, B1 => n101, B2 => n742, 
                           ZN => n828);
   U1279 : OAI21_X1 port map( B1 => n707, B2 => n325, A => n829, ZN => n3038);
   U1280 : AOI22_X1 port map( A1 => n709, A2 => d_in(27), B1 => d_link(27), B2 
                           => n710, ZN => n829);
   U1281 : NAND4_X1 port map( A1 => n830, A2 => n831, A3 => n832, A4 => n833, 
                           ZN => n3037);
   U1282 : AOI221_X1 port map( B1 => n715, B2 => registers_12_27_port, C1 => 
                           n716, C2 => registers_9_27_port, A => n834, ZN => 
                           n833);
   U1283 : OAI222_X1 port map( A1 => n423, A2 => n718, B1 => n9, B2 => n719, C1
                           => n233, C2 => n720, ZN => n834);
   U1284 : AOI221_X1 port map( B1 => n721, B2 => registers_4_27_port, C1 => 
                           n722, C2 => registers_20_27_port, A => n835, ZN => 
                           n832);
   U1285 : OAI22_X1 port map( A1 => n69, A2 => n724, B1 => n294, B2 => n725, ZN
                           => n835);
   U1286 : AOI221_X1 port map( B1 => n726, B2 => registers_15_27_port, C1 => 
                           n727, C2 => registers_30_27_port, A => n836, ZN => 
                           n831);
   U1287 : OAI222_X1 port map( A1 => n424, A2 => n729, B1 => n10, B2 => n730, 
                           C1 => n234, C2 => n731, ZN => n836);
   U1288 : AOI221_X1 port map( B1 => registers_31_27_port, B2 => n770, C1 => 
                           n771, C2 => n837, A => n838, ZN => n830);
   U1289 : OAI22_X1 port map( A1 => n2946, A2 => n774, B1 => n839, B2 => n776, 
                           ZN => n838);
   U1290 : INV_X1 port map( A => d_in(27), ZN => n839);
   U1291 : NAND4_X1 port map( A1 => n840, A2 => n841, A3 => n842, A4 => n843, 
                           ZN => n837);
   U1292 : AOI221_X1 port map( B1 => n760, B2 => registers_11_27_port, C1 => 
                           n761, C2 => registers_14_27_port, A => n844, ZN => 
                           n843);
   U1293 : OAI22_X1 port map( A1 => n360, A2 => n758, B1 => n104, B2 => n757, 
                           ZN => n844);
   U1294 : INV_X1 port map( A => n845, ZN => n842);
   U1295 : OAI221_X1 port map( B1 => n752, B2 => n170, C1 => n753, C2 => n486, 
                           A => n846, ZN => n845);
   U1296 : AOI22_X1 port map( A1 => registers_6_27_port, A2 => n756, B1 => 
                           registers_3_27_port, B2 => n755, ZN => n846);
   U1297 : INV_X1 port map( A => n847, ZN => n841);
   U1298 : OAI221_X1 port map( B1 => n747, B2 => n169, C1 => n748, C2 => n485, 
                           A => n848, ZN => n847);
   U1299 : AOI22_X1 port map( A1 => registers_25_27_port, A2 => n751, B1 => 
                           registers_28_27_port, B2 => n750, ZN => n848);
   U1300 : AOI221_X1 port map( B1 => n745, B2 => registers_22_27_port, C1 => 
                           n746, C2 => registers_19_27_port, A => n849, ZN => 
                           n840);
   U1301 : OAI22_X1 port map( A1 => n359, A2 => n743, B1 => n103, B2 => n742, 
                           ZN => n849);
   U1302 : OAI21_X1 port map( B1 => n707, B2 => n326, A => n850, ZN => n3036);
   U1303 : AOI22_X1 port map( A1 => n709, A2 => d_in(26), B1 => d_link(26), B2 
                           => n710, ZN => n850);
   U1304 : NAND4_X1 port map( A1 => n851, A2 => n852, A3 => n853, A4 => n854, 
                           ZN => n3035);
   U1305 : AOI221_X1 port map( B1 => n715, B2 => registers_12_26_port, C1 => 
                           n716, C2 => registers_9_26_port, A => n855, ZN => 
                           n854);
   U1306 : OAI222_X1 port map( A1 => n425, A2 => n718, B1 => n11, B2 => n719, 
                           C1 => n235, C2 => n720, ZN => n855);
   U1307 : AOI221_X1 port map( B1 => n721, B2 => registers_4_26_port, C1 => 
                           n722, C2 => registers_20_26_port, A => n856, ZN => 
                           n853);
   U1308 : OAI22_X1 port map( A1 => n70, A2 => n724, B1 => n295, B2 => n725, ZN
                           => n856);
   U1309 : AOI221_X1 port map( B1 => n726, B2 => registers_15_26_port, C1 => 
                           n727, C2 => registers_30_26_port, A => n857, ZN => 
                           n852);
   U1310 : OAI222_X1 port map( A1 => n426, A2 => n729, B1 => n12, B2 => n730, 
                           C1 => n236, C2 => n731, ZN => n857);
   U1311 : AOI221_X1 port map( B1 => registers_31_26_port, B2 => n770, C1 => 
                           n771, C2 => n858, A => n859, ZN => n851);
   U1312 : OAI22_X1 port map( A1 => n2945, A2 => n774, B1 => n860, B2 => n776, 
                           ZN => n859);
   U1313 : INV_X1 port map( A => d_in(26), ZN => n860);
   U1314 : NAND4_X1 port map( A1 => n861, A2 => n862, A3 => n863, A4 => n864, 
                           ZN => n858);
   U1315 : AOI221_X1 port map( B1 => n760, B2 => registers_11_26_port, C1 => 
                           n761, C2 => registers_14_26_port, A => n865, ZN => 
                           n864);
   U1316 : OAI22_X1 port map( A1 => n362, A2 => n758, B1 => n106, B2 => n757, 
                           ZN => n865);
   U1317 : INV_X1 port map( A => n866, ZN => n863);
   U1318 : OAI221_X1 port map( B1 => n752, B2 => n172, C1 => n753, C2 => n488, 
                           A => n867, ZN => n866);
   U1319 : AOI22_X1 port map( A1 => registers_6_26_port, A2 => n756, B1 => 
                           registers_3_26_port, B2 => n755, ZN => n867);
   U1320 : INV_X1 port map( A => n868, ZN => n862);
   U1321 : OAI221_X1 port map( B1 => n747, B2 => n171, C1 => n748, C2 => n487, 
                           A => n869, ZN => n868);
   U1322 : AOI22_X1 port map( A1 => registers_25_26_port, A2 => n751, B1 => 
                           registers_28_26_port, B2 => n750, ZN => n869);
   U1323 : AOI221_X1 port map( B1 => n745, B2 => registers_22_26_port, C1 => 
                           n746, C2 => registers_19_26_port, A => n870, ZN => 
                           n861);
   U1324 : OAI22_X1 port map( A1 => n361, A2 => n743, B1 => n105, B2 => n742, 
                           ZN => n870);
   U1325 : OAI21_X1 port map( B1 => n707, B2 => n327, A => n871, ZN => n3034);
   U1326 : AOI22_X1 port map( A1 => n709, A2 => d_in(25), B1 => d_link(25), B2 
                           => n710, ZN => n871);
   U1327 : NAND4_X1 port map( A1 => n872, A2 => n873, A3 => n874, A4 => n875, 
                           ZN => n3033);
   U1328 : AOI221_X1 port map( B1 => n715, B2 => registers_12_25_port, C1 => 
                           n716, C2 => registers_9_25_port, A => n876, ZN => 
                           n875);
   U1329 : OAI222_X1 port map( A1 => n427, A2 => n718, B1 => n13, B2 => n719, 
                           C1 => n237, C2 => n720, ZN => n876);
   U1330 : AOI221_X1 port map( B1 => n721, B2 => registers_4_25_port, C1 => 
                           n722, C2 => registers_20_25_port, A => n877, ZN => 
                           n874);
   U1331 : OAI22_X1 port map( A1 => n71, A2 => n724, B1 => n296, B2 => n725, ZN
                           => n877);
   U1332 : AOI221_X1 port map( B1 => n726, B2 => registers_15_25_port, C1 => 
                           n727, C2 => registers_30_25_port, A => n878, ZN => 
                           n873);
   U1333 : OAI222_X1 port map( A1 => n428, A2 => n729, B1 => n14, B2 => n730, 
                           C1 => n238, C2 => n731, ZN => n878);
   U1334 : AOI221_X1 port map( B1 => registers_31_25_port, B2 => n770, C1 => 
                           n771, C2 => n879, A => n880, ZN => n872);
   U1335 : OAI22_X1 port map( A1 => n2944, A2 => n774, B1 => n881, B2 => n776, 
                           ZN => n880);
   U1336 : INV_X1 port map( A => d_in(25), ZN => n881);
   U1337 : NAND4_X1 port map( A1 => n882, A2 => n883, A3 => n884, A4 => n885, 
                           ZN => n879);
   U1338 : AOI221_X1 port map( B1 => n760, B2 => registers_11_25_port, C1 => 
                           n761, C2 => registers_14_25_port, A => n886, ZN => 
                           n885);
   U1339 : OAI22_X1 port map( A1 => n364, A2 => n758, B1 => n108, B2 => n757, 
                           ZN => n886);
   U1340 : INV_X1 port map( A => n887, ZN => n884);
   U1341 : OAI221_X1 port map( B1 => n752, B2 => n174, C1 => n753, C2 => n490, 
                           A => n888, ZN => n887);
   U1342 : AOI22_X1 port map( A1 => registers_6_25_port, A2 => n756, B1 => 
                           registers_3_25_port, B2 => n755, ZN => n888);
   U1343 : INV_X1 port map( A => n889, ZN => n883);
   U1344 : OAI221_X1 port map( B1 => n747, B2 => n173, C1 => n748, C2 => n489, 
                           A => n890, ZN => n889);
   U1345 : AOI22_X1 port map( A1 => registers_25_25_port, A2 => n751, B1 => 
                           registers_28_25_port, B2 => n750, ZN => n890);
   U1346 : AOI221_X1 port map( B1 => n745, B2 => registers_22_25_port, C1 => 
                           n746, C2 => registers_19_25_port, A => n891, ZN => 
                           n882);
   U1347 : OAI22_X1 port map( A1 => n363, A2 => n743, B1 => n107, B2 => n742, 
                           ZN => n891);
   U1348 : OAI21_X1 port map( B1 => n707, B2 => n328, A => n892, ZN => n3032);
   U1349 : AOI22_X1 port map( A1 => n709, A2 => d_in(24), B1 => d_link(24), B2 
                           => n710, ZN => n892);
   U1350 : NAND4_X1 port map( A1 => n893, A2 => n894, A3 => n895, A4 => n896, 
                           ZN => n3031);
   U1351 : AOI221_X1 port map( B1 => n715, B2 => registers_12_24_port, C1 => 
                           n716, C2 => registers_9_24_port, A => n897, ZN => 
                           n896);
   U1352 : OAI222_X1 port map( A1 => n429, A2 => n718, B1 => n15, B2 => n719, 
                           C1 => n239, C2 => n720, ZN => n897);
   U1353 : AOI221_X1 port map( B1 => n721, B2 => registers_4_24_port, C1 => 
                           n722, C2 => registers_20_24_port, A => n898, ZN => 
                           n895);
   U1354 : OAI22_X1 port map( A1 => n72, A2 => n724, B1 => n297, B2 => n725, ZN
                           => n898);
   U1355 : AOI221_X1 port map( B1 => n726, B2 => registers_15_24_port, C1 => 
                           n727, C2 => registers_30_24_port, A => n899, ZN => 
                           n894);
   U1356 : OAI222_X1 port map( A1 => n430, A2 => n729, B1 => n16, B2 => n730, 
                           C1 => n240, C2 => n731, ZN => n899);
   U1357 : AOI221_X1 port map( B1 => registers_31_24_port, B2 => n770, C1 => 
                           n771, C2 => n900, A => n901, ZN => n893);
   U1358 : OAI22_X1 port map( A1 => n2943, A2 => n774, B1 => n902, B2 => n776, 
                           ZN => n901);
   U1359 : INV_X1 port map( A => d_in(24), ZN => n902);
   U1360 : NAND4_X1 port map( A1 => n903, A2 => n904, A3 => n905, A4 => n906, 
                           ZN => n900);
   U1361 : AOI221_X1 port map( B1 => n760, B2 => registers_11_24_port, C1 => 
                           n761, C2 => registers_14_24_port, A => n907, ZN => 
                           n906);
   U1362 : OAI22_X1 port map( A1 => n366, A2 => n758, B1 => n110, B2 => n757, 
                           ZN => n907);
   U1363 : INV_X1 port map( A => n908, ZN => n905);
   U1364 : OAI221_X1 port map( B1 => n752, B2 => n176, C1 => n753, C2 => n492, 
                           A => n909, ZN => n908);
   U1365 : AOI22_X1 port map( A1 => registers_6_24_port, A2 => n756, B1 => 
                           registers_3_24_port, B2 => n755, ZN => n909);
   U1366 : INV_X1 port map( A => n910, ZN => n904);
   U1367 : OAI221_X1 port map( B1 => n747, B2 => n175, C1 => n748, C2 => n491, 
                           A => n911, ZN => n910);
   U1368 : AOI22_X1 port map( A1 => registers_25_24_port, A2 => n751, B1 => 
                           registers_28_24_port, B2 => n750, ZN => n911);
   U1369 : AOI221_X1 port map( B1 => n745, B2 => registers_22_24_port, C1 => 
                           n746, C2 => registers_19_24_port, A => n912, ZN => 
                           n903);
   U1370 : OAI22_X1 port map( A1 => n365, A2 => n743, B1 => n109, B2 => n742, 
                           ZN => n912);
   U1371 : OAI21_X1 port map( B1 => n707, B2 => n329, A => n913, ZN => n3030);
   U1372 : AOI22_X1 port map( A1 => n709, A2 => d_in(23), B1 => d_link(23), B2 
                           => n710, ZN => n913);
   U1373 : NAND4_X1 port map( A1 => n914, A2 => n915, A3 => n916, A4 => n917, 
                           ZN => n3029);
   U1374 : AOI221_X1 port map( B1 => n715, B2 => registers_12_23_port, C1 => 
                           n716, C2 => registers_9_23_port, A => n918, ZN => 
                           n917);
   U1375 : OAI222_X1 port map( A1 => n431, A2 => n718, B1 => n17, B2 => n719, 
                           C1 => n241, C2 => n720, ZN => n918);
   U1376 : AOI221_X1 port map( B1 => n721, B2 => registers_4_23_port, C1 => 
                           n722, C2 => registers_20_23_port, A => n919, ZN => 
                           n916);
   U1377 : OAI22_X1 port map( A1 => n73, A2 => n724, B1 => n298, B2 => n725, ZN
                           => n919);
   U1378 : AOI221_X1 port map( B1 => n726, B2 => registers_15_23_port, C1 => 
                           n727, C2 => registers_30_23_port, A => n920, ZN => 
                           n915);
   U1379 : OAI222_X1 port map( A1 => n432, A2 => n729, B1 => n18_port, B2 => 
                           n730, C1 => n242, C2 => n731, ZN => n920);
   U1380 : AOI221_X1 port map( B1 => registers_31_23_port, B2 => n770, C1 => 
                           n771, C2 => n921, A => n922, ZN => n914);
   U1381 : OAI22_X1 port map( A1 => n2942, A2 => n774, B1 => n923, B2 => n776, 
                           ZN => n922);
   U1382 : INV_X1 port map( A => d_in(23), ZN => n923);
   U1383 : NAND4_X1 port map( A1 => n924, A2 => n925, A3 => n926, A4 => n927, 
                           ZN => n921);
   U1384 : AOI221_X1 port map( B1 => n760, B2 => registers_11_23_port, C1 => 
                           n761, C2 => registers_14_23_port, A => n928, ZN => 
                           n927);
   U1385 : OAI22_X1 port map( A1 => n368, A2 => n758, B1 => n112, B2 => n757, 
                           ZN => n928);
   U1386 : INV_X1 port map( A => n929, ZN => n926);
   U1387 : OAI221_X1 port map( B1 => n752, B2 => n178, C1 => n753, C2 => n494, 
                           A => n930, ZN => n929);
   U1388 : AOI22_X1 port map( A1 => registers_6_23_port, A2 => n756, B1 => 
                           registers_3_23_port, B2 => n755, ZN => n930);
   U1389 : INV_X1 port map( A => n931, ZN => n925);
   U1390 : OAI221_X1 port map( B1 => n747, B2 => n177, C1 => n748, C2 => n493, 
                           A => n932, ZN => n931);
   U1391 : AOI22_X1 port map( A1 => registers_25_23_port, A2 => n751, B1 => 
                           registers_28_23_port, B2 => n750, ZN => n932);
   U1392 : AOI221_X1 port map( B1 => n745, B2 => registers_22_23_port, C1 => 
                           n746, C2 => registers_19_23_port, A => n933, ZN => 
                           n924);
   U1393 : OAI22_X1 port map( A1 => n367, A2 => n743, B1 => n111, B2 => n742, 
                           ZN => n933);
   U1394 : OAI21_X1 port map( B1 => n707, B2 => n330, A => n934, ZN => n3028);
   U1395 : AOI22_X1 port map( A1 => n709, A2 => d_in(22), B1 => d_link(22), B2 
                           => n710, ZN => n934);
   U1396 : NAND4_X1 port map( A1 => n935, A2 => n936, A3 => n937, A4 => n938, 
                           ZN => n3027);
   U1397 : AOI221_X1 port map( B1 => n715, B2 => registers_12_22_port, C1 => 
                           n716, C2 => registers_9_22_port, A => n939, ZN => 
                           n938);
   U1398 : OAI222_X1 port map( A1 => n433, A2 => n718, B1 => n19, B2 => n719, 
                           C1 => n243, C2 => n720, ZN => n939);
   U1399 : AOI221_X1 port map( B1 => n721, B2 => registers_4_22_port, C1 => 
                           n722, C2 => registers_20_22_port, A => n940, ZN => 
                           n937);
   U1400 : OAI22_X1 port map( A1 => n74, A2 => n724, B1 => n299, B2 => n725, ZN
                           => n940);
   U1401 : AOI221_X1 port map( B1 => n726, B2 => registers_15_22_port, C1 => 
                           n727, C2 => registers_30_22_port, A => n941, ZN => 
                           n936);
   U1402 : OAI222_X1 port map( A1 => n434, A2 => n729, B1 => n20, B2 => n730, 
                           C1 => n244, C2 => n731, ZN => n941);
   U1403 : AOI221_X1 port map( B1 => registers_31_22_port, B2 => n770, C1 => 
                           n771, C2 => n942, A => n943, ZN => n935);
   U1404 : OAI22_X1 port map( A1 => n2941, A2 => n774, B1 => n944, B2 => n776, 
                           ZN => n943);
   U1405 : INV_X1 port map( A => d_in(22), ZN => n944);
   U1406 : NAND4_X1 port map( A1 => n945, A2 => n946, A3 => n947, A4 => n948, 
                           ZN => n942);
   U1407 : AOI221_X1 port map( B1 => n760, B2 => registers_11_22_port, C1 => 
                           n761, C2 => registers_14_22_port, A => n949, ZN => 
                           n948);
   U1408 : OAI22_X1 port map( A1 => n370, A2 => n758, B1 => n114, B2 => n757, 
                           ZN => n949);
   U1409 : INV_X1 port map( A => n950, ZN => n947);
   U1410 : OAI221_X1 port map( B1 => n752, B2 => n180, C1 => n753, C2 => n496, 
                           A => n951, ZN => n950);
   U1411 : AOI22_X1 port map( A1 => registers_6_22_port, A2 => n756, B1 => 
                           registers_3_22_port, B2 => n755, ZN => n951);
   U1412 : INV_X1 port map( A => n952, ZN => n946);
   U1413 : OAI221_X1 port map( B1 => n747, B2 => n179, C1 => n748, C2 => n495, 
                           A => n953, ZN => n952);
   U1414 : AOI22_X1 port map( A1 => registers_25_22_port, A2 => n751, B1 => 
                           registers_28_22_port, B2 => n750, ZN => n953);
   U1415 : AOI221_X1 port map( B1 => n745, B2 => registers_22_22_port, C1 => 
                           n746, C2 => registers_19_22_port, A => n954, ZN => 
                           n945);
   U1416 : OAI22_X1 port map( A1 => n369, A2 => n743, B1 => n113, B2 => n742, 
                           ZN => n954);
   U1417 : OAI21_X1 port map( B1 => n707, B2 => n331, A => n955, ZN => n3026);
   U1418 : AOI22_X1 port map( A1 => n709, A2 => d_in(21), B1 => d_link(21), B2 
                           => n710, ZN => n955);
   U1419 : NAND4_X1 port map( A1 => n956, A2 => n957, A3 => n958, A4 => n959, 
                           ZN => n3025);
   U1420 : AOI221_X1 port map( B1 => n715, B2 => registers_12_21_port, C1 => 
                           n716, C2 => registers_9_21_port, A => n960, ZN => 
                           n959);
   U1421 : OAI222_X1 port map( A1 => n435, A2 => n718, B1 => n21, B2 => n719, 
                           C1 => n245, C2 => n720, ZN => n960);
   U1422 : AOI221_X1 port map( B1 => n721, B2 => registers_4_21_port, C1 => 
                           n722, C2 => registers_20_21_port, A => n961, ZN => 
                           n958);
   U1423 : OAI22_X1 port map( A1 => n75, A2 => n724, B1 => n300, B2 => n725, ZN
                           => n961);
   U1424 : AOI221_X1 port map( B1 => n726, B2 => registers_15_21_port, C1 => 
                           n727, C2 => registers_30_21_port, A => n962, ZN => 
                           n957);
   U1425 : OAI222_X1 port map( A1 => n436, A2 => n729, B1 => n22, B2 => n730, 
                           C1 => n246, C2 => n731, ZN => n962);
   U1426 : AOI221_X1 port map( B1 => registers_31_21_port, B2 => n770, C1 => 
                           n771, C2 => n963, A => n964, ZN => n956);
   U1427 : OAI22_X1 port map( A1 => n2940, A2 => n774, B1 => n965, B2 => n776, 
                           ZN => n964);
   U1428 : INV_X1 port map( A => d_in(21), ZN => n965);
   U1429 : NAND4_X1 port map( A1 => n966, A2 => n967, A3 => n968, A4 => n969, 
                           ZN => n963);
   U1430 : AOI221_X1 port map( B1 => n760, B2 => registers_11_21_port, C1 => 
                           n761, C2 => registers_14_21_port, A => n970, ZN => 
                           n969);
   U1431 : OAI22_X1 port map( A1 => n372, A2 => n758, B1 => n116, B2 => n757, 
                           ZN => n970);
   U1432 : INV_X1 port map( A => n971, ZN => n968);
   U1433 : OAI221_X1 port map( B1 => n752, B2 => n182, C1 => n753, C2 => n498, 
                           A => n972, ZN => n971);
   U1434 : AOI22_X1 port map( A1 => registers_6_21_port, A2 => n756, B1 => 
                           registers_3_21_port, B2 => n755, ZN => n972);
   U1435 : INV_X1 port map( A => n973, ZN => n967);
   U1436 : OAI221_X1 port map( B1 => n747, B2 => n181, C1 => n748, C2 => n497, 
                           A => n974, ZN => n973);
   U1437 : AOI22_X1 port map( A1 => registers_25_21_port, A2 => n751, B1 => 
                           registers_28_21_port, B2 => n750, ZN => n974);
   U1438 : AOI221_X1 port map( B1 => n745, B2 => registers_22_21_port, C1 => 
                           n746, C2 => registers_19_21_port, A => n975, ZN => 
                           n966);
   U1439 : OAI22_X1 port map( A1 => n371, A2 => n743, B1 => n115, B2 => n742, 
                           ZN => n975);
   U1440 : OAI21_X1 port map( B1 => n707, B2 => n332, A => n976, ZN => n3024);
   U1441 : AOI22_X1 port map( A1 => n709, A2 => d_in(20), B1 => d_link(20), B2 
                           => n710, ZN => n976);
   U1442 : NAND4_X1 port map( A1 => n977, A2 => n978, A3 => n979, A4 => n980, 
                           ZN => n3023);
   U1443 : AOI221_X1 port map( B1 => n715, B2 => registers_12_20_port, C1 => 
                           n716, C2 => registers_9_20_port, A => n981, ZN => 
                           n980);
   U1444 : OAI222_X1 port map( A1 => n437, A2 => n718, B1 => n23, B2 => n719, 
                           C1 => n247, C2 => n720, ZN => n981);
   U1445 : AOI221_X1 port map( B1 => n721, B2 => registers_4_20_port, C1 => 
                           n722, C2 => registers_20_20_port, A => n982, ZN => 
                           n979);
   U1446 : OAI22_X1 port map( A1 => n76, A2 => n724, B1 => n301, B2 => n725, ZN
                           => n982);
   U1447 : AOI221_X1 port map( B1 => n726, B2 => registers_15_20_port, C1 => 
                           n727, C2 => registers_30_20_port, A => n983, ZN => 
                           n978);
   U1448 : OAI222_X1 port map( A1 => n438, A2 => n729, B1 => n24, B2 => n730, 
                           C1 => n248, C2 => n731, ZN => n983);
   U1449 : AOI221_X1 port map( B1 => registers_31_20_port, B2 => n770, C1 => 
                           n771, C2 => n984, A => n985, ZN => n977);
   U1450 : OAI22_X1 port map( A1 => n2939, A2 => n774, B1 => n986, B2 => n776, 
                           ZN => n985);
   U1451 : INV_X1 port map( A => d_in(20), ZN => n986);
   U1452 : NAND4_X1 port map( A1 => n987, A2 => n988, A3 => n989, A4 => n990, 
                           ZN => n984);
   U1453 : AOI221_X1 port map( B1 => n760, B2 => registers_11_20_port, C1 => 
                           n761, C2 => registers_14_20_port, A => n991, ZN => 
                           n990);
   U1454 : OAI22_X1 port map( A1 => n374, A2 => n758, B1 => n118, B2 => n757, 
                           ZN => n991);
   U1455 : INV_X1 port map( A => n992, ZN => n989);
   U1456 : OAI221_X1 port map( B1 => n752, B2 => n184, C1 => n753, C2 => n500, 
                           A => n993, ZN => n992);
   U1457 : AOI22_X1 port map( A1 => registers_6_20_port, A2 => n756, B1 => 
                           registers_3_20_port, B2 => n755, ZN => n993);
   U1458 : INV_X1 port map( A => n994, ZN => n988);
   U1459 : OAI221_X1 port map( B1 => n747, B2 => n183, C1 => n748, C2 => n499, 
                           A => n995, ZN => n994);
   U1460 : AOI22_X1 port map( A1 => registers_25_20_port, A2 => n751, B1 => 
                           registers_28_20_port, B2 => n750, ZN => n995);
   U1461 : AOI221_X1 port map( B1 => n745, B2 => registers_22_20_port, C1 => 
                           n746, C2 => registers_19_20_port, A => n996, ZN => 
                           n987);
   U1462 : OAI22_X1 port map( A1 => n373, A2 => n743, B1 => n117, B2 => n742, 
                           ZN => n996);
   U1463 : OAI21_X1 port map( B1 => n707, B2 => n333, A => n997, ZN => n3022);
   U1464 : AOI22_X1 port map( A1 => n709, A2 => d_in(19), B1 => d_link(19), B2 
                           => n710, ZN => n997);
   U1465 : NAND4_X1 port map( A1 => n998, A2 => n999, A3 => n1000, A4 => n1001,
                           ZN => n3021);
   U1466 : AOI221_X1 port map( B1 => n715, B2 => registers_12_19_port, C1 => 
                           n716, C2 => registers_9_19_port, A => n1002, ZN => 
                           n1001);
   U1467 : OAI222_X1 port map( A1 => n439, A2 => n718, B1 => n25, B2 => n719, 
                           C1 => n249, C2 => n720, ZN => n1002);
   U1468 : AOI221_X1 port map( B1 => n721, B2 => registers_4_19_port, C1 => 
                           n722, C2 => registers_20_19_port, A => n1003, ZN => 
                           n1000);
   U1469 : OAI22_X1 port map( A1 => n77, A2 => n724, B1 => n302, B2 => n725, ZN
                           => n1003);
   U1470 : AOI221_X1 port map( B1 => n726, B2 => registers_15_19_port, C1 => 
                           n727, C2 => registers_30_19_port, A => n1004, ZN => 
                           n999);
   U1471 : OAI222_X1 port map( A1 => n440, A2 => n729, B1 => n26, B2 => n730, 
                           C1 => n250, C2 => n731, ZN => n1004);
   U1472 : AOI221_X1 port map( B1 => registers_31_19_port, B2 => n770, C1 => 
                           n771, C2 => n1005, A => n1006, ZN => n998);
   U1473 : OAI22_X1 port map( A1 => n2938, A2 => n774, B1 => n1007, B2 => n776,
                           ZN => n1006);
   U1474 : INV_X1 port map( A => d_in(19), ZN => n1007);
   U1475 : NAND4_X1 port map( A1 => n1008, A2 => n1009, A3 => n1010, A4 => 
                           n1011, ZN => n1005);
   U1476 : AOI221_X1 port map( B1 => n760, B2 => registers_11_19_port, C1 => 
                           n761, C2 => registers_14_19_port, A => n1012, ZN => 
                           n1011);
   U1477 : OAI22_X1 port map( A1 => n376, A2 => n758, B1 => n120, B2 => n757, 
                           ZN => n1012);
   U1478 : INV_X1 port map( A => n1013, ZN => n1010);
   U1479 : OAI221_X1 port map( B1 => n752, B2 => n186, C1 => n753, C2 => n502, 
                           A => n1014, ZN => n1013);
   U1480 : AOI22_X1 port map( A1 => registers_6_19_port, A2 => n756, B1 => 
                           registers_3_19_port, B2 => n755, ZN => n1014);
   U1481 : INV_X1 port map( A => n1015, ZN => n1009);
   U1482 : OAI221_X1 port map( B1 => n747, B2 => n185, C1 => n748, C2 => n501, 
                           A => n1016, ZN => n1015);
   U1483 : AOI22_X1 port map( A1 => registers_25_19_port, A2 => n751, B1 => 
                           registers_28_19_port, B2 => n750, ZN => n1016);
   U1484 : AOI221_X1 port map( B1 => n745, B2 => registers_22_19_port, C1 => 
                           n746, C2 => registers_19_19_port, A => n1017, ZN => 
                           n1008);
   U1485 : OAI22_X1 port map( A1 => n375, A2 => n743, B1 => n119, B2 => n742, 
                           ZN => n1017);
   U1486 : OAI21_X1 port map( B1 => n707, B2 => n334, A => n1018, ZN => n3020);
   U1487 : AOI22_X1 port map( A1 => n709, A2 => d_in(18), B1 => d_link(18), B2 
                           => n710, ZN => n1018);
   U1488 : NAND4_X1 port map( A1 => n1019, A2 => n1020, A3 => n1021, A4 => 
                           n1022, ZN => n3019);
   U1489 : AOI221_X1 port map( B1 => n715, B2 => registers_12_18_port, C1 => 
                           n716, C2 => registers_9_18_port, A => n1023, ZN => 
                           n1022);
   U1490 : OAI222_X1 port map( A1 => n441, A2 => n718, B1 => n27, B2 => n719, 
                           C1 => n251, C2 => n720, ZN => n1023);
   U1491 : AOI221_X1 port map( B1 => n721, B2 => registers_4_18_port, C1 => 
                           n722, C2 => registers_20_18_port, A => n1024, ZN => 
                           n1021);
   U1492 : OAI22_X1 port map( A1 => n78, A2 => n724, B1 => n303, B2 => n725, ZN
                           => n1024);
   U1493 : AOI221_X1 port map( B1 => n726, B2 => registers_15_18_port, C1 => 
                           n727, C2 => registers_30_18_port, A => n1025, ZN => 
                           n1020);
   U1494 : OAI222_X1 port map( A1 => n442, A2 => n729, B1 => n28, B2 => n730, 
                           C1 => n252, C2 => n731, ZN => n1025);
   U1495 : AOI221_X1 port map( B1 => registers_31_18_port, B2 => n770, C1 => 
                           n771, C2 => n1026, A => n1027, ZN => n1019);
   U1496 : OAI22_X1 port map( A1 => n2937, A2 => n774, B1 => n1028, B2 => n776,
                           ZN => n1027);
   U1497 : INV_X1 port map( A => d_in(18), ZN => n1028);
   U1498 : NAND4_X1 port map( A1 => n1029, A2 => n1030, A3 => n1031, A4 => 
                           n1032, ZN => n1026);
   U1499 : AOI221_X1 port map( B1 => n760, B2 => registers_11_18_port, C1 => 
                           n761, C2 => registers_14_18_port, A => n1033, ZN => 
                           n1032);
   U1500 : OAI22_X1 port map( A1 => n378, A2 => n758, B1 => n122, B2 => n757, 
                           ZN => n1033);
   U1501 : INV_X1 port map( A => n1034, ZN => n1031);
   U1502 : OAI221_X1 port map( B1 => n752, B2 => n188, C1 => n753, C2 => n504, 
                           A => n1035, ZN => n1034);
   U1503 : AOI22_X1 port map( A1 => registers_6_18_port, A2 => n756, B1 => 
                           registers_3_18_port, B2 => n755, ZN => n1035);
   U1504 : INV_X1 port map( A => n1036, ZN => n1030);
   U1505 : OAI221_X1 port map( B1 => n747, B2 => n187, C1 => n748, C2 => n503, 
                           A => n1037, ZN => n1036);
   U1506 : AOI22_X1 port map( A1 => registers_25_18_port, A2 => n751, B1 => 
                           registers_28_18_port, B2 => n750, ZN => n1037);
   U1507 : AOI221_X1 port map( B1 => n745, B2 => registers_22_18_port, C1 => 
                           n746, C2 => registers_19_18_port, A => n1038, ZN => 
                           n1029);
   U1508 : OAI22_X1 port map( A1 => n377, A2 => n743, B1 => n121, B2 => n742, 
                           ZN => n1038);
   U1509 : OAI21_X1 port map( B1 => n707, B2 => n335, A => n1039, ZN => n3018);
   U1510 : AOI22_X1 port map( A1 => n709, A2 => d_in(17), B1 => d_link(17), B2 
                           => n710, ZN => n1039);
   U1511 : NAND4_X1 port map( A1 => n1040, A2 => n1041, A3 => n1042, A4 => 
                           n1043, ZN => n3017);
   U1512 : AOI221_X1 port map( B1 => n715, B2 => registers_12_17_port, C1 => 
                           n716, C2 => registers_9_17_port, A => n1044, ZN => 
                           n1043);
   U1513 : OAI222_X1 port map( A1 => n443, A2 => n718, B1 => n29, B2 => n719, 
                           C1 => n253, C2 => n720, ZN => n1044);
   U1514 : AOI221_X1 port map( B1 => n721, B2 => registers_4_17_port, C1 => 
                           n722, C2 => registers_20_17_port, A => n1045, ZN => 
                           n1042);
   U1515 : OAI22_X1 port map( A1 => n79, A2 => n724, B1 => n304, B2 => n725, ZN
                           => n1045);
   U1516 : AOI221_X1 port map( B1 => n726, B2 => registers_15_17_port, C1 => 
                           n727, C2 => registers_30_17_port, A => n1046, ZN => 
                           n1041);
   U1517 : OAI222_X1 port map( A1 => n444, A2 => n729, B1 => n30, B2 => n730, 
                           C1 => n254, C2 => n731, ZN => n1046);
   U1518 : AOI221_X1 port map( B1 => registers_31_17_port, B2 => n770, C1 => 
                           n771, C2 => n1047, A => n1048, ZN => n1040);
   U1519 : OAI22_X1 port map( A1 => n2936, A2 => n774, B1 => n1049, B2 => n776,
                           ZN => n1048);
   U1520 : INV_X1 port map( A => d_in(17), ZN => n1049);
   U1521 : NAND4_X1 port map( A1 => n1050, A2 => n1051, A3 => n1052, A4 => 
                           n1053, ZN => n1047);
   U1522 : AOI221_X1 port map( B1 => n760, B2 => registers_11_17_port, C1 => 
                           n761, C2 => registers_14_17_port, A => n1054, ZN => 
                           n1053);
   U1523 : OAI22_X1 port map( A1 => n380, A2 => n758, B1 => n124, B2 => n757, 
                           ZN => n1054);
   U1524 : INV_X1 port map( A => n1055, ZN => n1052);
   U1525 : OAI221_X1 port map( B1 => n752, B2 => n190, C1 => n753, C2 => n506, 
                           A => n1056, ZN => n1055);
   U1526 : AOI22_X1 port map( A1 => registers_6_17_port, A2 => n756, B1 => 
                           registers_3_17_port, B2 => n755, ZN => n1056);
   U1527 : INV_X1 port map( A => n1057, ZN => n1051);
   U1528 : OAI221_X1 port map( B1 => n747, B2 => n189, C1 => n748, C2 => n505, 
                           A => n1058, ZN => n1057);
   U1529 : AOI22_X1 port map( A1 => registers_25_17_port, A2 => n751, B1 => 
                           registers_28_17_port, B2 => n750, ZN => n1058);
   U1530 : AOI221_X1 port map( B1 => n745, B2 => registers_22_17_port, C1 => 
                           n746, C2 => registers_19_17_port, A => n1059, ZN => 
                           n1050);
   U1531 : OAI22_X1 port map( A1 => n379, A2 => n743, B1 => n123, B2 => n742, 
                           ZN => n1059);
   U1532 : OAI21_X1 port map( B1 => n707, B2 => n336, A => n1060, ZN => n3016);
   U1533 : AOI22_X1 port map( A1 => n709, A2 => d_in(16), B1 => d_link(16), B2 
                           => n710, ZN => n1060);
   U1534 : NAND4_X1 port map( A1 => n1061, A2 => n1062, A3 => n1063, A4 => 
                           n1064, ZN => n3015);
   U1535 : AOI221_X1 port map( B1 => n715, B2 => registers_12_16_port, C1 => 
                           n716, C2 => registers_9_16_port, A => n1065, ZN => 
                           n1064);
   U1536 : OAI222_X1 port map( A1 => n445, A2 => n718, B1 => n31, B2 => n719, 
                           C1 => n255, C2 => n720, ZN => n1065);
   U1537 : AOI221_X1 port map( B1 => n721, B2 => registers_4_16_port, C1 => 
                           n722, C2 => registers_20_16_port, A => n1066, ZN => 
                           n1063);
   U1538 : OAI22_X1 port map( A1 => n80, A2 => n724, B1 => n305, B2 => n725, ZN
                           => n1066);
   U1539 : AOI221_X1 port map( B1 => n726, B2 => registers_15_16_port, C1 => 
                           n727, C2 => registers_30_16_port, A => n1067, ZN => 
                           n1062);
   U1540 : OAI222_X1 port map( A1 => n446, A2 => n729, B1 => n32, B2 => n730, 
                           C1 => n256, C2 => n731, ZN => n1067);
   U1541 : AOI221_X1 port map( B1 => registers_31_16_port, B2 => n770, C1 => 
                           n771, C2 => n1068, A => n1069, ZN => n1061);
   U1542 : OAI22_X1 port map( A1 => n2935, A2 => n774, B1 => n1070, B2 => n776,
                           ZN => n1069);
   U1543 : INV_X1 port map( A => d_in(16), ZN => n1070);
   U1544 : NAND4_X1 port map( A1 => n1071, A2 => n1072, A3 => n1073, A4 => 
                           n1074, ZN => n1068);
   U1545 : AOI221_X1 port map( B1 => n760, B2 => registers_11_16_port, C1 => 
                           n761, C2 => registers_14_16_port, A => n1075, ZN => 
                           n1074);
   U1546 : OAI22_X1 port map( A1 => n382, A2 => n758, B1 => n126, B2 => n757, 
                           ZN => n1075);
   U1547 : INV_X1 port map( A => n1076, ZN => n1073);
   U1548 : OAI221_X1 port map( B1 => n752, B2 => n192, C1 => n753, C2 => n508, 
                           A => n1077, ZN => n1076);
   U1549 : AOI22_X1 port map( A1 => registers_6_16_port, A2 => n756, B1 => 
                           registers_3_16_port, B2 => n755, ZN => n1077);
   U1550 : INV_X1 port map( A => n1078, ZN => n1072);
   U1551 : OAI221_X1 port map( B1 => n747, B2 => n191, C1 => n748, C2 => n507, 
                           A => n1079, ZN => n1078);
   U1552 : AOI22_X1 port map( A1 => registers_25_16_port, A2 => n751, B1 => 
                           registers_28_16_port, B2 => n750, ZN => n1079);
   U1553 : AOI221_X1 port map( B1 => n745, B2 => registers_22_16_port, C1 => 
                           n746, C2 => registers_19_16_port, A => n1080, ZN => 
                           n1071);
   U1554 : OAI22_X1 port map( A1 => n381, A2 => n743, B1 => n125, B2 => n742, 
                           ZN => n1080);
   U1555 : OAI21_X1 port map( B1 => n707, B2 => n337, A => n1081, ZN => n3014);
   U1556 : AOI22_X1 port map( A1 => n709, A2 => d_in(15), B1 => d_link(15), B2 
                           => n710, ZN => n1081);
   U1557 : NAND4_X1 port map( A1 => n1082, A2 => n1083, A3 => n1084, A4 => 
                           n1085, ZN => n3013);
   U1558 : AOI221_X1 port map( B1 => n715, B2 => registers_12_15_port, C1 => 
                           n716, C2 => registers_9_15_port, A => n1086, ZN => 
                           n1085);
   U1559 : OAI222_X1 port map( A1 => n447, A2 => n718, B1 => n33, B2 => n719, 
                           C1 => n257, C2 => n720, ZN => n1086);
   U1560 : AOI221_X1 port map( B1 => n721, B2 => registers_4_15_port, C1 => 
                           n722, C2 => registers_20_15_port, A => n1087, ZN => 
                           n1084);
   U1561 : OAI22_X1 port map( A1 => n81, A2 => n724, B1 => n306, B2 => n725, ZN
                           => n1087);
   U1562 : AOI221_X1 port map( B1 => n726, B2 => registers_15_15_port, C1 => 
                           n727, C2 => registers_30_15_port, A => n1088, ZN => 
                           n1083);
   U1563 : OAI222_X1 port map( A1 => n448, A2 => n729, B1 => n34, B2 => n730, 
                           C1 => n258, C2 => n731, ZN => n1088);
   U1564 : AOI221_X1 port map( B1 => registers_31_15_port, B2 => n770, C1 => 
                           n771, C2 => n1089, A => n1090, ZN => n1082);
   U1565 : OAI22_X1 port map( A1 => n2934, A2 => n774, B1 => n1091, B2 => n776,
                           ZN => n1090);
   U1566 : INV_X1 port map( A => d_in(15), ZN => n1091);
   U1567 : NAND4_X1 port map( A1 => n1092, A2 => n1093, A3 => n1094, A4 => 
                           n1095, ZN => n1089);
   U1568 : AOI221_X1 port map( B1 => n760, B2 => registers_11_15_port, C1 => 
                           n761, C2 => registers_14_15_port, A => n1096, ZN => 
                           n1095);
   U1569 : OAI22_X1 port map( A1 => n384, A2 => n758, B1 => n128, B2 => n757, 
                           ZN => n1096);
   U1570 : INV_X1 port map( A => n1097, ZN => n1094);
   U1571 : OAI221_X1 port map( B1 => n752, B2 => n194, C1 => n753, C2 => n510, 
                           A => n1098, ZN => n1097);
   U1572 : AOI22_X1 port map( A1 => registers_6_15_port, A2 => n756, B1 => 
                           registers_3_15_port, B2 => n755, ZN => n1098);
   U1573 : INV_X1 port map( A => n1099, ZN => n1093);
   U1574 : OAI221_X1 port map( B1 => n747, B2 => n193, C1 => n748, C2 => n509, 
                           A => n1100, ZN => n1099);
   U1575 : AOI22_X1 port map( A1 => registers_25_15_port, A2 => n751, B1 => 
                           registers_28_15_port, B2 => n750, ZN => n1100);
   U1576 : AOI221_X1 port map( B1 => n745, B2 => registers_22_15_port, C1 => 
                           n746, C2 => registers_19_15_port, A => n1101, ZN => 
                           n1092);
   U1577 : OAI22_X1 port map( A1 => n383, A2 => n743, B1 => n127, B2 => n742, 
                           ZN => n1101);
   U1578 : OAI21_X1 port map( B1 => n707, B2 => n338, A => n1102, ZN => n3012);
   U1579 : AOI22_X1 port map( A1 => n709, A2 => d_in(14), B1 => d_link(14), B2 
                           => n710, ZN => n1102);
   U1580 : NAND4_X1 port map( A1 => n1103, A2 => n1104, A3 => n1105, A4 => 
                           n1106, ZN => n3011);
   U1581 : AOI221_X1 port map( B1 => n715, B2 => registers_12_14_port, C1 => 
                           n716, C2 => registers_9_14_port, A => n1107, ZN => 
                           n1106);
   U1582 : OAI222_X1 port map( A1 => n449, A2 => n718, B1 => n35, B2 => n719, 
                           C1 => n259, C2 => n720, ZN => n1107);
   U1583 : AOI221_X1 port map( B1 => n721, B2 => registers_4_14_port, C1 => 
                           n722, C2 => registers_20_14_port, A => n1108, ZN => 
                           n1105);
   U1584 : OAI22_X1 port map( A1 => n82, A2 => n724, B1 => n307, B2 => n725, ZN
                           => n1108);
   U1585 : AOI221_X1 port map( B1 => n726, B2 => registers_15_14_port, C1 => 
                           n727, C2 => registers_30_14_port, A => n1109, ZN => 
                           n1104);
   U1586 : OAI222_X1 port map( A1 => n450, A2 => n729, B1 => n36, B2 => n730, 
                           C1 => n260, C2 => n731, ZN => n1109);
   U1587 : AOI221_X1 port map( B1 => registers_31_14_port, B2 => n770, C1 => 
                           n771, C2 => n1110, A => n1111, ZN => n1103);
   U1588 : OAI22_X1 port map( A1 => n2933, A2 => n774, B1 => n1112, B2 => n776,
                           ZN => n1111);
   U1589 : INV_X1 port map( A => d_in(14), ZN => n1112);
   U1590 : NAND4_X1 port map( A1 => n1113, A2 => n1114, A3 => n1115, A4 => 
                           n1116, ZN => n1110);
   U1591 : AOI221_X1 port map( B1 => n760, B2 => registers_11_14_port, C1 => 
                           n761, C2 => registers_14_14_port, A => n1117, ZN => 
                           n1116);
   U1592 : OAI22_X1 port map( A1 => n386, A2 => n758, B1 => n130, B2 => n757, 
                           ZN => n1117);
   U1593 : INV_X1 port map( A => n1118, ZN => n1115);
   U1594 : OAI221_X1 port map( B1 => n752, B2 => n196, C1 => n753, C2 => n512, 
                           A => n1119, ZN => n1118);
   U1595 : AOI22_X1 port map( A1 => registers_6_14_port, A2 => n756, B1 => 
                           registers_3_14_port, B2 => n755, ZN => n1119);
   U1596 : INV_X1 port map( A => n1120, ZN => n1114);
   U1597 : OAI221_X1 port map( B1 => n747, B2 => n195, C1 => n748, C2 => n511, 
                           A => n1121, ZN => n1120);
   U1598 : AOI22_X1 port map( A1 => registers_25_14_port, A2 => n751, B1 => 
                           registers_28_14_port, B2 => n750, ZN => n1121);
   U1599 : AOI221_X1 port map( B1 => n745, B2 => registers_22_14_port, C1 => 
                           n746, C2 => registers_19_14_port, A => n1122, ZN => 
                           n1113);
   U1600 : OAI22_X1 port map( A1 => n385, A2 => n743, B1 => n129, B2 => n742, 
                           ZN => n1122);
   U1601 : OAI21_X1 port map( B1 => n707, B2 => n339, A => n1123, ZN => n3010);
   U1602 : AOI22_X1 port map( A1 => n709, A2 => d_in(13), B1 => d_link(13), B2 
                           => n710, ZN => n1123);
   U1603 : NAND4_X1 port map( A1 => n1124, A2 => n1125, A3 => n1126, A4 => 
                           n1127, ZN => n3009);
   U1604 : AOI221_X1 port map( B1 => n715, B2 => registers_12_13_port, C1 => 
                           n716, C2 => registers_9_13_port, A => n1128, ZN => 
                           n1127);
   U1605 : OAI222_X1 port map( A1 => n451, A2 => n718, B1 => n37, B2 => n719, 
                           C1 => n261, C2 => n720, ZN => n1128);
   U1606 : AOI221_X1 port map( B1 => n721, B2 => registers_4_13_port, C1 => 
                           n722, C2 => registers_20_13_port, A => n1129, ZN => 
                           n1126);
   U1607 : OAI22_X1 port map( A1 => n83, A2 => n724, B1 => n308, B2 => n725, ZN
                           => n1129);
   U1608 : AOI221_X1 port map( B1 => n726, B2 => registers_15_13_port, C1 => 
                           n727, C2 => registers_30_13_port, A => n1130, ZN => 
                           n1125);
   U1609 : OAI222_X1 port map( A1 => n452, A2 => n729, B1 => n38, B2 => n730, 
                           C1 => n262, C2 => n731, ZN => n1130);
   U1610 : AOI221_X1 port map( B1 => registers_31_13_port, B2 => n770, C1 => 
                           n771, C2 => n1131, A => n1132, ZN => n1124);
   U1611 : OAI22_X1 port map( A1 => n2932, A2 => n774, B1 => n1133, B2 => n776,
                           ZN => n1132);
   U1612 : INV_X1 port map( A => d_in(13), ZN => n1133);
   U1613 : NAND4_X1 port map( A1 => n1134, A2 => n1135, A3 => n1136, A4 => 
                           n1137, ZN => n1131);
   U1614 : AOI221_X1 port map( B1 => n760, B2 => registers_11_13_port, C1 => 
                           n761, C2 => registers_14_13_port, A => n1138, ZN => 
                           n1137);
   U1615 : OAI22_X1 port map( A1 => n388, A2 => n758, B1 => n132, B2 => n757, 
                           ZN => n1138);
   U1616 : INV_X1 port map( A => n1139, ZN => n1136);
   U1617 : OAI221_X1 port map( B1 => n752, B2 => n198, C1 => n753, C2 => n514, 
                           A => n1140, ZN => n1139);
   U1618 : AOI22_X1 port map( A1 => registers_6_13_port, A2 => n756, B1 => 
                           registers_3_13_port, B2 => n755, ZN => n1140);
   U1619 : INV_X1 port map( A => n1141, ZN => n1135);
   U1620 : OAI221_X1 port map( B1 => n747, B2 => n197, C1 => n748, C2 => n513, 
                           A => n1142, ZN => n1141);
   U1621 : AOI22_X1 port map( A1 => registers_25_13_port, A2 => n751, B1 => 
                           registers_28_13_port, B2 => n750, ZN => n1142);
   U1622 : AOI221_X1 port map( B1 => n745, B2 => registers_22_13_port, C1 => 
                           n746, C2 => registers_19_13_port, A => n1143, ZN => 
                           n1134);
   U1623 : OAI22_X1 port map( A1 => n387, A2 => n743, B1 => n131, B2 => n742, 
                           ZN => n1143);
   U1624 : OAI21_X1 port map( B1 => n707, B2 => n340, A => n1144, ZN => n3008);
   U1625 : AOI22_X1 port map( A1 => n709, A2 => d_in(12), B1 => d_link(12), B2 
                           => n710, ZN => n1144);
   U1626 : NAND4_X1 port map( A1 => n1145, A2 => n1146, A3 => n1147, A4 => 
                           n1148, ZN => n3007);
   U1627 : AOI221_X1 port map( B1 => n715, B2 => registers_12_12_port, C1 => 
                           n716, C2 => registers_9_12_port, A => n1149, ZN => 
                           n1148);
   U1628 : OAI222_X1 port map( A1 => n453, A2 => n718, B1 => n39, B2 => n719, 
                           C1 => n263, C2 => n720, ZN => n1149);
   U1629 : AOI221_X1 port map( B1 => n721, B2 => registers_4_12_port, C1 => 
                           n722, C2 => registers_20_12_port, A => n1150, ZN => 
                           n1147);
   U1630 : OAI22_X1 port map( A1 => n84, A2 => n724, B1 => n309, B2 => n725, ZN
                           => n1150);
   U1631 : AOI221_X1 port map( B1 => n726, B2 => registers_15_12_port, C1 => 
                           n727, C2 => registers_30_12_port, A => n1151, ZN => 
                           n1146);
   U1632 : OAI222_X1 port map( A1 => n454, A2 => n729, B1 => n40, B2 => n730, 
                           C1 => n264, C2 => n731, ZN => n1151);
   U1633 : AOI221_X1 port map( B1 => registers_31_12_port, B2 => n770, C1 => 
                           n771, C2 => n1152, A => n1153, ZN => n1145);
   U1634 : OAI22_X1 port map( A1 => n2931, A2 => n774, B1 => n1154, B2 => n776,
                           ZN => n1153);
   U1635 : INV_X1 port map( A => d_in(12), ZN => n1154);
   U1636 : NAND4_X1 port map( A1 => n1155, A2 => n1156, A3 => n1157, A4 => 
                           n1158, ZN => n1152);
   U1637 : AOI221_X1 port map( B1 => n760, B2 => registers_11_12_port, C1 => 
                           n761, C2 => registers_14_12_port, A => n1159, ZN => 
                           n1158);
   U1638 : OAI22_X1 port map( A1 => n390, A2 => n758, B1 => n134, B2 => n757, 
                           ZN => n1159);
   U1639 : INV_X1 port map( A => n1160, ZN => n1157);
   U1640 : OAI221_X1 port map( B1 => n752, B2 => n200, C1 => n753, C2 => n516, 
                           A => n1161, ZN => n1160);
   U1641 : AOI22_X1 port map( A1 => registers_6_12_port, A2 => n756, B1 => 
                           registers_3_12_port, B2 => n755, ZN => n1161);
   U1642 : INV_X1 port map( A => n1162, ZN => n1156);
   U1643 : OAI221_X1 port map( B1 => n747, B2 => n199, C1 => n748, C2 => n515, 
                           A => n1163, ZN => n1162);
   U1644 : AOI22_X1 port map( A1 => registers_25_12_port, A2 => n751, B1 => 
                           registers_28_12_port, B2 => n750, ZN => n1163);
   U1645 : AOI221_X1 port map( B1 => n745, B2 => registers_22_12_port, C1 => 
                           n746, C2 => registers_19_12_port, A => n1164, ZN => 
                           n1155);
   U1646 : OAI22_X1 port map( A1 => n389, A2 => n743, B1 => n133, B2 => n742, 
                           ZN => n1164);
   U1647 : OAI21_X1 port map( B1 => n707, B2 => n341, A => n1165, ZN => n3006);
   U1648 : AOI22_X1 port map( A1 => n709, A2 => d_in(11), B1 => d_link(11), B2 
                           => n710, ZN => n1165);
   U1649 : NAND4_X1 port map( A1 => n1166, A2 => n1167, A3 => n1168, A4 => 
                           n1169, ZN => n3005);
   U1650 : AOI221_X1 port map( B1 => n715, B2 => registers_12_11_port, C1 => 
                           n716, C2 => registers_9_11_port, A => n1170, ZN => 
                           n1169);
   U1651 : OAI222_X1 port map( A1 => n455, A2 => n718, B1 => n41, B2 => n719, 
                           C1 => n265, C2 => n720, ZN => n1170);
   U1652 : AOI221_X1 port map( B1 => n721, B2 => registers_4_11_port, C1 => 
                           n722, C2 => registers_20_11_port, A => n1171, ZN => 
                           n1168);
   U1653 : OAI22_X1 port map( A1 => n85, A2 => n724, B1 => n310, B2 => n725, ZN
                           => n1171);
   U1654 : AOI221_X1 port map( B1 => n726, B2 => registers_15_11_port, C1 => 
                           n727, C2 => registers_30_11_port, A => n1172, ZN => 
                           n1167);
   U1655 : OAI222_X1 port map( A1 => n456, A2 => n729, B1 => n42, B2 => n730, 
                           C1 => n266, C2 => n731, ZN => n1172);
   U1656 : AOI221_X1 port map( B1 => registers_31_11_port, B2 => n770, C1 => 
                           n771, C2 => n1173, A => n1174, ZN => n1166);
   U1657 : OAI22_X1 port map( A1 => n2930, A2 => n774, B1 => n1175, B2 => n776,
                           ZN => n1174);
   U1658 : INV_X1 port map( A => d_in(11), ZN => n1175);
   U1659 : NAND4_X1 port map( A1 => n1176, A2 => n1177, A3 => n1178, A4 => 
                           n1179, ZN => n1173);
   U1660 : AOI221_X1 port map( B1 => n760, B2 => registers_11_11_port, C1 => 
                           n761, C2 => registers_14_11_port, A => n1180, ZN => 
                           n1179);
   U1661 : OAI22_X1 port map( A1 => n392, A2 => n758, B1 => n136, B2 => n757, 
                           ZN => n1180);
   U1662 : INV_X1 port map( A => n1181, ZN => n1178);
   U1663 : OAI221_X1 port map( B1 => n752, B2 => n202, C1 => n753, C2 => n518, 
                           A => n1182, ZN => n1181);
   U1664 : AOI22_X1 port map( A1 => registers_6_11_port, A2 => n756, B1 => 
                           registers_3_11_port, B2 => n755, ZN => n1182);
   U1665 : INV_X1 port map( A => n1183, ZN => n1177);
   U1666 : OAI221_X1 port map( B1 => n747, B2 => n201, C1 => n748, C2 => n517, 
                           A => n1184, ZN => n1183);
   U1667 : AOI22_X1 port map( A1 => registers_25_11_port, A2 => n751, B1 => 
                           registers_28_11_port, B2 => n750, ZN => n1184);
   U1668 : AOI221_X1 port map( B1 => n745, B2 => registers_22_11_port, C1 => 
                           n746, C2 => registers_19_11_port, A => n1185, ZN => 
                           n1176);
   U1669 : OAI22_X1 port map( A1 => n391, A2 => n743, B1 => n135, B2 => n742, 
                           ZN => n1185);
   U1670 : OAI21_X1 port map( B1 => n707, B2 => n342, A => n1186, ZN => n3004);
   U1671 : AOI22_X1 port map( A1 => n709, A2 => d_in(10), B1 => d_link(10), B2 
                           => n710, ZN => n1186);
   U1672 : NAND4_X1 port map( A1 => n1187, A2 => n1188, A3 => n1189, A4 => 
                           n1190, ZN => n3003);
   U1673 : AOI221_X1 port map( B1 => n715, B2 => registers_12_10_port, C1 => 
                           n716, C2 => registers_9_10_port, A => n1191, ZN => 
                           n1190);
   U1674 : OAI222_X1 port map( A1 => n457, A2 => n718, B1 => n43, B2 => n719, 
                           C1 => n267, C2 => n720, ZN => n1191);
   U1675 : AOI221_X1 port map( B1 => n721, B2 => registers_4_10_port, C1 => 
                           n722, C2 => registers_20_10_port, A => n1192, ZN => 
                           n1189);
   U1676 : OAI22_X1 port map( A1 => n86, A2 => n724, B1 => n311, B2 => n725, ZN
                           => n1192);
   U1677 : AOI221_X1 port map( B1 => n726, B2 => registers_15_10_port, C1 => 
                           n727, C2 => registers_30_10_port, A => n1193, ZN => 
                           n1188);
   U1678 : OAI222_X1 port map( A1 => n458, A2 => n729, B1 => n44, B2 => n730, 
                           C1 => n268, C2 => n731, ZN => n1193);
   U1679 : AOI221_X1 port map( B1 => registers_31_10_port, B2 => n770, C1 => 
                           n771, C2 => n1194, A => n1195, ZN => n1187);
   U1680 : OAI22_X1 port map( A1 => n2929, A2 => n774, B1 => n1196, B2 => n776,
                           ZN => n1195);
   U1681 : INV_X1 port map( A => d_in(10), ZN => n1196);
   U1682 : NAND4_X1 port map( A1 => n1197, A2 => n1198, A3 => n1199, A4 => 
                           n1200, ZN => n1194);
   U1683 : AOI221_X1 port map( B1 => n760, B2 => registers_11_10_port, C1 => 
                           n761, C2 => registers_14_10_port, A => n1201, ZN => 
                           n1200);
   U1684 : OAI22_X1 port map( A1 => n394, A2 => n758, B1 => n138, B2 => n757, 
                           ZN => n1201);
   U1685 : INV_X1 port map( A => n1202, ZN => n1199);
   U1686 : OAI221_X1 port map( B1 => n752, B2 => n204, C1 => n753, C2 => n520, 
                           A => n1203, ZN => n1202);
   U1687 : AOI22_X1 port map( A1 => registers_6_10_port, A2 => n756, B1 => 
                           registers_3_10_port, B2 => n755, ZN => n1203);
   U1688 : INV_X1 port map( A => n1204, ZN => n1198);
   U1689 : OAI221_X1 port map( B1 => n747, B2 => n203, C1 => n748, C2 => n519, 
                           A => n1205, ZN => n1204);
   U1690 : AOI22_X1 port map( A1 => registers_25_10_port, A2 => n751, B1 => 
                           registers_28_10_port, B2 => n750, ZN => n1205);
   U1691 : AOI221_X1 port map( B1 => n745, B2 => registers_22_10_port, C1 => 
                           n746, C2 => registers_19_10_port, A => n1206, ZN => 
                           n1197);
   U1692 : OAI22_X1 port map( A1 => n393, A2 => n743, B1 => n137, B2 => n742, 
                           ZN => n1206);
   U1693 : OAI21_X1 port map( B1 => n707, B2 => n343, A => n1207, ZN => n3002);
   U1694 : AOI22_X1 port map( A1 => n709, A2 => d_in(9), B1 => d_link(9), B2 =>
                           n710, ZN => n1207);
   U1695 : NAND4_X1 port map( A1 => n1208, A2 => n1209, A3 => n1210, A4 => 
                           n1211, ZN => n3001);
   U1696 : AOI221_X1 port map( B1 => n715, B2 => registers_12_9_port, C1 => 
                           n716, C2 => registers_9_9_port, A => n1212, ZN => 
                           n1211);
   U1697 : OAI222_X1 port map( A1 => n459, A2 => n718, B1 => n45, B2 => n719, 
                           C1 => n269, C2 => n720, ZN => n1212);
   U1698 : AOI221_X1 port map( B1 => n721, B2 => registers_4_9_port, C1 => n722
                           , C2 => registers_20_9_port, A => n1213, ZN => n1210
                           );
   U1699 : OAI22_X1 port map( A1 => n87, A2 => n724, B1 => n312, B2 => n725, ZN
                           => n1213);
   U1700 : AOI221_X1 port map( B1 => n726, B2 => registers_15_9_port, C1 => 
                           n727, C2 => registers_30_9_port, A => n1214, ZN => 
                           n1209);
   U1701 : OAI222_X1 port map( A1 => n460, A2 => n729, B1 => n46, B2 => n730, 
                           C1 => n270, C2 => n731, ZN => n1214);
   U1702 : AOI221_X1 port map( B1 => registers_31_9_port, B2 => n770, C1 => 
                           n771, C2 => n1215, A => n1216, ZN => n1208);
   U1703 : OAI22_X1 port map( A1 => n2928, A2 => n774, B1 => n1217, B2 => n776,
                           ZN => n1216);
   U1704 : INV_X1 port map( A => d_in(9), ZN => n1217);
   U1705 : NAND4_X1 port map( A1 => n1218, A2 => n1219, A3 => n1220, A4 => 
                           n1221, ZN => n1215);
   U1706 : AOI221_X1 port map( B1 => n760, B2 => registers_11_9_port, C1 => 
                           n761, C2 => registers_14_9_port, A => n1222, ZN => 
                           n1221);
   U1707 : OAI22_X1 port map( A1 => n396, A2 => n758, B1 => n140, B2 => n757, 
                           ZN => n1222);
   U1708 : INV_X1 port map( A => n1223, ZN => n1220);
   U1709 : OAI221_X1 port map( B1 => n752, B2 => n206, C1 => n753, C2 => n522, 
                           A => n1224, ZN => n1223);
   U1710 : AOI22_X1 port map( A1 => registers_6_9_port, A2 => n756, B1 => 
                           registers_3_9_port, B2 => n755, ZN => n1224);
   U1711 : INV_X1 port map( A => n1225, ZN => n1219);
   U1712 : OAI221_X1 port map( B1 => n747, B2 => n205, C1 => n748, C2 => n521, 
                           A => n1226, ZN => n1225);
   U1713 : AOI22_X1 port map( A1 => registers_25_9_port, A2 => n751, B1 => 
                           registers_28_9_port, B2 => n750, ZN => n1226);
   U1714 : AOI221_X1 port map( B1 => n745, B2 => registers_22_9_port, C1 => 
                           n746, C2 => registers_19_9_port, A => n1227, ZN => 
                           n1218);
   U1715 : OAI22_X1 port map( A1 => n395, A2 => n743, B1 => n139, B2 => n742, 
                           ZN => n1227);
   U1716 : OAI21_X1 port map( B1 => n707, B2 => n344, A => n1228, ZN => n3000);
   U1717 : AOI22_X1 port map( A1 => n709, A2 => d_in(8), B1 => d_link(8), B2 =>
                           n710, ZN => n1228);
   U1718 : NAND4_X1 port map( A1 => n1229, A2 => n1230, A3 => n1231, A4 => 
                           n1232, ZN => n2999);
   U1719 : AOI221_X1 port map( B1 => n715, B2 => registers_12_8_port, C1 => 
                           n716, C2 => registers_9_8_port, A => n1233, ZN => 
                           n1232);
   U1720 : OAI222_X1 port map( A1 => n461, A2 => n718, B1 => n47, B2 => n719, 
                           C1 => n271, C2 => n720, ZN => n1233);
   U1721 : AOI221_X1 port map( B1 => n721, B2 => registers_4_8_port, C1 => n722
                           , C2 => registers_20_8_port, A => n1234, ZN => n1231
                           );
   U1722 : OAI22_X1 port map( A1 => n88, A2 => n724, B1 => n313, B2 => n725, ZN
                           => n1234);
   U1723 : AOI221_X1 port map( B1 => n726, B2 => registers_15_8_port, C1 => 
                           n727, C2 => registers_30_8_port, A => n1235, ZN => 
                           n1230);
   U1724 : OAI222_X1 port map( A1 => n462, A2 => n729, B1 => n48, B2 => n730, 
                           C1 => n272, C2 => n731, ZN => n1235);
   U1725 : AOI221_X1 port map( B1 => registers_31_8_port, B2 => n770, C1 => 
                           n771, C2 => n1236, A => n1237, ZN => n1229);
   U1726 : OAI22_X1 port map( A1 => n2927, A2 => n774, B1 => n1238, B2 => n776,
                           ZN => n1237);
   U1727 : INV_X1 port map( A => d_in(8), ZN => n1238);
   U1728 : NAND4_X1 port map( A1 => n1239, A2 => n1240, A3 => n1241, A4 => 
                           n1242, ZN => n1236);
   U1729 : AOI221_X1 port map( B1 => n760, B2 => registers_11_8_port, C1 => 
                           n761, C2 => registers_14_8_port, A => n1243, ZN => 
                           n1242);
   U1730 : OAI22_X1 port map( A1 => n398, A2 => n758, B1 => n142, B2 => n757, 
                           ZN => n1243);
   U1731 : INV_X1 port map( A => n1244, ZN => n1241);
   U1732 : OAI221_X1 port map( B1 => n752, B2 => n208, C1 => n753, C2 => n524, 
                           A => n1245, ZN => n1244);
   U1733 : AOI22_X1 port map( A1 => registers_6_8_port, A2 => n756, B1 => 
                           registers_3_8_port, B2 => n755, ZN => n1245);
   U1734 : INV_X1 port map( A => n1246, ZN => n1240);
   U1735 : OAI221_X1 port map( B1 => n747, B2 => n207, C1 => n748, C2 => n523, 
                           A => n1247, ZN => n1246);
   U1736 : AOI22_X1 port map( A1 => registers_25_8_port, A2 => n751, B1 => 
                           registers_28_8_port, B2 => n750, ZN => n1247);
   U1737 : AOI221_X1 port map( B1 => n745, B2 => registers_22_8_port, C1 => 
                           n746, C2 => registers_19_8_port, A => n1248, ZN => 
                           n1239);
   U1738 : OAI22_X1 port map( A1 => n397, A2 => n743, B1 => n141, B2 => n742, 
                           ZN => n1248);
   U1739 : OAI21_X1 port map( B1 => n707, B2 => n345, A => n1249, ZN => n2998);
   U1740 : AOI22_X1 port map( A1 => n709, A2 => d_in(7), B1 => d_link(7), B2 =>
                           n710, ZN => n1249);
   U1741 : NAND4_X1 port map( A1 => n1250, A2 => n1251, A3 => n1252, A4 => 
                           n1253, ZN => n2997);
   U1742 : AOI221_X1 port map( B1 => n715, B2 => registers_12_7_port, C1 => 
                           n716, C2 => registers_9_7_port, A => n1254, ZN => 
                           n1253);
   U1743 : OAI222_X1 port map( A1 => n463, A2 => n718, B1 => n49, B2 => n719, 
                           C1 => n273, C2 => n720, ZN => n1254);
   U1744 : AOI221_X1 port map( B1 => n721, B2 => registers_4_7_port, C1 => n722
                           , C2 => registers_20_7_port, A => n1255, ZN => n1252
                           );
   U1745 : OAI22_X1 port map( A1 => n89, A2 => n724, B1 => n314, B2 => n725, ZN
                           => n1255);
   U1746 : AOI221_X1 port map( B1 => n726, B2 => registers_15_7_port, C1 => 
                           n727, C2 => registers_30_7_port, A => n1256, ZN => 
                           n1251);
   U1747 : OAI222_X1 port map( A1 => n464, A2 => n729, B1 => n50, B2 => n730, 
                           C1 => n274, C2 => n731, ZN => n1256);
   U1748 : AOI221_X1 port map( B1 => registers_31_7_port, B2 => n770, C1 => 
                           n771, C2 => n1257, A => n1258, ZN => n1250);
   U1749 : OAI22_X1 port map( A1 => n2926, A2 => n774, B1 => n1259, B2 => n776,
                           ZN => n1258);
   U1750 : INV_X1 port map( A => d_in(7), ZN => n1259);
   U1751 : NAND4_X1 port map( A1 => n1260, A2 => n1261, A3 => n1262, A4 => 
                           n1263, ZN => n1257);
   U1752 : AOI221_X1 port map( B1 => n760, B2 => registers_11_7_port, C1 => 
                           n761, C2 => registers_14_7_port, A => n1264, ZN => 
                           n1263);
   U1753 : OAI22_X1 port map( A1 => n400, A2 => n758, B1 => n144, B2 => n757, 
                           ZN => n1264);
   U1754 : INV_X1 port map( A => n1265, ZN => n1262);
   U1755 : OAI221_X1 port map( B1 => n752, B2 => n210, C1 => n753, C2 => n526, 
                           A => n1266, ZN => n1265);
   U1756 : AOI22_X1 port map( A1 => registers_6_7_port, A2 => n756, B1 => 
                           registers_3_7_port, B2 => n755, ZN => n1266);
   U1757 : INV_X1 port map( A => n1267, ZN => n1261);
   U1758 : OAI221_X1 port map( B1 => n747, B2 => n209, C1 => n748, C2 => n525, 
                           A => n1268, ZN => n1267);
   U1759 : AOI22_X1 port map( A1 => registers_25_7_port, A2 => n751, B1 => 
                           registers_28_7_port, B2 => n750, ZN => n1268);
   U1760 : AOI221_X1 port map( B1 => n745, B2 => registers_22_7_port, C1 => 
                           n746, C2 => registers_19_7_port, A => n1269, ZN => 
                           n1260);
   U1761 : OAI22_X1 port map( A1 => n399, A2 => n743, B1 => n143, B2 => n742, 
                           ZN => n1269);
   U1762 : OAI21_X1 port map( B1 => n707, B2 => n346, A => n1270, ZN => n2996);
   U1763 : AOI22_X1 port map( A1 => n709, A2 => d_in(6), B1 => d_link(6), B2 =>
                           n710, ZN => n1270);
   U1764 : NAND4_X1 port map( A1 => n1271, A2 => n1272, A3 => n1273, A4 => 
                           n1274, ZN => n2995);
   U1765 : AOI221_X1 port map( B1 => n715, B2 => registers_12_6_port, C1 => 
                           n716, C2 => registers_9_6_port, A => n1275, ZN => 
                           n1274);
   U1766 : OAI222_X1 port map( A1 => n465, A2 => n718, B1 => n51, B2 => n719, 
                           C1 => n275, C2 => n720, ZN => n1275);
   U1767 : AOI221_X1 port map( B1 => n721, B2 => registers_4_6_port, C1 => n722
                           , C2 => registers_20_6_port, A => n1276, ZN => n1273
                           );
   U1768 : OAI22_X1 port map( A1 => n90, A2 => n724, B1 => n315, B2 => n725, ZN
                           => n1276);
   U1769 : AOI221_X1 port map( B1 => n726, B2 => registers_15_6_port, C1 => 
                           n727, C2 => registers_30_6_port, A => n1277, ZN => 
                           n1272);
   U1770 : OAI222_X1 port map( A1 => n466, A2 => n729, B1 => n52, B2 => n730, 
                           C1 => n276, C2 => n731, ZN => n1277);
   U1771 : AOI221_X1 port map( B1 => registers_31_6_port, B2 => n770, C1 => 
                           n771, C2 => n1278, A => n1279, ZN => n1271);
   U1772 : OAI22_X1 port map( A1 => n2925, A2 => n774, B1 => n1280, B2 => n776,
                           ZN => n1279);
   U1773 : INV_X1 port map( A => d_in(6), ZN => n1280);
   U1774 : NAND4_X1 port map( A1 => n1281, A2 => n1282, A3 => n1283, A4 => 
                           n1284, ZN => n1278);
   U1775 : AOI221_X1 port map( B1 => n760, B2 => registers_11_6_port, C1 => 
                           n761, C2 => registers_14_6_port, A => n1285, ZN => 
                           n1284);
   U1776 : OAI22_X1 port map( A1 => n402, A2 => n758, B1 => n146, B2 => n757, 
                           ZN => n1285);
   U1777 : INV_X1 port map( A => n1286, ZN => n1283);
   U1778 : OAI221_X1 port map( B1 => n752, B2 => n212, C1 => n753, C2 => n528, 
                           A => n1287, ZN => n1286);
   U1779 : AOI22_X1 port map( A1 => registers_6_6_port, A2 => n756, B1 => 
                           registers_3_6_port, B2 => n755, ZN => n1287);
   U1780 : INV_X1 port map( A => n1288, ZN => n1282);
   U1781 : OAI221_X1 port map( B1 => n747, B2 => n211, C1 => n748, C2 => n527, 
                           A => n1289, ZN => n1288);
   U1782 : AOI22_X1 port map( A1 => registers_25_6_port, A2 => n751, B1 => 
                           registers_28_6_port, B2 => n750, ZN => n1289);
   U1783 : AOI221_X1 port map( B1 => n745, B2 => registers_22_6_port, C1 => 
                           n746, C2 => registers_19_6_port, A => n1290, ZN => 
                           n1281);
   U1784 : OAI22_X1 port map( A1 => n401, A2 => n743, B1 => n145, B2 => n742, 
                           ZN => n1290);
   U1785 : OAI21_X1 port map( B1 => n707, B2 => n347, A => n1291, ZN => n2994);
   U1786 : AOI22_X1 port map( A1 => n709, A2 => d_in(5), B1 => d_link(5), B2 =>
                           n710, ZN => n1291);
   U1787 : NAND4_X1 port map( A1 => n1292, A2 => n1293, A3 => n1294, A4 => 
                           n1295, ZN => n2993);
   U1788 : AOI221_X1 port map( B1 => n715, B2 => registers_12_5_port, C1 => 
                           n716, C2 => registers_9_5_port, A => n1296, ZN => 
                           n1295);
   U1789 : OAI222_X1 port map( A1 => n467, A2 => n718, B1 => n53, B2 => n719, 
                           C1 => n277, C2 => n720, ZN => n1296);
   U1790 : AOI221_X1 port map( B1 => n721, B2 => registers_4_5_port, C1 => n722
                           , C2 => registers_20_5_port, A => n1297, ZN => n1294
                           );
   U1791 : OAI22_X1 port map( A1 => n91, A2 => n724, B1 => n316, B2 => n725, ZN
                           => n1297);
   U1792 : AOI221_X1 port map( B1 => n726, B2 => registers_15_5_port, C1 => 
                           n727, C2 => registers_30_5_port, A => n1298, ZN => 
                           n1293);
   U1793 : OAI222_X1 port map( A1 => n468, A2 => n729, B1 => n54, B2 => n730, 
                           C1 => n278, C2 => n731, ZN => n1298);
   U1794 : AOI221_X1 port map( B1 => registers_31_5_port, B2 => n770, C1 => 
                           n771, C2 => n1299, A => n1300, ZN => n1292);
   U1795 : OAI22_X1 port map( A1 => n2924, A2 => n774, B1 => n1301, B2 => n776,
                           ZN => n1300);
   U1796 : INV_X1 port map( A => d_in(5), ZN => n1301);
   U1797 : NAND4_X1 port map( A1 => n1302, A2 => n1303, A3 => n1304, A4 => 
                           n1305, ZN => n1299);
   U1798 : AOI221_X1 port map( B1 => n760, B2 => registers_11_5_port, C1 => 
                           n761, C2 => registers_14_5_port, A => n1306, ZN => 
                           n1305);
   U1799 : OAI22_X1 port map( A1 => n404, A2 => n758, B1 => n148, B2 => n757, 
                           ZN => n1306);
   U1800 : INV_X1 port map( A => n1307, ZN => n1304);
   U1801 : OAI221_X1 port map( B1 => n752, B2 => n214, C1 => n753, C2 => n530, 
                           A => n1308, ZN => n1307);
   U1802 : AOI22_X1 port map( A1 => registers_6_5_port, A2 => n756, B1 => 
                           registers_3_5_port, B2 => n755, ZN => n1308);
   U1803 : INV_X1 port map( A => n1309, ZN => n1303);
   U1804 : OAI221_X1 port map( B1 => n747, B2 => n213, C1 => n748, C2 => n529, 
                           A => n1310, ZN => n1309);
   U1805 : AOI22_X1 port map( A1 => registers_25_5_port, A2 => n751, B1 => 
                           registers_28_5_port, B2 => n750, ZN => n1310);
   U1806 : AOI221_X1 port map( B1 => n745, B2 => registers_22_5_port, C1 => 
                           n746, C2 => registers_19_5_port, A => n1311, ZN => 
                           n1302);
   U1807 : OAI22_X1 port map( A1 => n403, A2 => n743, B1 => n147, B2 => n742, 
                           ZN => n1311);
   U1808 : OAI21_X1 port map( B1 => n707, B2 => n348, A => n1312, ZN => n2992);
   U1809 : AOI22_X1 port map( A1 => n709, A2 => d_in(4), B1 => d_link(4), B2 =>
                           n710, ZN => n1312);
   U1810 : NAND4_X1 port map( A1 => n1313, A2 => n1314, A3 => n1315, A4 => 
                           n1316, ZN => n2991);
   U1811 : AOI221_X1 port map( B1 => n715, B2 => registers_12_4_port, C1 => 
                           n716, C2 => registers_9_4_port, A => n1317, ZN => 
                           n1316);
   U1812 : OAI222_X1 port map( A1 => n469, A2 => n718, B1 => n55, B2 => n719, 
                           C1 => n279, C2 => n720, ZN => n1317);
   U1813 : AOI221_X1 port map( B1 => n721, B2 => registers_4_4_port, C1 => n722
                           , C2 => registers_20_4_port, A => n1318, ZN => n1315
                           );
   U1814 : OAI22_X1 port map( A1 => n92, A2 => n724, B1 => n317, B2 => n725, ZN
                           => n1318);
   U1815 : AOI221_X1 port map( B1 => n726, B2 => registers_15_4_port, C1 => 
                           n727, C2 => registers_30_4_port, A => n1319, ZN => 
                           n1314);
   U1816 : OAI222_X1 port map( A1 => n470, A2 => n729, B1 => n56, B2 => n730, 
                           C1 => n280, C2 => n731, ZN => n1319);
   U1817 : AOI221_X1 port map( B1 => registers_31_4_port, B2 => n770, C1 => 
                           n771, C2 => n1320, A => n1321, ZN => n1313);
   U1818 : OAI22_X1 port map( A1 => n2923, A2 => n774, B1 => n1322, B2 => n776,
                           ZN => n1321);
   U1819 : INV_X1 port map( A => d_in(4), ZN => n1322);
   U1820 : NAND4_X1 port map( A1 => n1323, A2 => n1324, A3 => n1325, A4 => 
                           n1326, ZN => n1320);
   U1821 : AOI221_X1 port map( B1 => n760, B2 => registers_11_4_port, C1 => 
                           n761, C2 => registers_14_4_port, A => n1327, ZN => 
                           n1326);
   U1822 : OAI22_X1 port map( A1 => n406, A2 => n758, B1 => n150, B2 => n757, 
                           ZN => n1327);
   U1823 : INV_X1 port map( A => n1328, ZN => n1325);
   U1824 : OAI221_X1 port map( B1 => n752, B2 => n216, C1 => n753, C2 => n532, 
                           A => n1329, ZN => n1328);
   U1825 : AOI22_X1 port map( A1 => registers_6_4_port, A2 => n756, B1 => 
                           registers_3_4_port, B2 => n755, ZN => n1329);
   U1826 : INV_X1 port map( A => n1330, ZN => n1324);
   U1827 : OAI221_X1 port map( B1 => n747, B2 => n215, C1 => n748, C2 => n531, 
                           A => n1331, ZN => n1330);
   U1828 : AOI22_X1 port map( A1 => registers_25_4_port, A2 => n751, B1 => 
                           registers_28_4_port, B2 => n750, ZN => n1331);
   U1829 : AOI221_X1 port map( B1 => n745, B2 => registers_22_4_port, C1 => 
                           n746, C2 => registers_19_4_port, A => n1332, ZN => 
                           n1323);
   U1830 : OAI22_X1 port map( A1 => n405, A2 => n743, B1 => n149, B2 => n742, 
                           ZN => n1332);
   U1831 : OAI21_X1 port map( B1 => n707, B2 => n349, A => n1333, ZN => n2990);
   U1832 : AOI22_X1 port map( A1 => n709, A2 => d_in(3), B1 => d_link(3), B2 =>
                           n710, ZN => n1333);
   U1833 : NAND4_X1 port map( A1 => n1334, A2 => n1335, A3 => n1336, A4 => 
                           n1337, ZN => n2989);
   U1834 : AOI221_X1 port map( B1 => n715, B2 => registers_12_3_port, C1 => 
                           n716, C2 => registers_9_3_port, A => n1338, ZN => 
                           n1337);
   U1835 : OAI222_X1 port map( A1 => n471, A2 => n718, B1 => n57, B2 => n719, 
                           C1 => n281, C2 => n720, ZN => n1338);
   U1836 : AOI221_X1 port map( B1 => n721, B2 => registers_4_3_port, C1 => n722
                           , C2 => registers_20_3_port, A => n1339, ZN => n1336
                           );
   U1837 : OAI22_X1 port map( A1 => n93, A2 => n724, B1 => n318, B2 => n725, ZN
                           => n1339);
   U1838 : AOI221_X1 port map( B1 => n726, B2 => registers_15_3_port, C1 => 
                           n727, C2 => registers_30_3_port, A => n1340, ZN => 
                           n1335);
   U1839 : OAI222_X1 port map( A1 => n472, A2 => n729, B1 => n58, B2 => n730, 
                           C1 => n282, C2 => n731, ZN => n1340);
   U1840 : AOI221_X1 port map( B1 => registers_31_3_port, B2 => n770, C1 => 
                           n771, C2 => n1341, A => n1342, ZN => n1334);
   U1841 : OAI22_X1 port map( A1 => n2922, A2 => n774, B1 => n1343, B2 => n776,
                           ZN => n1342);
   U1842 : INV_X1 port map( A => d_in(3), ZN => n1343);
   U1843 : NAND4_X1 port map( A1 => n1344, A2 => n1345, A3 => n1346, A4 => 
                           n1347, ZN => n1341);
   U1844 : AOI221_X1 port map( B1 => n760, B2 => registers_11_3_port, C1 => 
                           n761, C2 => registers_14_3_port, A => n1348, ZN => 
                           n1347);
   U1845 : OAI22_X1 port map( A1 => n408, A2 => n758, B1 => n152, B2 => n757, 
                           ZN => n1348);
   U1846 : INV_X1 port map( A => n1349, ZN => n1346);
   U1847 : OAI221_X1 port map( B1 => n752, B2 => n218, C1 => n753, C2 => n534, 
                           A => n1350, ZN => n1349);
   U1848 : AOI22_X1 port map( A1 => registers_6_3_port, A2 => n756, B1 => 
                           registers_3_3_port, B2 => n755, ZN => n1350);
   U1849 : INV_X1 port map( A => n1351, ZN => n1345);
   U1850 : OAI221_X1 port map( B1 => n747, B2 => n217, C1 => n748, C2 => n533, 
                           A => n1352, ZN => n1351);
   U1851 : AOI22_X1 port map( A1 => registers_25_3_port, A2 => n751, B1 => 
                           registers_28_3_port, B2 => n750, ZN => n1352);
   U1852 : AOI221_X1 port map( B1 => n745, B2 => registers_22_3_port, C1 => 
                           n746, C2 => registers_19_3_port, A => n1353, ZN => 
                           n1344);
   U1853 : OAI22_X1 port map( A1 => n407, A2 => n743, B1 => n151, B2 => n742, 
                           ZN => n1353);
   U1854 : OAI21_X1 port map( B1 => n707, B2 => n350, A => n1354, ZN => n2988);
   U1855 : AOI22_X1 port map( A1 => n709, A2 => d_in(2), B1 => d_link(2), B2 =>
                           n710, ZN => n1354);
   U1856 : NAND4_X1 port map( A1 => n1355, A2 => n1356, A3 => n1357, A4 => 
                           n1358, ZN => n2987);
   U1857 : AOI221_X1 port map( B1 => n715, B2 => registers_12_2_port, C1 => 
                           n716, C2 => registers_9_2_port, A => n1359, ZN => 
                           n1358);
   U1858 : OAI222_X1 port map( A1 => n473, A2 => n718, B1 => n59, B2 => n719, 
                           C1 => n283, C2 => n720, ZN => n1359);
   U1859 : AOI221_X1 port map( B1 => n721, B2 => registers_4_2_port, C1 => n722
                           , C2 => registers_20_2_port, A => n1360, ZN => n1357
                           );
   U1860 : OAI22_X1 port map( A1 => n94, A2 => n724, B1 => n319, B2 => n725, ZN
                           => n1360);
   U1861 : AOI221_X1 port map( B1 => n726, B2 => registers_15_2_port, C1 => 
                           n727, C2 => registers_30_2_port, A => n1361, ZN => 
                           n1356);
   U1862 : OAI222_X1 port map( A1 => n474, A2 => n729, B1 => n60, B2 => n730, 
                           C1 => n284, C2 => n731, ZN => n1361);
   U1863 : AOI221_X1 port map( B1 => registers_31_2_port, B2 => n770, C1 => 
                           n771, C2 => n1362, A => n1363, ZN => n1355);
   U1864 : OAI22_X1 port map( A1 => n2921, A2 => n774, B1 => n1364, B2 => n776,
                           ZN => n1363);
   U1865 : INV_X1 port map( A => d_in(2), ZN => n1364);
   U1866 : NAND4_X1 port map( A1 => n1365, A2 => n1366, A3 => n1367, A4 => 
                           n1368, ZN => n1362);
   U1867 : AOI221_X1 port map( B1 => n760, B2 => registers_11_2_port, C1 => 
                           n761, C2 => registers_14_2_port, A => n1369, ZN => 
                           n1368);
   U1868 : OAI22_X1 port map( A1 => n410, A2 => n758, B1 => n154, B2 => n757, 
                           ZN => n1369);
   U1869 : INV_X1 port map( A => n1370, ZN => n1367);
   U1870 : OAI221_X1 port map( B1 => n752, B2 => n220, C1 => n753, C2 => n536, 
                           A => n1371, ZN => n1370);
   U1871 : AOI22_X1 port map( A1 => registers_6_2_port, A2 => n756, B1 => 
                           registers_3_2_port, B2 => n755, ZN => n1371);
   U1872 : INV_X1 port map( A => n1372, ZN => n1366);
   U1873 : OAI221_X1 port map( B1 => n747, B2 => n219, C1 => n748, C2 => n535, 
                           A => n1373, ZN => n1372);
   U1874 : AOI22_X1 port map( A1 => registers_25_2_port, A2 => n751, B1 => 
                           registers_28_2_port, B2 => n750, ZN => n1373);
   U1875 : AOI221_X1 port map( B1 => n745, B2 => registers_22_2_port, C1 => 
                           n746, C2 => registers_19_2_port, A => n1374, ZN => 
                           n1365);
   U1876 : OAI22_X1 port map( A1 => n409, A2 => n743, B1 => n153, B2 => n742, 
                           ZN => n1374);
   U1877 : OAI21_X1 port map( B1 => n707, B2 => n351, A => n1375, ZN => n2986);
   U1878 : AOI22_X1 port map( A1 => n709, A2 => d_in(1), B1 => d_link(1), B2 =>
                           n710, ZN => n1375);
   U1879 : NAND4_X1 port map( A1 => n1376, A2 => n1377, A3 => n1378, A4 => 
                           n1379, ZN => n2985);
   U1880 : AOI221_X1 port map( B1 => n715, B2 => registers_12_1_port, C1 => 
                           n716, C2 => registers_9_1_port, A => n1380, ZN => 
                           n1379);
   U1881 : OAI222_X1 port map( A1 => n475, A2 => n718, B1 => n61, B2 => n719, 
                           C1 => n285, C2 => n720, ZN => n1380);
   U1882 : AOI221_X1 port map( B1 => n721, B2 => registers_4_1_port, C1 => n722
                           , C2 => registers_20_1_port, A => n1381, ZN => n1378
                           );
   U1883 : OAI22_X1 port map( A1 => n95, A2 => n724, B1 => n320, B2 => n725, ZN
                           => n1381);
   U1884 : AOI221_X1 port map( B1 => n726, B2 => registers_15_1_port, C1 => 
                           n727, C2 => registers_30_1_port, A => n1382, ZN => 
                           n1377);
   U1885 : OAI222_X1 port map( A1 => n476, A2 => n729, B1 => n62, B2 => n730, 
                           C1 => n286, C2 => n731, ZN => n1382);
   U1886 : AOI221_X1 port map( B1 => registers_31_1_port, B2 => n770, C1 => 
                           n771, C2 => n1383, A => n1384, ZN => n1376);
   U1887 : OAI22_X1 port map( A1 => n2920, A2 => n774, B1 => n1385, B2 => n776,
                           ZN => n1384);
   U1888 : INV_X1 port map( A => d_in(1), ZN => n1385);
   U1889 : NAND4_X1 port map( A1 => n1386, A2 => n1387, A3 => n1388, A4 => 
                           n1389, ZN => n1383);
   U1890 : AOI221_X1 port map( B1 => n760, B2 => registers_11_1_port, C1 => 
                           n761, C2 => registers_14_1_port, A => n1390, ZN => 
                           n1389);
   U1891 : OAI22_X1 port map( A1 => n412, A2 => n758, B1 => n156, B2 => n757, 
                           ZN => n1390);
   U1892 : INV_X1 port map( A => n1391, ZN => n1388);
   U1893 : OAI221_X1 port map( B1 => n752, B2 => n222, C1 => n753, C2 => n538, 
                           A => n1392, ZN => n1391);
   U1894 : AOI22_X1 port map( A1 => registers_6_1_port, A2 => n756, B1 => 
                           registers_3_1_port, B2 => n755, ZN => n1392);
   U1895 : INV_X1 port map( A => n1393, ZN => n1387);
   U1896 : OAI221_X1 port map( B1 => n747, B2 => n221, C1 => n748, C2 => n537, 
                           A => n1394, ZN => n1393);
   U1897 : AOI22_X1 port map( A1 => registers_25_1_port, A2 => n751, B1 => 
                           registers_28_1_port, B2 => n750, ZN => n1394);
   U1898 : AOI221_X1 port map( B1 => n745, B2 => registers_22_1_port, C1 => 
                           n746, C2 => registers_19_1_port, A => n1395, ZN => 
                           n1386);
   U1899 : OAI22_X1 port map( A1 => n411, A2 => n743, B1 => n155, B2 => n742, 
                           ZN => n1395);
   U1900 : OAI21_X1 port map( B1 => n707, B2 => n352, A => n1396, ZN => n2984);
   U1901 : AOI22_X1 port map( A1 => n709, A2 => d_in(0), B1 => d_link(0), B2 =>
                           n710, ZN => n1396);
   U1902 : AOI22_X1 port map( A1 => en, A2 => link_en, B1 => n663, B2 => n702, 
                           ZN => n1397);
   U1903 : AND3_X1 port map( A1 => wr_addr(3), A2 => wr_addr(2), A3 => n690, ZN
                           => n702);
   U1904 : AND3_X1 port map( A1 => wr_en, A2 => en, A3 => wr_addr(4), ZN => 
                           n690);
   U1905 : NOR2_X1 port map( A1 => n706, A2 => n704, ZN => n663);
   U1906 : INV_X1 port map( A => wr_addr(0), ZN => n704);
   U1907 : INV_X1 port map( A => wr_addr(1), ZN => n706);
   U1908 : NAND4_X1 port map( A1 => n1398, A2 => n1399, A3 => n1400, A4 => 
                           n1401, ZN => n2983);
   U1909 : AOI221_X1 port map( B1 => n715, B2 => registers_12_0_port, C1 => 
                           n716, C2 => registers_9_0_port, A => n1402, ZN => 
                           n1401);
   U1910 : OAI222_X1 port map( A1 => n477, A2 => n718, B1 => n63, B2 => n719, 
                           C1 => n287, C2 => n720, ZN => n1402);
   U1911 : AOI221_X1 port map( B1 => n721, B2 => registers_4_0_port, C1 => n722
                           , C2 => registers_20_0_port, A => n1409, ZN => n1400
                           );
   U1912 : OAI22_X1 port map( A1 => n96, A2 => n724, B1 => n321, B2 => n725, ZN
                           => n1409);
   U1913 : AND2_X1 port map( A1 => n1411, A2 => n771, ZN => n1404);
   U1914 : AOI221_X1 port map( B1 => n726, B2 => registers_15_0_port, C1 => 
                           n727, C2 => registers_30_0_port, A => n1413, ZN => 
                           n1399);
   U1915 : OAI222_X1 port map( A1 => n478, A2 => n729, B1 => n64, B2 => n730, 
                           C1 => n288, C2 => n731, ZN => n1413);
   U1916 : AND2_X1 port map( A1 => n1414, A2 => n771, ZN => n1407);
   U1917 : AOI221_X1 port map( B1 => registers_31_0_port, B2 => n770, C1 => 
                           n771, C2 => n1419, A => n1420, ZN => n1398);
   U1918 : OAI22_X1 port map( A1 => n2919, A2 => n774, B1 => n1421, B2 => n776,
                           ZN => n1420);
   U1919 : NOR2_X1 port map( A1 => n1422, A2 => n733, ZN => n732);
   U1920 : INV_X1 port map( A => d_in(0), ZN => n1421);
   U1921 : NAND4_X1 port map( A1 => n1423, A2 => n1424, A3 => n1425, A4 => 
                           n1426, ZN => n1419);
   U1922 : AOI221_X1 port map( B1 => n760, B2 => registers_11_0_port, C1 => 
                           n761, C2 => registers_14_0_port, A => n1427, ZN => 
                           n1426);
   U1923 : OAI22_X1 port map( A1 => n414, A2 => n758, B1 => n158, B2 => n757, 
                           ZN => n1427);
   U1924 : NOR3_X1 port map( A1 => rd2_addr(0), A2 => rd2_addr(4), A3 => n1428,
                           ZN => n1408);
   U1925 : NOR3_X1 port map( A1 => n1429, A2 => rd2_addr(4), A3 => n1428, ZN =>
                           n1406);
   U1926 : INV_X1 port map( A => n1430, ZN => n1425);
   U1927 : OAI221_X1 port map( B1 => n752, B2 => n224, C1 => n753, C2 => n540, 
                           A => n1431, ZN => n1430);
   U1928 : AOI22_X1 port map( A1 => registers_6_0_port, A2 => n756, B1 => 
                           registers_3_0_port, B2 => n755, ZN => n1431);
   U1929 : NOR3_X1 port map( A1 => rd2_addr(3), A2 => rd2_addr(4), A3 => 
                           rd2_addr(0), ZN => n1412);
   U1930 : INV_X1 port map( A => n1432, ZN => n1424);
   U1931 : OAI221_X1 port map( B1 => n747, B2 => n223, C1 => n748, C2 => n539, 
                           A => n1433, ZN => n1432);
   U1932 : AOI22_X1 port map( A1 => registers_25_0_port, A2 => n751, B1 => 
                           registers_28_0_port, B2 => n750, ZN => n1433);
   U1933 : NOR2_X1 port map( A1 => n1434, A2 => rd2_addr(1), ZN => n1414);
   U1934 : NOR3_X1 port map( A1 => n1435, A2 => rd2_addr(0), A3 => n1428, ZN =>
                           n1415);
   U1935 : AOI221_X1 port map( B1 => n745, B2 => registers_22_0_port, C1 => 
                           n746, C2 => registers_19_0_port, A => n1436, ZN => 
                           n1423);
   U1936 : OAI22_X1 port map( A1 => n413, A2 => n743, B1 => n157, B2 => n742, 
                           ZN => n1436);
   U1937 : NOR2_X1 port map( A1 => rd2_addr(1), A2 => rd2_addr(2), ZN => n1411)
                           ;
   U1938 : NOR3_X1 port map( A1 => rd2_addr(3), A2 => rd2_addr(4), A3 => n1429,
                           ZN => n1410);
   U1939 : NOR3_X1 port map( A1 => n1429, A2 => rd2_addr(3), A3 => n1435, ZN =>
                           n1405);
   U1940 : NOR2_X1 port map( A1 => n1437, A2 => rd2_addr(2), ZN => n1416);
   U1941 : NOR3_X1 port map( A1 => rd2_addr(0), A2 => rd2_addr(3), A3 => n1435,
                           ZN => n1403);
   U1942 : NAND3_X1 port map( A1 => n1417, A2 => n771, A3 => n1418, ZN => n737)
                           ;
   U1943 : NOR2_X1 port map( A1 => n1434, A2 => n1437, ZN => n1418);
   U1944 : INV_X1 port map( A => rd2_addr(1), ZN => n1437);
   U1945 : NAND2_X1 port map( A1 => n774, A2 => n1422, ZN => n736);
   U1946 : NAND4_X1 port map( A1 => n1438, A2 => n1439, A3 => n1440, A4 => 
                           n1441, ZN => n1422);
   U1947 : NOR3_X1 port map( A1 => n1442, A2 => n684, A3 => n1443, ZN => n1441)
                           ;
   U1948 : XOR2_X1 port map( A => wr_addr(1), B => rd2_addr(1), Z => n1443);
   U1949 : XOR2_X1 port map( A => wr_addr(0), B => rd2_addr(0), Z => n1442);
   U1950 : XOR2_X1 port map( A => n1428, B => wr_addr(3), Z => n1440);
   U1951 : XOR2_X1 port map( A => wr_addr(4), B => n1435, Z => n1439);
   U1952 : XOR2_X1 port map( A => n1434, B => wr_addr(2), Z => n1438);
   U1953 : INV_X1 port map( A => rd2_addr(2), ZN => n1434);
   U1954 : NAND3_X1 port map( A1 => rd2_en, A2 => en, A3 => rst, ZN => n733);
   U1955 : NOR3_X1 port map( A1 => n1435, A2 => n1429, A3 => n1428, ZN => n1417
                           );
   U1956 : INV_X1 port map( A => rd2_addr(3), ZN => n1428);
   U1957 : INV_X1 port map( A => rd2_addr(0), ZN => n1429);
   U1958 : INV_X1 port map( A => rd2_addr(4), ZN => n1435);
   U1959 : NAND4_X1 port map( A1 => n1444, A2 => n1445, A3 => n1446, A4 => 
                           n1447, ZN => n2982);
   U1960 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_31_port, C1 => 
                           n1449, C2 => registers_9_31_port, A => n1450, ZN => 
                           n1447);
   U1961 : OAI222_X1 port map( A1 => n415, A2 => n1451, B1 => n1, B2 => n1452, 
                           C1 => n225, C2 => n1453, ZN => n1450);
   U1962 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_31_port, C1 => 
                           n1455, C2 => registers_20_31_port, A => n1456, ZN =>
                           n1446);
   U1963 : OAI22_X1 port map( A1 => n65, A2 => n1457, B1 => n290, B2 => n1458, 
                           ZN => n1456);
   U1964 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_31_port, C1 => 
                           n1460, C2 => registers_30_31_port, A => n1461, ZN =>
                           n1445);
   U1965 : OAI222_X1 port map( A1 => n416, A2 => n1462, B1 => n2, B2 => n1463, 
                           C1 => n226, C2 => n1464, ZN => n1461);
   U1966 : AOI221_X1 port map( B1 => n1465, B2 => d_in(31), C1 => n1466, C2 => 
                           d_out1_31_port, A => n1467, ZN => n1444);
   U1967 : OAI22_X1 port map( A1 => n1468, A2 => n1469, B1 => n289, B2 => n1470
                           , ZN => n1467);
   U1968 : NOR4_X1 port map( A1 => n1471, A2 => n1472, A3 => n1473, A4 => n1474
                           , ZN => n1468);
   U1969 : OAI221_X1 port map( B1 => n159, B2 => n1475, C1 => n541, C2 => n1476
                           , A => n1477, ZN => n1474);
   U1970 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_31_port, B1 => 
                           n1479, B2 => registers_19_31_port, ZN => n1477);
   U1971 : OAI221_X1 port map( B1 => n160, B2 => n1480, C1 => n542, C2 => n1481
                           , A => n1482, ZN => n1473);
   U1972 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_31_port, B1 => 
                           n1484, B2 => registers_25_31_port, ZN => n1482);
   U1973 : OAI221_X1 port map( B1 => n161, B2 => n1485, C1 => n543, C2 => n1486
                           , A => n1487, ZN => n1472);
   U1974 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_31_port, B1 => 
                           n1489, B2 => registers_6_31_port, ZN => n1487);
   U1975 : OAI221_X1 port map( B1 => n162, B2 => n1490, C1 => n544, C2 => n1491
                           , A => n1492, ZN => n1471);
   U1976 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_31_port, B1 => 
                           n1494, B2 => registers_14_31_port, ZN => n1492);
   U1977 : NAND4_X1 port map( A1 => n1495, A2 => n1496, A3 => n1497, A4 => 
                           n1498, ZN => n2981);
   U1978 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_30_port, C1 => 
                           n1449, C2 => registers_9_30_port, A => n1499, ZN => 
                           n1498);
   U1979 : OAI222_X1 port map( A1 => n417, A2 => n1451, B1 => n3, B2 => n1452, 
                           C1 => n227, C2 => n1453, ZN => n1499);
   U1980 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_30_port, C1 => 
                           n1455, C2 => registers_20_30_port, A => n1500, ZN =>
                           n1497);
   U1981 : OAI22_X1 port map( A1 => n66, A2 => n1457, B1 => n291, B2 => n1458, 
                           ZN => n1500);
   U1982 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_30_port, C1 => 
                           n1460, C2 => registers_30_30_port, A => n1501, ZN =>
                           n1496);
   U1983 : OAI222_X1 port map( A1 => n418, A2 => n1462, B1 => n4, B2 => n1463, 
                           C1 => n228, C2 => n1464, ZN => n1501);
   U1984 : AOI221_X1 port map( B1 => n1465, B2 => d_in(30), C1 => n1466, C2 => 
                           d_out1_30_port, A => n1502, ZN => n1495);
   U1985 : OAI22_X1 port map( A1 => n1503, A2 => n1469, B1 => n322, B2 => n1470
                           , ZN => n1502);
   U1986 : NOR4_X1 port map( A1 => n1504, A2 => n1505, A3 => n1506, A4 => n1507
                           , ZN => n1503);
   U1987 : OAI221_X1 port map( B1 => n97, B2 => n1475, C1 => n353, C2 => n1476,
                           A => n1508, ZN => n1507);
   U1988 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_30_port, B1 => 
                           n1479, B2 => registers_19_30_port, ZN => n1508);
   U1989 : OAI221_X1 port map( B1 => n163, B2 => n1480, C1 => n479, C2 => n1481
                           , A => n1509, ZN => n1506);
   U1990 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_30_port, B1 => 
                           n1484, B2 => registers_25_30_port, ZN => n1509);
   U1991 : OAI221_X1 port map( B1 => n164, B2 => n1485, C1 => n480, C2 => n1486
                           , A => n1510, ZN => n1505);
   U1992 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_30_port, B1 => 
                           n1489, B2 => registers_6_30_port, ZN => n1510);
   U1993 : OAI221_X1 port map( B1 => n98, B2 => n1490, C1 => n354, C2 => n1491,
                           A => n1511, ZN => n1504);
   U1994 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_30_port, B1 => 
                           n1494, B2 => registers_14_30_port, ZN => n1511);
   U1995 : NAND4_X1 port map( A1 => n1512, A2 => n1513, A3 => n1514, A4 => 
                           n1515, ZN => n2980);
   U1996 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_29_port, C1 => 
                           n1449, C2 => registers_9_29_port, A => n1516, ZN => 
                           n1515);
   U1997 : OAI222_X1 port map( A1 => n419, A2 => n1451, B1 => n5, B2 => n1452, 
                           C1 => n229, C2 => n1453, ZN => n1516);
   U1998 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_29_port, C1 => 
                           n1455, C2 => registers_20_29_port, A => n1517, ZN =>
                           n1514);
   U1999 : OAI22_X1 port map( A1 => n67, A2 => n1457, B1 => n292, B2 => n1458, 
                           ZN => n1517);
   U2000 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_29_port, C1 => 
                           n1460, C2 => registers_30_29_port, A => n1518, ZN =>
                           n1513);
   U2001 : OAI222_X1 port map( A1 => n420, A2 => n1462, B1 => n6, B2 => n1463, 
                           C1 => n230, C2 => n1464, ZN => n1518);
   U2002 : AOI221_X1 port map( B1 => n1465, B2 => d_in(29), C1 => n1466, C2 => 
                           d_out1_29_port, A => n1519, ZN => n1512);
   U2003 : OAI22_X1 port map( A1 => n1520, A2 => n1469, B1 => n323, B2 => n1470
                           , ZN => n1519);
   U2004 : NOR4_X1 port map( A1 => n1521, A2 => n1522, A3 => n1523, A4 => n1524
                           , ZN => n1520);
   U2005 : OAI221_X1 port map( B1 => n99, B2 => n1475, C1 => n355, C2 => n1476,
                           A => n1525, ZN => n1524);
   U2006 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_29_port, B1 => 
                           n1479, B2 => registers_19_29_port, ZN => n1525);
   U2007 : OAI221_X1 port map( B1 => n165, B2 => n1480, C1 => n481, C2 => n1481
                           , A => n1526, ZN => n1523);
   U2008 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_29_port, B1 => 
                           n1484, B2 => registers_25_29_port, ZN => n1526);
   U2009 : OAI221_X1 port map( B1 => n166, B2 => n1485, C1 => n482, C2 => n1486
                           , A => n1527, ZN => n1522);
   U2010 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_29_port, B1 => 
                           n1489, B2 => registers_6_29_port, ZN => n1527);
   U2011 : OAI221_X1 port map( B1 => n100, B2 => n1490, C1 => n356, C2 => n1491
                           , A => n1528, ZN => n1521);
   U2012 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_29_port, B1 => 
                           n1494, B2 => registers_14_29_port, ZN => n1528);
   U2013 : NAND4_X1 port map( A1 => n1529, A2 => n1530, A3 => n1531, A4 => 
                           n1532, ZN => n2979);
   U2014 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_28_port, C1 => 
                           n1449, C2 => registers_9_28_port, A => n1533, ZN => 
                           n1532);
   U2015 : OAI222_X1 port map( A1 => n421, A2 => n1451, B1 => n7, B2 => n1452, 
                           C1 => n231, C2 => n1453, ZN => n1533);
   U2016 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_28_port, C1 => 
                           n1455, C2 => registers_20_28_port, A => n1534, ZN =>
                           n1531);
   U2017 : OAI22_X1 port map( A1 => n68, A2 => n1457, B1 => n293, B2 => n1458, 
                           ZN => n1534);
   U2018 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_28_port, C1 => 
                           n1460, C2 => registers_30_28_port, A => n1535, ZN =>
                           n1530);
   U2019 : OAI222_X1 port map( A1 => n422, A2 => n1462, B1 => n8, B2 => n1463, 
                           C1 => n232, C2 => n1464, ZN => n1535);
   U2020 : AOI221_X1 port map( B1 => n1465, B2 => d_in(28), C1 => n1466, C2 => 
                           d_out1_28_port, A => n1536, ZN => n1529);
   U2021 : OAI22_X1 port map( A1 => n1537, A2 => n1469, B1 => n324, B2 => n1470
                           , ZN => n1536);
   U2022 : NOR4_X1 port map( A1 => n1538, A2 => n1539, A3 => n1540, A4 => n1541
                           , ZN => n1537);
   U2023 : OAI221_X1 port map( B1 => n101, B2 => n1475, C1 => n357, C2 => n1476
                           , A => n1542, ZN => n1541);
   U2024 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_28_port, B1 => 
                           n1479, B2 => registers_19_28_port, ZN => n1542);
   U2025 : OAI221_X1 port map( B1 => n167, B2 => n1480, C1 => n483, C2 => n1481
                           , A => n1543, ZN => n1540);
   U2026 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_28_port, B1 => 
                           n1484, B2 => registers_25_28_port, ZN => n1543);
   U2027 : OAI221_X1 port map( B1 => n168, B2 => n1485, C1 => n484, C2 => n1486
                           , A => n1544, ZN => n1539);
   U2028 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_28_port, B1 => 
                           n1489, B2 => registers_6_28_port, ZN => n1544);
   U2029 : OAI221_X1 port map( B1 => n102, B2 => n1490, C1 => n358, C2 => n1491
                           , A => n1545, ZN => n1538);
   U2030 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_28_port, B1 => 
                           n1494, B2 => registers_14_28_port, ZN => n1545);
   U2031 : NAND4_X1 port map( A1 => n1546, A2 => n1547, A3 => n1548, A4 => 
                           n1549, ZN => n2978);
   U2032 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_27_port, C1 => 
                           n1449, C2 => registers_9_27_port, A => n1550, ZN => 
                           n1549);
   U2033 : OAI222_X1 port map( A1 => n423, A2 => n1451, B1 => n9, B2 => n1452, 
                           C1 => n233, C2 => n1453, ZN => n1550);
   U2034 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_27_port, C1 => 
                           n1455, C2 => registers_20_27_port, A => n1551, ZN =>
                           n1548);
   U2035 : OAI22_X1 port map( A1 => n69, A2 => n1457, B1 => n294, B2 => n1458, 
                           ZN => n1551);
   U2036 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_27_port, C1 => 
                           n1460, C2 => registers_30_27_port, A => n1552, ZN =>
                           n1547);
   U2037 : OAI222_X1 port map( A1 => n424, A2 => n1462, B1 => n10, B2 => n1463,
                           C1 => n234, C2 => n1464, ZN => n1552);
   U2038 : AOI221_X1 port map( B1 => n1465, B2 => d_in(27), C1 => n1466, C2 => 
                           d_out1_27_port, A => n1553, ZN => n1546);
   U2039 : OAI22_X1 port map( A1 => n1554, A2 => n1469, B1 => n325, B2 => n1470
                           , ZN => n1553);
   U2040 : NOR4_X1 port map( A1 => n1555, A2 => n1556, A3 => n1557, A4 => n1558
                           , ZN => n1554);
   U2041 : OAI221_X1 port map( B1 => n103, B2 => n1475, C1 => n359, C2 => n1476
                           , A => n1559, ZN => n1558);
   U2042 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_27_port, B1 => 
                           n1479, B2 => registers_19_27_port, ZN => n1559);
   U2043 : OAI221_X1 port map( B1 => n169, B2 => n1480, C1 => n485, C2 => n1481
                           , A => n1560, ZN => n1557);
   U2044 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_27_port, B1 => 
                           n1484, B2 => registers_25_27_port, ZN => n1560);
   U2045 : OAI221_X1 port map( B1 => n170, B2 => n1485, C1 => n486, C2 => n1486
                           , A => n1561, ZN => n1556);
   U2046 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_27_port, B1 => 
                           n1489, B2 => registers_6_27_port, ZN => n1561);
   U2047 : OAI221_X1 port map( B1 => n104, B2 => n1490, C1 => n360, C2 => n1491
                           , A => n1562, ZN => n1555);
   U2048 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_27_port, B1 => 
                           n1494, B2 => registers_14_27_port, ZN => n1562);
   U2049 : NAND4_X1 port map( A1 => n1563, A2 => n1564, A3 => n1565, A4 => 
                           n1566, ZN => n2977);
   U2050 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_26_port, C1 => 
                           n1449, C2 => registers_9_26_port, A => n1567, ZN => 
                           n1566);
   U2051 : OAI222_X1 port map( A1 => n425, A2 => n1451, B1 => n11, B2 => n1452,
                           C1 => n235, C2 => n1453, ZN => n1567);
   U2052 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_26_port, C1 => 
                           n1455, C2 => registers_20_26_port, A => n1568, ZN =>
                           n1565);
   U2053 : OAI22_X1 port map( A1 => n70, A2 => n1457, B1 => n295, B2 => n1458, 
                           ZN => n1568);
   U2054 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_26_port, C1 => 
                           n1460, C2 => registers_30_26_port, A => n1569, ZN =>
                           n1564);
   U2055 : OAI222_X1 port map( A1 => n426, A2 => n1462, B1 => n12, B2 => n1463,
                           C1 => n236, C2 => n1464, ZN => n1569);
   U2056 : AOI221_X1 port map( B1 => n1465, B2 => d_in(26), C1 => n1466, C2 => 
                           d_out1_26_port, A => n1570, ZN => n1563);
   U2057 : OAI22_X1 port map( A1 => n1571, A2 => n1469, B1 => n326, B2 => n1470
                           , ZN => n1570);
   U2058 : NOR4_X1 port map( A1 => n1572, A2 => n1573, A3 => n1574, A4 => n1575
                           , ZN => n1571);
   U2059 : OAI221_X1 port map( B1 => n105, B2 => n1475, C1 => n361, C2 => n1476
                           , A => n1576, ZN => n1575);
   U2060 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_26_port, B1 => 
                           n1479, B2 => registers_19_26_port, ZN => n1576);
   U2061 : OAI221_X1 port map( B1 => n171, B2 => n1480, C1 => n487, C2 => n1481
                           , A => n1577, ZN => n1574);
   U2062 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_26_port, B1 => 
                           n1484, B2 => registers_25_26_port, ZN => n1577);
   U2063 : OAI221_X1 port map( B1 => n172, B2 => n1485, C1 => n488, C2 => n1486
                           , A => n1578, ZN => n1573);
   U2064 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_26_port, B1 => 
                           n1489, B2 => registers_6_26_port, ZN => n1578);
   U2065 : OAI221_X1 port map( B1 => n106, B2 => n1490, C1 => n362, C2 => n1491
                           , A => n1579, ZN => n1572);
   U2066 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_26_port, B1 => 
                           n1494, B2 => registers_14_26_port, ZN => n1579);
   U2067 : NAND4_X1 port map( A1 => n1580, A2 => n1581, A3 => n1582, A4 => 
                           n1583, ZN => n2976);
   U2068 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_25_port, C1 => 
                           n1449, C2 => registers_9_25_port, A => n1584, ZN => 
                           n1583);
   U2069 : OAI222_X1 port map( A1 => n427, A2 => n1451, B1 => n13, B2 => n1452,
                           C1 => n237, C2 => n1453, ZN => n1584);
   U2070 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_25_port, C1 => 
                           n1455, C2 => registers_20_25_port, A => n1585, ZN =>
                           n1582);
   U2071 : OAI22_X1 port map( A1 => n71, A2 => n1457, B1 => n296, B2 => n1458, 
                           ZN => n1585);
   U2072 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_25_port, C1 => 
                           n1460, C2 => registers_30_25_port, A => n1586, ZN =>
                           n1581);
   U2073 : OAI222_X1 port map( A1 => n428, A2 => n1462, B1 => n14, B2 => n1463,
                           C1 => n238, C2 => n1464, ZN => n1586);
   U2074 : AOI221_X1 port map( B1 => n1465, B2 => d_in(25), C1 => n1466, C2 => 
                           d_out1_25_port, A => n1587, ZN => n1580);
   U2075 : OAI22_X1 port map( A1 => n1588, A2 => n1469, B1 => n327, B2 => n1470
                           , ZN => n1587);
   U2076 : NOR4_X1 port map( A1 => n1589, A2 => n1590, A3 => n1591, A4 => n1592
                           , ZN => n1588);
   U2077 : OAI221_X1 port map( B1 => n107, B2 => n1475, C1 => n363, C2 => n1476
                           , A => n1593, ZN => n1592);
   U2078 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_25_port, B1 => 
                           n1479, B2 => registers_19_25_port, ZN => n1593);
   U2079 : OAI221_X1 port map( B1 => n173, B2 => n1480, C1 => n489, C2 => n1481
                           , A => n1594, ZN => n1591);
   U2080 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_25_port, B1 => 
                           n1484, B2 => registers_25_25_port, ZN => n1594);
   U2081 : OAI221_X1 port map( B1 => n174, B2 => n1485, C1 => n490, C2 => n1486
                           , A => n1595, ZN => n1590);
   U2082 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_25_port, B1 => 
                           n1489, B2 => registers_6_25_port, ZN => n1595);
   U2083 : OAI221_X1 port map( B1 => n108, B2 => n1490, C1 => n364, C2 => n1491
                           , A => n1596, ZN => n1589);
   U2084 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_25_port, B1 => 
                           n1494, B2 => registers_14_25_port, ZN => n1596);
   U2085 : NAND4_X1 port map( A1 => n1597, A2 => n1598, A3 => n1599, A4 => 
                           n1600, ZN => n2975);
   U2086 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_24_port, C1 => 
                           n1449, C2 => registers_9_24_port, A => n1601, ZN => 
                           n1600);
   U2087 : OAI222_X1 port map( A1 => n429, A2 => n1451, B1 => n15, B2 => n1452,
                           C1 => n239, C2 => n1453, ZN => n1601);
   U2088 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_24_port, C1 => 
                           n1455, C2 => registers_20_24_port, A => n1602, ZN =>
                           n1599);
   U2089 : OAI22_X1 port map( A1 => n72, A2 => n1457, B1 => n297, B2 => n1458, 
                           ZN => n1602);
   U2090 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_24_port, C1 => 
                           n1460, C2 => registers_30_24_port, A => n1603, ZN =>
                           n1598);
   U2091 : OAI222_X1 port map( A1 => n430, A2 => n1462, B1 => n16, B2 => n1463,
                           C1 => n240, C2 => n1464, ZN => n1603);
   U2092 : AOI221_X1 port map( B1 => n1465, B2 => d_in(24), C1 => n1466, C2 => 
                           d_out1_24_port, A => n1604, ZN => n1597);
   U2093 : OAI22_X1 port map( A1 => n1605, A2 => n1469, B1 => n328, B2 => n1470
                           , ZN => n1604);
   U2094 : NOR4_X1 port map( A1 => n1606, A2 => n1607, A3 => n1608, A4 => n1609
                           , ZN => n1605);
   U2095 : OAI221_X1 port map( B1 => n109, B2 => n1475, C1 => n365, C2 => n1476
                           , A => n1610, ZN => n1609);
   U2096 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_24_port, B1 => 
                           n1479, B2 => registers_19_24_port, ZN => n1610);
   U2097 : OAI221_X1 port map( B1 => n175, B2 => n1480, C1 => n491, C2 => n1481
                           , A => n1611, ZN => n1608);
   U2098 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_24_port, B1 => 
                           n1484, B2 => registers_25_24_port, ZN => n1611);
   U2099 : OAI221_X1 port map( B1 => n176, B2 => n1485, C1 => n492, C2 => n1486
                           , A => n1612, ZN => n1607);
   U2100 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_24_port, B1 => 
                           n1489, B2 => registers_6_24_port, ZN => n1612);
   U2101 : OAI221_X1 port map( B1 => n110, B2 => n1490, C1 => n366, C2 => n1491
                           , A => n1613, ZN => n1606);
   U2102 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_24_port, B1 => 
                           n1494, B2 => registers_14_24_port, ZN => n1613);
   U2103 : NAND4_X1 port map( A1 => n1614, A2 => n1615, A3 => n1616, A4 => 
                           n1617, ZN => n2974);
   U2104 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_23_port, C1 => 
                           n1449, C2 => registers_9_23_port, A => n1618, ZN => 
                           n1617);
   U2105 : OAI222_X1 port map( A1 => n431, A2 => n1451, B1 => n17, B2 => n1452,
                           C1 => n241, C2 => n1453, ZN => n1618);
   U2106 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_23_port, C1 => 
                           n1455, C2 => registers_20_23_port, A => n1619, ZN =>
                           n1616);
   U2107 : OAI22_X1 port map( A1 => n73, A2 => n1457, B1 => n298, B2 => n1458, 
                           ZN => n1619);
   U2108 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_23_port, C1 => 
                           n1460, C2 => registers_30_23_port, A => n1620, ZN =>
                           n1615);
   U2109 : OAI222_X1 port map( A1 => n432, A2 => n1462, B1 => n18_port, B2 => 
                           n1463, C1 => n242, C2 => n1464, ZN => n1620);
   U2110 : AOI221_X1 port map( B1 => n1465, B2 => d_in(23), C1 => n1466, C2 => 
                           d_out1_23_port, A => n1621, ZN => n1614);
   U2111 : OAI22_X1 port map( A1 => n1622, A2 => n1469, B1 => n329, B2 => n1470
                           , ZN => n1621);
   U2112 : NOR4_X1 port map( A1 => n1623, A2 => n1624, A3 => n1625, A4 => n1626
                           , ZN => n1622);
   U2113 : OAI221_X1 port map( B1 => n111, B2 => n1475, C1 => n367, C2 => n1476
                           , A => n1627, ZN => n1626);
   U2114 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_23_port, B1 => 
                           n1479, B2 => registers_19_23_port, ZN => n1627);
   U2115 : OAI221_X1 port map( B1 => n177, B2 => n1480, C1 => n493, C2 => n1481
                           , A => n1628, ZN => n1625);
   U2116 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_23_port, B1 => 
                           n1484, B2 => registers_25_23_port, ZN => n1628);
   U2117 : OAI221_X1 port map( B1 => n178, B2 => n1485, C1 => n494, C2 => n1486
                           , A => n1629, ZN => n1624);
   U2118 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_23_port, B1 => 
                           n1489, B2 => registers_6_23_port, ZN => n1629);
   U2119 : OAI221_X1 port map( B1 => n112, B2 => n1490, C1 => n368, C2 => n1491
                           , A => n1630, ZN => n1623);
   U2120 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_23_port, B1 => 
                           n1494, B2 => registers_14_23_port, ZN => n1630);
   U2121 : NAND4_X1 port map( A1 => n1631, A2 => n1632, A3 => n1633, A4 => 
                           n1634, ZN => n2973);
   U2122 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_22_port, C1 => 
                           n1449, C2 => registers_9_22_port, A => n1635, ZN => 
                           n1634);
   U2123 : OAI222_X1 port map( A1 => n433, A2 => n1451, B1 => n19, B2 => n1452,
                           C1 => n243, C2 => n1453, ZN => n1635);
   U2124 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_22_port, C1 => 
                           n1455, C2 => registers_20_22_port, A => n1636, ZN =>
                           n1633);
   U2125 : OAI22_X1 port map( A1 => n74, A2 => n1457, B1 => n299, B2 => n1458, 
                           ZN => n1636);
   U2126 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_22_port, C1 => 
                           n1460, C2 => registers_30_22_port, A => n1637, ZN =>
                           n1632);
   U2127 : OAI222_X1 port map( A1 => n434, A2 => n1462, B1 => n20, B2 => n1463,
                           C1 => n244, C2 => n1464, ZN => n1637);
   U2128 : AOI221_X1 port map( B1 => n1465, B2 => d_in(22), C1 => n1466, C2 => 
                           d_out1_22_port, A => n1638, ZN => n1631);
   U2129 : OAI22_X1 port map( A1 => n1639, A2 => n1469, B1 => n330, B2 => n1470
                           , ZN => n1638);
   U2130 : NOR4_X1 port map( A1 => n1640, A2 => n1641, A3 => n1642, A4 => n1643
                           , ZN => n1639);
   U2131 : OAI221_X1 port map( B1 => n113, B2 => n1475, C1 => n369, C2 => n1476
                           , A => n1644, ZN => n1643);
   U2132 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_22_port, B1 => 
                           n1479, B2 => registers_19_22_port, ZN => n1644);
   U2133 : OAI221_X1 port map( B1 => n179, B2 => n1480, C1 => n495, C2 => n1481
                           , A => n1645, ZN => n1642);
   U2134 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_22_port, B1 => 
                           n1484, B2 => registers_25_22_port, ZN => n1645);
   U2135 : OAI221_X1 port map( B1 => n180, B2 => n1485, C1 => n496, C2 => n1486
                           , A => n1646, ZN => n1641);
   U2136 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_22_port, B1 => 
                           n1489, B2 => registers_6_22_port, ZN => n1646);
   U2137 : OAI221_X1 port map( B1 => n114, B2 => n1490, C1 => n370, C2 => n1491
                           , A => n1647, ZN => n1640);
   U2138 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_22_port, B1 => 
                           n1494, B2 => registers_14_22_port, ZN => n1647);
   U2139 : NAND4_X1 port map( A1 => n1648, A2 => n1649, A3 => n1650, A4 => 
                           n1651, ZN => n2972);
   U2140 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_21_port, C1 => 
                           n1449, C2 => registers_9_21_port, A => n1652, ZN => 
                           n1651);
   U2141 : OAI222_X1 port map( A1 => n435, A2 => n1451, B1 => n21, B2 => n1452,
                           C1 => n245, C2 => n1453, ZN => n1652);
   U2142 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_21_port, C1 => 
                           n1455, C2 => registers_20_21_port, A => n1653, ZN =>
                           n1650);
   U2143 : OAI22_X1 port map( A1 => n75, A2 => n1457, B1 => n300, B2 => n1458, 
                           ZN => n1653);
   U2144 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_21_port, C1 => 
                           n1460, C2 => registers_30_21_port, A => n1654, ZN =>
                           n1649);
   U2145 : OAI222_X1 port map( A1 => n436, A2 => n1462, B1 => n22, B2 => n1463,
                           C1 => n246, C2 => n1464, ZN => n1654);
   U2146 : AOI221_X1 port map( B1 => n1465, B2 => d_in(21), C1 => n1466, C2 => 
                           d_out1_21_port, A => n1655, ZN => n1648);
   U2147 : OAI22_X1 port map( A1 => n1656, A2 => n1469, B1 => n331, B2 => n1470
                           , ZN => n1655);
   U2148 : NOR4_X1 port map( A1 => n1657, A2 => n1658, A3 => n1659, A4 => n1660
                           , ZN => n1656);
   U2149 : OAI221_X1 port map( B1 => n115, B2 => n1475, C1 => n371, C2 => n1476
                           , A => n1661, ZN => n1660);
   U2150 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_21_port, B1 => 
                           n1479, B2 => registers_19_21_port, ZN => n1661);
   U2151 : OAI221_X1 port map( B1 => n181, B2 => n1480, C1 => n497, C2 => n1481
                           , A => n1662, ZN => n1659);
   U2152 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_21_port, B1 => 
                           n1484, B2 => registers_25_21_port, ZN => n1662);
   U2153 : OAI221_X1 port map( B1 => n182, B2 => n1485, C1 => n498, C2 => n1486
                           , A => n1663, ZN => n1658);
   U2154 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_21_port, B1 => 
                           n1489, B2 => registers_6_21_port, ZN => n1663);
   U2155 : OAI221_X1 port map( B1 => n116, B2 => n1490, C1 => n372, C2 => n1491
                           , A => n1664, ZN => n1657);
   U2156 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_21_port, B1 => 
                           n1494, B2 => registers_14_21_port, ZN => n1664);
   U2157 : NAND4_X1 port map( A1 => n1665, A2 => n1666, A3 => n1667, A4 => 
                           n1668, ZN => n2971);
   U2158 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_20_port, C1 => 
                           n1449, C2 => registers_9_20_port, A => n1669, ZN => 
                           n1668);
   U2159 : OAI222_X1 port map( A1 => n437, A2 => n1451, B1 => n23, B2 => n1452,
                           C1 => n247, C2 => n1453, ZN => n1669);
   U2160 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_20_port, C1 => 
                           n1455, C2 => registers_20_20_port, A => n1670, ZN =>
                           n1667);
   U2161 : OAI22_X1 port map( A1 => n76, A2 => n1457, B1 => n301, B2 => n1458, 
                           ZN => n1670);
   U2162 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_20_port, C1 => 
                           n1460, C2 => registers_30_20_port, A => n1671, ZN =>
                           n1666);
   U2163 : OAI222_X1 port map( A1 => n438, A2 => n1462, B1 => n24, B2 => n1463,
                           C1 => n248, C2 => n1464, ZN => n1671);
   U2164 : AOI221_X1 port map( B1 => n1465, B2 => d_in(20), C1 => n1466, C2 => 
                           d_out1_20_port, A => n1672, ZN => n1665);
   U2165 : OAI22_X1 port map( A1 => n1673, A2 => n1469, B1 => n332, B2 => n1470
                           , ZN => n1672);
   U2166 : NOR4_X1 port map( A1 => n1674, A2 => n1675, A3 => n1676, A4 => n1677
                           , ZN => n1673);
   U2167 : OAI221_X1 port map( B1 => n117, B2 => n1475, C1 => n373, C2 => n1476
                           , A => n1678, ZN => n1677);
   U2168 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_20_port, B1 => 
                           n1479, B2 => registers_19_20_port, ZN => n1678);
   U2169 : OAI221_X1 port map( B1 => n183, B2 => n1480, C1 => n499, C2 => n1481
                           , A => n1679, ZN => n1676);
   U2170 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_20_port, B1 => 
                           n1484, B2 => registers_25_20_port, ZN => n1679);
   U2171 : OAI221_X1 port map( B1 => n184, B2 => n1485, C1 => n500, C2 => n1486
                           , A => n1680, ZN => n1675);
   U2172 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_20_port, B1 => 
                           n1489, B2 => registers_6_20_port, ZN => n1680);
   U2173 : OAI221_X1 port map( B1 => n118, B2 => n1490, C1 => n374, C2 => n1491
                           , A => n1681, ZN => n1674);
   U2174 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_20_port, B1 => 
                           n1494, B2 => registers_14_20_port, ZN => n1681);
   U2175 : NAND4_X1 port map( A1 => n1682, A2 => n1683, A3 => n1684, A4 => 
                           n1685, ZN => n2970);
   U2176 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_19_port, C1 => 
                           n1449, C2 => registers_9_19_port, A => n1686, ZN => 
                           n1685);
   U2177 : OAI222_X1 port map( A1 => n439, A2 => n1451, B1 => n25, B2 => n1452,
                           C1 => n249, C2 => n1453, ZN => n1686);
   U2178 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_19_port, C1 => 
                           n1455, C2 => registers_20_19_port, A => n1687, ZN =>
                           n1684);
   U2179 : OAI22_X1 port map( A1 => n77, A2 => n1457, B1 => n302, B2 => n1458, 
                           ZN => n1687);
   U2180 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_19_port, C1 => 
                           n1460, C2 => registers_30_19_port, A => n1688, ZN =>
                           n1683);
   U2181 : OAI222_X1 port map( A1 => n440, A2 => n1462, B1 => n26, B2 => n1463,
                           C1 => n250, C2 => n1464, ZN => n1688);
   U2182 : AOI221_X1 port map( B1 => n1465, B2 => d_in(19), C1 => n1466, C2 => 
                           d_out1_19_port, A => n1689, ZN => n1682);
   U2183 : OAI22_X1 port map( A1 => n1690, A2 => n1469, B1 => n333, B2 => n1470
                           , ZN => n1689);
   U2184 : NOR4_X1 port map( A1 => n1691, A2 => n1692, A3 => n1693, A4 => n1694
                           , ZN => n1690);
   U2185 : OAI221_X1 port map( B1 => n119, B2 => n1475, C1 => n375, C2 => n1476
                           , A => n1695, ZN => n1694);
   U2186 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_19_port, B1 => 
                           n1479, B2 => registers_19_19_port, ZN => n1695);
   U2187 : OAI221_X1 port map( B1 => n185, B2 => n1480, C1 => n501, C2 => n1481
                           , A => n1696, ZN => n1693);
   U2188 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_19_port, B1 => 
                           n1484, B2 => registers_25_19_port, ZN => n1696);
   U2189 : OAI221_X1 port map( B1 => n186, B2 => n1485, C1 => n502, C2 => n1486
                           , A => n1697, ZN => n1692);
   U2190 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_19_port, B1 => 
                           n1489, B2 => registers_6_19_port, ZN => n1697);
   U2191 : OAI221_X1 port map( B1 => n120, B2 => n1490, C1 => n376, C2 => n1491
                           , A => n1698, ZN => n1691);
   U2192 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_19_port, B1 => 
                           n1494, B2 => registers_14_19_port, ZN => n1698);
   U2193 : NAND4_X1 port map( A1 => n1699, A2 => n1700, A3 => n1701, A4 => 
                           n1702, ZN => n2969);
   U2194 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_18_port, C1 => 
                           n1449, C2 => registers_9_18_port, A => n1703, ZN => 
                           n1702);
   U2195 : OAI222_X1 port map( A1 => n441, A2 => n1451, B1 => n27, B2 => n1452,
                           C1 => n251, C2 => n1453, ZN => n1703);
   U2196 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_18_port, C1 => 
                           n1455, C2 => registers_20_18_port, A => n1704, ZN =>
                           n1701);
   U2197 : OAI22_X1 port map( A1 => n78, A2 => n1457, B1 => n303, B2 => n1458, 
                           ZN => n1704);
   U2198 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_18_port, C1 => 
                           n1460, C2 => registers_30_18_port, A => n1705, ZN =>
                           n1700);
   U2199 : OAI222_X1 port map( A1 => n442, A2 => n1462, B1 => n28, B2 => n1463,
                           C1 => n252, C2 => n1464, ZN => n1705);
   U2200 : AOI221_X1 port map( B1 => n1465, B2 => d_in(18), C1 => n1466, C2 => 
                           d_out1_18_port, A => n1706, ZN => n1699);
   U2201 : OAI22_X1 port map( A1 => n1707, A2 => n1469, B1 => n334, B2 => n1470
                           , ZN => n1706);
   U2202 : NOR4_X1 port map( A1 => n1708, A2 => n1709, A3 => n1710, A4 => n1711
                           , ZN => n1707);
   U2203 : OAI221_X1 port map( B1 => n121, B2 => n1475, C1 => n377, C2 => n1476
                           , A => n1712, ZN => n1711);
   U2204 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_18_port, B1 => 
                           n1479, B2 => registers_19_18_port, ZN => n1712);
   U2205 : OAI221_X1 port map( B1 => n187, B2 => n1480, C1 => n503, C2 => n1481
                           , A => n1713, ZN => n1710);
   U2206 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_18_port, B1 => 
                           n1484, B2 => registers_25_18_port, ZN => n1713);
   U2207 : OAI221_X1 port map( B1 => n188, B2 => n1485, C1 => n504, C2 => n1486
                           , A => n1714, ZN => n1709);
   U2208 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_18_port, B1 => 
                           n1489, B2 => registers_6_18_port, ZN => n1714);
   U2209 : OAI221_X1 port map( B1 => n122, B2 => n1490, C1 => n378, C2 => n1491
                           , A => n1715, ZN => n1708);
   U2210 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_18_port, B1 => 
                           n1494, B2 => registers_14_18_port, ZN => n1715);
   U2211 : NAND4_X1 port map( A1 => n1716, A2 => n1717, A3 => n1718, A4 => 
                           n1719, ZN => n2968);
   U2212 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_17_port, C1 => 
                           n1449, C2 => registers_9_17_port, A => n1720, ZN => 
                           n1719);
   U2213 : OAI222_X1 port map( A1 => n443, A2 => n1451, B1 => n29, B2 => n1452,
                           C1 => n253, C2 => n1453, ZN => n1720);
   U2214 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_17_port, C1 => 
                           n1455, C2 => registers_20_17_port, A => n1721, ZN =>
                           n1718);
   U2215 : OAI22_X1 port map( A1 => n79, A2 => n1457, B1 => n304, B2 => n1458, 
                           ZN => n1721);
   U2216 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_17_port, C1 => 
                           n1460, C2 => registers_30_17_port, A => n1722, ZN =>
                           n1717);
   U2217 : OAI222_X1 port map( A1 => n444, A2 => n1462, B1 => n30, B2 => n1463,
                           C1 => n254, C2 => n1464, ZN => n1722);
   U2218 : AOI221_X1 port map( B1 => n1465, B2 => d_in(17), C1 => n1466, C2 => 
                           d_out1_17_port, A => n1723, ZN => n1716);
   U2219 : OAI22_X1 port map( A1 => n1724, A2 => n1469, B1 => n335, B2 => n1470
                           , ZN => n1723);
   U2220 : NOR4_X1 port map( A1 => n1725, A2 => n1726, A3 => n1727, A4 => n1728
                           , ZN => n1724);
   U2221 : OAI221_X1 port map( B1 => n123, B2 => n1475, C1 => n379, C2 => n1476
                           , A => n1729, ZN => n1728);
   U2222 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_17_port, B1 => 
                           n1479, B2 => registers_19_17_port, ZN => n1729);
   U2223 : OAI221_X1 port map( B1 => n189, B2 => n1480, C1 => n505, C2 => n1481
                           , A => n1730, ZN => n1727);
   U2224 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_17_port, B1 => 
                           n1484, B2 => registers_25_17_port, ZN => n1730);
   U2225 : OAI221_X1 port map( B1 => n190, B2 => n1485, C1 => n506, C2 => n1486
                           , A => n1731, ZN => n1726);
   U2226 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_17_port, B1 => 
                           n1489, B2 => registers_6_17_port, ZN => n1731);
   U2227 : OAI221_X1 port map( B1 => n124, B2 => n1490, C1 => n380, C2 => n1491
                           , A => n1732, ZN => n1725);
   U2228 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_17_port, B1 => 
                           n1494, B2 => registers_14_17_port, ZN => n1732);
   U2229 : NAND4_X1 port map( A1 => n1733, A2 => n1734, A3 => n1735, A4 => 
                           n1736, ZN => n2967);
   U2230 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_16_port, C1 => 
                           n1449, C2 => registers_9_16_port, A => n1737, ZN => 
                           n1736);
   U2231 : OAI222_X1 port map( A1 => n445, A2 => n1451, B1 => n31, B2 => n1452,
                           C1 => n255, C2 => n1453, ZN => n1737);
   U2232 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_16_port, C1 => 
                           n1455, C2 => registers_20_16_port, A => n1738, ZN =>
                           n1735);
   U2233 : OAI22_X1 port map( A1 => n80, A2 => n1457, B1 => n305, B2 => n1458, 
                           ZN => n1738);
   U2234 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_16_port, C1 => 
                           n1460, C2 => registers_30_16_port, A => n1739, ZN =>
                           n1734);
   U2235 : OAI222_X1 port map( A1 => n446, A2 => n1462, B1 => n32, B2 => n1463,
                           C1 => n256, C2 => n1464, ZN => n1739);
   U2236 : AOI221_X1 port map( B1 => n1465, B2 => d_in(16), C1 => n1466, C2 => 
                           d_out1_16_port, A => n1740, ZN => n1733);
   U2237 : OAI22_X1 port map( A1 => n1741, A2 => n1469, B1 => n336, B2 => n1470
                           , ZN => n1740);
   U2238 : NOR4_X1 port map( A1 => n1742, A2 => n1743, A3 => n1744, A4 => n1745
                           , ZN => n1741);
   U2239 : OAI221_X1 port map( B1 => n125, B2 => n1475, C1 => n381, C2 => n1476
                           , A => n1746, ZN => n1745);
   U2240 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_16_port, B1 => 
                           n1479, B2 => registers_19_16_port, ZN => n1746);
   U2241 : OAI221_X1 port map( B1 => n191, B2 => n1480, C1 => n507, C2 => n1481
                           , A => n1747, ZN => n1744);
   U2242 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_16_port, B1 => 
                           n1484, B2 => registers_25_16_port, ZN => n1747);
   U2243 : OAI221_X1 port map( B1 => n192, B2 => n1485, C1 => n508, C2 => n1486
                           , A => n1748, ZN => n1743);
   U2244 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_16_port, B1 => 
                           n1489, B2 => registers_6_16_port, ZN => n1748);
   U2245 : OAI221_X1 port map( B1 => n126, B2 => n1490, C1 => n382, C2 => n1491
                           , A => n1749, ZN => n1742);
   U2246 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_16_port, B1 => 
                           n1494, B2 => registers_14_16_port, ZN => n1749);
   U2247 : NAND4_X1 port map( A1 => n1750, A2 => n1751, A3 => n1752, A4 => 
                           n1753, ZN => n2966);
   U2248 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_15_port, C1 => 
                           n1449, C2 => registers_9_15_port, A => n1754, ZN => 
                           n1753);
   U2249 : OAI222_X1 port map( A1 => n447, A2 => n1451, B1 => n33, B2 => n1452,
                           C1 => n257, C2 => n1453, ZN => n1754);
   U2250 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_15_port, C1 => 
                           n1455, C2 => registers_20_15_port, A => n1755, ZN =>
                           n1752);
   U2251 : OAI22_X1 port map( A1 => n81, A2 => n1457, B1 => n306, B2 => n1458, 
                           ZN => n1755);
   U2252 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_15_port, C1 => 
                           n1460, C2 => registers_30_15_port, A => n1756, ZN =>
                           n1751);
   U2253 : OAI222_X1 port map( A1 => n448, A2 => n1462, B1 => n34, B2 => n1463,
                           C1 => n258, C2 => n1464, ZN => n1756);
   U2254 : AOI221_X1 port map( B1 => n1465, B2 => d_in(15), C1 => n1466, C2 => 
                           d_out1_15_port, A => n1757, ZN => n1750);
   U2255 : OAI22_X1 port map( A1 => n1758, A2 => n1469, B1 => n337, B2 => n1470
                           , ZN => n1757);
   U2256 : NOR4_X1 port map( A1 => n1759, A2 => n1760, A3 => n1761, A4 => n1762
                           , ZN => n1758);
   U2257 : OAI221_X1 port map( B1 => n127, B2 => n1475, C1 => n383, C2 => n1476
                           , A => n1763, ZN => n1762);
   U2258 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_15_port, B1 => 
                           n1479, B2 => registers_19_15_port, ZN => n1763);
   U2259 : OAI221_X1 port map( B1 => n193, B2 => n1480, C1 => n509, C2 => n1481
                           , A => n1764, ZN => n1761);
   U2260 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_15_port, B1 => 
                           n1484, B2 => registers_25_15_port, ZN => n1764);
   U2261 : OAI221_X1 port map( B1 => n194, B2 => n1485, C1 => n510, C2 => n1486
                           , A => n1765, ZN => n1760);
   U2262 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_15_port, B1 => 
                           n1489, B2 => registers_6_15_port, ZN => n1765);
   U2263 : OAI221_X1 port map( B1 => n128, B2 => n1490, C1 => n384, C2 => n1491
                           , A => n1766, ZN => n1759);
   U2264 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_15_port, B1 => 
                           n1494, B2 => registers_14_15_port, ZN => n1766);
   U2265 : NAND4_X1 port map( A1 => n1767, A2 => n1768, A3 => n1769, A4 => 
                           n1770, ZN => n2965);
   U2266 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_14_port, C1 => 
                           n1449, C2 => registers_9_14_port, A => n1771, ZN => 
                           n1770);
   U2267 : OAI222_X1 port map( A1 => n449, A2 => n1451, B1 => n35, B2 => n1452,
                           C1 => n259, C2 => n1453, ZN => n1771);
   U2268 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_14_port, C1 => 
                           n1455, C2 => registers_20_14_port, A => n1772, ZN =>
                           n1769);
   U2269 : OAI22_X1 port map( A1 => n82, A2 => n1457, B1 => n307, B2 => n1458, 
                           ZN => n1772);
   U2270 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_14_port, C1 => 
                           n1460, C2 => registers_30_14_port, A => n1773, ZN =>
                           n1768);
   U2271 : OAI222_X1 port map( A1 => n450, A2 => n1462, B1 => n36, B2 => n1463,
                           C1 => n260, C2 => n1464, ZN => n1773);
   U2272 : AOI221_X1 port map( B1 => n1465, B2 => d_in(14), C1 => n1466, C2 => 
                           d_out1_14_port, A => n1774, ZN => n1767);
   U2273 : OAI22_X1 port map( A1 => n1775, A2 => n1469, B1 => n338, B2 => n1470
                           , ZN => n1774);
   U2274 : NOR4_X1 port map( A1 => n1776, A2 => n1777, A3 => n1778, A4 => n1779
                           , ZN => n1775);
   U2275 : OAI221_X1 port map( B1 => n129, B2 => n1475, C1 => n385, C2 => n1476
                           , A => n1780, ZN => n1779);
   U2276 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_14_port, B1 => 
                           n1479, B2 => registers_19_14_port, ZN => n1780);
   U2277 : OAI221_X1 port map( B1 => n195, B2 => n1480, C1 => n511, C2 => n1481
                           , A => n1781, ZN => n1778);
   U2278 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_14_port, B1 => 
                           n1484, B2 => registers_25_14_port, ZN => n1781);
   U2279 : OAI221_X1 port map( B1 => n196, B2 => n1485, C1 => n512, C2 => n1486
                           , A => n1782, ZN => n1777);
   U2280 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_14_port, B1 => 
                           n1489, B2 => registers_6_14_port, ZN => n1782);
   U2281 : OAI221_X1 port map( B1 => n130, B2 => n1490, C1 => n386, C2 => n1491
                           , A => n1783, ZN => n1776);
   U2282 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_14_port, B1 => 
                           n1494, B2 => registers_14_14_port, ZN => n1783);
   U2283 : NAND4_X1 port map( A1 => n1784, A2 => n1785, A3 => n1786, A4 => 
                           n1787, ZN => n2964);
   U2284 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_13_port, C1 => 
                           n1449, C2 => registers_9_13_port, A => n1788, ZN => 
                           n1787);
   U2285 : OAI222_X1 port map( A1 => n451, A2 => n1451, B1 => n37, B2 => n1452,
                           C1 => n261, C2 => n1453, ZN => n1788);
   U2286 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_13_port, C1 => 
                           n1455, C2 => registers_20_13_port, A => n1789, ZN =>
                           n1786);
   U2287 : OAI22_X1 port map( A1 => n83, A2 => n1457, B1 => n308, B2 => n1458, 
                           ZN => n1789);
   U2288 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_13_port, C1 => 
                           n1460, C2 => registers_30_13_port, A => n1790, ZN =>
                           n1785);
   U2289 : OAI222_X1 port map( A1 => n452, A2 => n1462, B1 => n38, B2 => n1463,
                           C1 => n262, C2 => n1464, ZN => n1790);
   U2290 : AOI221_X1 port map( B1 => n1465, B2 => d_in(13), C1 => n1466, C2 => 
                           d_out1_13_port, A => n1791, ZN => n1784);
   U2291 : OAI22_X1 port map( A1 => n1792, A2 => n1469, B1 => n339, B2 => n1470
                           , ZN => n1791);
   U2292 : NOR4_X1 port map( A1 => n1793, A2 => n1794, A3 => n1795, A4 => n1796
                           , ZN => n1792);
   U2293 : OAI221_X1 port map( B1 => n131, B2 => n1475, C1 => n387, C2 => n1476
                           , A => n1797, ZN => n1796);
   U2294 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_13_port, B1 => 
                           n1479, B2 => registers_19_13_port, ZN => n1797);
   U2295 : OAI221_X1 port map( B1 => n197, B2 => n1480, C1 => n513, C2 => n1481
                           , A => n1798, ZN => n1795);
   U2296 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_13_port, B1 => 
                           n1484, B2 => registers_25_13_port, ZN => n1798);
   U2297 : OAI221_X1 port map( B1 => n198, B2 => n1485, C1 => n514, C2 => n1486
                           , A => n1799, ZN => n1794);
   U2298 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_13_port, B1 => 
                           n1489, B2 => registers_6_13_port, ZN => n1799);
   U2299 : OAI221_X1 port map( B1 => n132, B2 => n1490, C1 => n388, C2 => n1491
                           , A => n1800, ZN => n1793);
   U2300 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_13_port, B1 => 
                           n1494, B2 => registers_14_13_port, ZN => n1800);
   U2301 : NAND4_X1 port map( A1 => n1801, A2 => n1802, A3 => n1803, A4 => 
                           n1804, ZN => n2963);
   U2302 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_12_port, C1 => 
                           n1449, C2 => registers_9_12_port, A => n1805, ZN => 
                           n1804);
   U2303 : OAI222_X1 port map( A1 => n453, A2 => n1451, B1 => n39, B2 => n1452,
                           C1 => n263, C2 => n1453, ZN => n1805);
   U2304 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_12_port, C1 => 
                           n1455, C2 => registers_20_12_port, A => n1806, ZN =>
                           n1803);
   U2305 : OAI22_X1 port map( A1 => n84, A2 => n1457, B1 => n309, B2 => n1458, 
                           ZN => n1806);
   U2306 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_12_port, C1 => 
                           n1460, C2 => registers_30_12_port, A => n1807, ZN =>
                           n1802);
   U2307 : OAI222_X1 port map( A1 => n454, A2 => n1462, B1 => n40, B2 => n1463,
                           C1 => n264, C2 => n1464, ZN => n1807);
   U2308 : AOI221_X1 port map( B1 => n1465, B2 => d_in(12), C1 => n1466, C2 => 
                           d_out1_12_port, A => n1808, ZN => n1801);
   U2309 : OAI22_X1 port map( A1 => n1809, A2 => n1469, B1 => n340, B2 => n1470
                           , ZN => n1808);
   U2310 : NOR4_X1 port map( A1 => n1810, A2 => n1811, A3 => n1812, A4 => n1813
                           , ZN => n1809);
   U2311 : OAI221_X1 port map( B1 => n133, B2 => n1475, C1 => n389, C2 => n1476
                           , A => n1814, ZN => n1813);
   U2312 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_12_port, B1 => 
                           n1479, B2 => registers_19_12_port, ZN => n1814);
   U2313 : OAI221_X1 port map( B1 => n199, B2 => n1480, C1 => n515, C2 => n1481
                           , A => n1815, ZN => n1812);
   U2314 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_12_port, B1 => 
                           n1484, B2 => registers_25_12_port, ZN => n1815);
   U2315 : OAI221_X1 port map( B1 => n200, B2 => n1485, C1 => n516, C2 => n1486
                           , A => n1816, ZN => n1811);
   U2316 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_12_port, B1 => 
                           n1489, B2 => registers_6_12_port, ZN => n1816);
   U2317 : OAI221_X1 port map( B1 => n134, B2 => n1490, C1 => n390, C2 => n1491
                           , A => n1817, ZN => n1810);
   U2318 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_12_port, B1 => 
                           n1494, B2 => registers_14_12_port, ZN => n1817);
   U2319 : NAND4_X1 port map( A1 => n1818, A2 => n1819, A3 => n1820, A4 => 
                           n1821, ZN => n2962);
   U2320 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_11_port, C1 => 
                           n1449, C2 => registers_9_11_port, A => n1822, ZN => 
                           n1821);
   U2321 : OAI222_X1 port map( A1 => n455, A2 => n1451, B1 => n41, B2 => n1452,
                           C1 => n265, C2 => n1453, ZN => n1822);
   U2322 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_11_port, C1 => 
                           n1455, C2 => registers_20_11_port, A => n1823, ZN =>
                           n1820);
   U2323 : OAI22_X1 port map( A1 => n85, A2 => n1457, B1 => n310, B2 => n1458, 
                           ZN => n1823);
   U2324 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_11_port, C1 => 
                           n1460, C2 => registers_30_11_port, A => n1824, ZN =>
                           n1819);
   U2325 : OAI222_X1 port map( A1 => n456, A2 => n1462, B1 => n42, B2 => n1463,
                           C1 => n266, C2 => n1464, ZN => n1824);
   U2326 : AOI221_X1 port map( B1 => n1465, B2 => d_in(11), C1 => n1466, C2 => 
                           d_out1_11_port, A => n1825, ZN => n1818);
   U2327 : OAI22_X1 port map( A1 => n1826, A2 => n1469, B1 => n341, B2 => n1470
                           , ZN => n1825);
   U2328 : NOR4_X1 port map( A1 => n1827, A2 => n1828, A3 => n1829, A4 => n1830
                           , ZN => n1826);
   U2329 : OAI221_X1 port map( B1 => n135, B2 => n1475, C1 => n391, C2 => n1476
                           , A => n1831, ZN => n1830);
   U2330 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_11_port, B1 => 
                           n1479, B2 => registers_19_11_port, ZN => n1831);
   U2331 : OAI221_X1 port map( B1 => n201, B2 => n1480, C1 => n517, C2 => n1481
                           , A => n1832, ZN => n1829);
   U2332 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_11_port, B1 => 
                           n1484, B2 => registers_25_11_port, ZN => n1832);
   U2333 : OAI221_X1 port map( B1 => n202, B2 => n1485, C1 => n518, C2 => n1486
                           , A => n1833, ZN => n1828);
   U2334 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_11_port, B1 => 
                           n1489, B2 => registers_6_11_port, ZN => n1833);
   U2335 : OAI221_X1 port map( B1 => n136, B2 => n1490, C1 => n392, C2 => n1491
                           , A => n1834, ZN => n1827);
   U2336 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_11_port, B1 => 
                           n1494, B2 => registers_14_11_port, ZN => n1834);
   U2337 : NAND4_X1 port map( A1 => n1835, A2 => n1836, A3 => n1837, A4 => 
                           n1838, ZN => n2961);
   U2338 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_10_port, C1 => 
                           n1449, C2 => registers_9_10_port, A => n1839, ZN => 
                           n1838);
   U2339 : OAI222_X1 port map( A1 => n457, A2 => n1451, B1 => n43, B2 => n1452,
                           C1 => n267, C2 => n1453, ZN => n1839);
   U2340 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_10_port, C1 => 
                           n1455, C2 => registers_20_10_port, A => n1840, ZN =>
                           n1837);
   U2341 : OAI22_X1 port map( A1 => n86, A2 => n1457, B1 => n311, B2 => n1458, 
                           ZN => n1840);
   U2342 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_10_port, C1 => 
                           n1460, C2 => registers_30_10_port, A => n1841, ZN =>
                           n1836);
   U2343 : OAI222_X1 port map( A1 => n458, A2 => n1462, B1 => n44, B2 => n1463,
                           C1 => n268, C2 => n1464, ZN => n1841);
   U2344 : AOI221_X1 port map( B1 => n1465, B2 => d_in(10), C1 => n1466, C2 => 
                           d_out1_10_port, A => n1842, ZN => n1835);
   U2345 : OAI22_X1 port map( A1 => n1843, A2 => n1469, B1 => n342, B2 => n1470
                           , ZN => n1842);
   U2346 : NOR4_X1 port map( A1 => n1844, A2 => n1845, A3 => n1846, A4 => n1847
                           , ZN => n1843);
   U2347 : OAI221_X1 port map( B1 => n137, B2 => n1475, C1 => n393, C2 => n1476
                           , A => n1848, ZN => n1847);
   U2348 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_10_port, B1 => 
                           n1479, B2 => registers_19_10_port, ZN => n1848);
   U2349 : OAI221_X1 port map( B1 => n203, B2 => n1480, C1 => n519, C2 => n1481
                           , A => n1849, ZN => n1846);
   U2350 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_10_port, B1 => 
                           n1484, B2 => registers_25_10_port, ZN => n1849);
   U2351 : OAI221_X1 port map( B1 => n204, B2 => n1485, C1 => n520, C2 => n1486
                           , A => n1850, ZN => n1845);
   U2352 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_10_port, B1 => 
                           n1489, B2 => registers_6_10_port, ZN => n1850);
   U2353 : OAI221_X1 port map( B1 => n138, B2 => n1490, C1 => n394, C2 => n1491
                           , A => n1851, ZN => n1844);
   U2354 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_10_port, B1 => 
                           n1494, B2 => registers_14_10_port, ZN => n1851);
   U2355 : NAND4_X1 port map( A1 => n1852, A2 => n1853, A3 => n1854, A4 => 
                           n1855, ZN => n2960);
   U2356 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_9_port, C1 => 
                           n1449, C2 => registers_9_9_port, A => n1856, ZN => 
                           n1855);
   U2357 : OAI222_X1 port map( A1 => n459, A2 => n1451, B1 => n45, B2 => n1452,
                           C1 => n269, C2 => n1453, ZN => n1856);
   U2358 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_9_port, C1 => 
                           n1455, C2 => registers_20_9_port, A => n1857, ZN => 
                           n1854);
   U2359 : OAI22_X1 port map( A1 => n87, A2 => n1457, B1 => n312, B2 => n1458, 
                           ZN => n1857);
   U2360 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_9_port, C1 => 
                           n1460, C2 => registers_30_9_port, A => n1858, ZN => 
                           n1853);
   U2361 : OAI222_X1 port map( A1 => n460, A2 => n1462, B1 => n46, B2 => n1463,
                           C1 => n270, C2 => n1464, ZN => n1858);
   U2362 : AOI221_X1 port map( B1 => n1465, B2 => d_in(9), C1 => n1466, C2 => 
                           d_out1_9_port, A => n1859, ZN => n1852);
   U2363 : OAI22_X1 port map( A1 => n1860, A2 => n1469, B1 => n343, B2 => n1470
                           , ZN => n1859);
   U2364 : NOR4_X1 port map( A1 => n1861, A2 => n1862, A3 => n1863, A4 => n1864
                           , ZN => n1860);
   U2365 : OAI221_X1 port map( B1 => n139, B2 => n1475, C1 => n395, C2 => n1476
                           , A => n1865, ZN => n1864);
   U2366 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_9_port, B1 => 
                           n1479, B2 => registers_19_9_port, ZN => n1865);
   U2367 : OAI221_X1 port map( B1 => n205, B2 => n1480, C1 => n521, C2 => n1481
                           , A => n1866, ZN => n1863);
   U2368 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_9_port, B1 => 
                           n1484, B2 => registers_25_9_port, ZN => n1866);
   U2369 : OAI221_X1 port map( B1 => n206, B2 => n1485, C1 => n522, C2 => n1486
                           , A => n1867, ZN => n1862);
   U2370 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_9_port, B1 => 
                           n1489, B2 => registers_6_9_port, ZN => n1867);
   U2371 : OAI221_X1 port map( B1 => n140, B2 => n1490, C1 => n396, C2 => n1491
                           , A => n1868, ZN => n1861);
   U2372 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_9_port, B1 => 
                           n1494, B2 => registers_14_9_port, ZN => n1868);
   U2373 : NAND4_X1 port map( A1 => n1869, A2 => n1870, A3 => n1871, A4 => 
                           n1872, ZN => n2959);
   U2374 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_8_port, C1 => 
                           n1449, C2 => registers_9_8_port, A => n1873, ZN => 
                           n1872);
   U2375 : OAI222_X1 port map( A1 => n461, A2 => n1451, B1 => n47, B2 => n1452,
                           C1 => n271, C2 => n1453, ZN => n1873);
   U2376 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_8_port, C1 => 
                           n1455, C2 => registers_20_8_port, A => n1874, ZN => 
                           n1871);
   U2377 : OAI22_X1 port map( A1 => n88, A2 => n1457, B1 => n313, B2 => n1458, 
                           ZN => n1874);
   U2378 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_8_port, C1 => 
                           n1460, C2 => registers_30_8_port, A => n1875, ZN => 
                           n1870);
   U2379 : OAI222_X1 port map( A1 => n462, A2 => n1462, B1 => n48, B2 => n1463,
                           C1 => n272, C2 => n1464, ZN => n1875);
   U2380 : AOI221_X1 port map( B1 => n1465, B2 => d_in(8), C1 => n1466, C2 => 
                           d_out1_8_port, A => n1876, ZN => n1869);
   U2381 : OAI22_X1 port map( A1 => n1877, A2 => n1469, B1 => n344, B2 => n1470
                           , ZN => n1876);
   U2382 : NOR4_X1 port map( A1 => n1878, A2 => n1879, A3 => n1880, A4 => n1881
                           , ZN => n1877);
   U2383 : OAI221_X1 port map( B1 => n141, B2 => n1475, C1 => n397, C2 => n1476
                           , A => n1882, ZN => n1881);
   U2384 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_8_port, B1 => 
                           n1479, B2 => registers_19_8_port, ZN => n1882);
   U2385 : OAI221_X1 port map( B1 => n207, B2 => n1480, C1 => n523, C2 => n1481
                           , A => n1883, ZN => n1880);
   U2386 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_8_port, B1 => 
                           n1484, B2 => registers_25_8_port, ZN => n1883);
   U2387 : OAI221_X1 port map( B1 => n208, B2 => n1485, C1 => n524, C2 => n1486
                           , A => n1884, ZN => n1879);
   U2388 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_8_port, B1 => 
                           n1489, B2 => registers_6_8_port, ZN => n1884);
   U2389 : OAI221_X1 port map( B1 => n142, B2 => n1490, C1 => n398, C2 => n1491
                           , A => n1885, ZN => n1878);
   U2390 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_8_port, B1 => 
                           n1494, B2 => registers_14_8_port, ZN => n1885);
   U2391 : NAND4_X1 port map( A1 => n1886, A2 => n1887, A3 => n1888, A4 => 
                           n1889, ZN => n2958);
   U2392 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_7_port, C1 => 
                           n1449, C2 => registers_9_7_port, A => n1890, ZN => 
                           n1889);
   U2393 : OAI222_X1 port map( A1 => n463, A2 => n1451, B1 => n49, B2 => n1452,
                           C1 => n273, C2 => n1453, ZN => n1890);
   U2394 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_7_port, C1 => 
                           n1455, C2 => registers_20_7_port, A => n1891, ZN => 
                           n1888);
   U2395 : OAI22_X1 port map( A1 => n89, A2 => n1457, B1 => n314, B2 => n1458, 
                           ZN => n1891);
   U2396 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_7_port, C1 => 
                           n1460, C2 => registers_30_7_port, A => n1892, ZN => 
                           n1887);
   U2397 : OAI222_X1 port map( A1 => n464, A2 => n1462, B1 => n50, B2 => n1463,
                           C1 => n274, C2 => n1464, ZN => n1892);
   U2398 : AOI221_X1 port map( B1 => n1465, B2 => d_in(7), C1 => n1466, C2 => 
                           d_out1_7_port, A => n1893, ZN => n1886);
   U2399 : OAI22_X1 port map( A1 => n1894, A2 => n1469, B1 => n345, B2 => n1470
                           , ZN => n1893);
   U2400 : NOR4_X1 port map( A1 => n1895, A2 => n1896, A3 => n1897, A4 => n1898
                           , ZN => n1894);
   U2401 : OAI221_X1 port map( B1 => n143, B2 => n1475, C1 => n399, C2 => n1476
                           , A => n1899, ZN => n1898);
   U2402 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_7_port, B1 => 
                           n1479, B2 => registers_19_7_port, ZN => n1899);
   U2403 : OAI221_X1 port map( B1 => n209, B2 => n1480, C1 => n525, C2 => n1481
                           , A => n1900, ZN => n1897);
   U2404 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_7_port, B1 => 
                           n1484, B2 => registers_25_7_port, ZN => n1900);
   U2405 : OAI221_X1 port map( B1 => n210, B2 => n1485, C1 => n526, C2 => n1486
                           , A => n1901, ZN => n1896);
   U2406 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_7_port, B1 => 
                           n1489, B2 => registers_6_7_port, ZN => n1901);
   U2407 : OAI221_X1 port map( B1 => n144, B2 => n1490, C1 => n400, C2 => n1491
                           , A => n1902, ZN => n1895);
   U2408 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_7_port, B1 => 
                           n1494, B2 => registers_14_7_port, ZN => n1902);
   U2409 : NAND4_X1 port map( A1 => n1903, A2 => n1904, A3 => n1905, A4 => 
                           n1906, ZN => n2957);
   U2410 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_6_port, C1 => 
                           n1449, C2 => registers_9_6_port, A => n1907, ZN => 
                           n1906);
   U2411 : OAI222_X1 port map( A1 => n465, A2 => n1451, B1 => n51, B2 => n1452,
                           C1 => n275, C2 => n1453, ZN => n1907);
   U2412 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_6_port, C1 => 
                           n1455, C2 => registers_20_6_port, A => n1908, ZN => 
                           n1905);
   U2413 : OAI22_X1 port map( A1 => n90, A2 => n1457, B1 => n315, B2 => n1458, 
                           ZN => n1908);
   U2414 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_6_port, C1 => 
                           n1460, C2 => registers_30_6_port, A => n1909, ZN => 
                           n1904);
   U2415 : OAI222_X1 port map( A1 => n466, A2 => n1462, B1 => n52, B2 => n1463,
                           C1 => n276, C2 => n1464, ZN => n1909);
   U2416 : AOI221_X1 port map( B1 => n1465, B2 => d_in(6), C1 => n1466, C2 => 
                           d_out1_6_port, A => n1910, ZN => n1903);
   U2417 : OAI22_X1 port map( A1 => n1911, A2 => n1469, B1 => n346, B2 => n1470
                           , ZN => n1910);
   U2418 : NOR4_X1 port map( A1 => n1912, A2 => n1913, A3 => n1914, A4 => n1915
                           , ZN => n1911);
   U2419 : OAI221_X1 port map( B1 => n145, B2 => n1475, C1 => n401, C2 => n1476
                           , A => n1916, ZN => n1915);
   U2420 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_6_port, B1 => 
                           n1479, B2 => registers_19_6_port, ZN => n1916);
   U2421 : OAI221_X1 port map( B1 => n211, B2 => n1480, C1 => n527, C2 => n1481
                           , A => n1917, ZN => n1914);
   U2422 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_6_port, B1 => 
                           n1484, B2 => registers_25_6_port, ZN => n1917);
   U2423 : OAI221_X1 port map( B1 => n212, B2 => n1485, C1 => n528, C2 => n1486
                           , A => n1918, ZN => n1913);
   U2424 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_6_port, B1 => 
                           n1489, B2 => registers_6_6_port, ZN => n1918);
   U2425 : OAI221_X1 port map( B1 => n146, B2 => n1490, C1 => n402, C2 => n1491
                           , A => n1919, ZN => n1912);
   U2426 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_6_port, B1 => 
                           n1494, B2 => registers_14_6_port, ZN => n1919);
   U2427 : NAND4_X1 port map( A1 => n1920, A2 => n1921, A3 => n1922, A4 => 
                           n1923, ZN => n2956);
   U2428 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_5_port, C1 => 
                           n1449, C2 => registers_9_5_port, A => n1924, ZN => 
                           n1923);
   U2429 : OAI222_X1 port map( A1 => n467, A2 => n1451, B1 => n53, B2 => n1452,
                           C1 => n277, C2 => n1453, ZN => n1924);
   U2430 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_5_port, C1 => 
                           n1455, C2 => registers_20_5_port, A => n1925, ZN => 
                           n1922);
   U2431 : OAI22_X1 port map( A1 => n91, A2 => n1457, B1 => n316, B2 => n1458, 
                           ZN => n1925);
   U2432 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_5_port, C1 => 
                           n1460, C2 => registers_30_5_port, A => n1926, ZN => 
                           n1921);
   U2433 : OAI222_X1 port map( A1 => n468, A2 => n1462, B1 => n54, B2 => n1463,
                           C1 => n278, C2 => n1464, ZN => n1926);
   U2434 : AOI221_X1 port map( B1 => n1465, B2 => d_in(5), C1 => n1466, C2 => 
                           d_out1_5_port, A => n1927, ZN => n1920);
   U2435 : OAI22_X1 port map( A1 => n1928, A2 => n1469, B1 => n347, B2 => n1470
                           , ZN => n1927);
   U2436 : NOR4_X1 port map( A1 => n1929, A2 => n1930, A3 => n1931, A4 => n1932
                           , ZN => n1928);
   U2437 : OAI221_X1 port map( B1 => n147, B2 => n1475, C1 => n403, C2 => n1476
                           , A => n1933, ZN => n1932);
   U2438 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_5_port, B1 => 
                           n1479, B2 => registers_19_5_port, ZN => n1933);
   U2439 : OAI221_X1 port map( B1 => n213, B2 => n1480, C1 => n529, C2 => n1481
                           , A => n1934, ZN => n1931);
   U2440 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_5_port, B1 => 
                           n1484, B2 => registers_25_5_port, ZN => n1934);
   U2441 : OAI221_X1 port map( B1 => n214, B2 => n1485, C1 => n530, C2 => n1486
                           , A => n1935, ZN => n1930);
   U2442 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_5_port, B1 => 
                           n1489, B2 => registers_6_5_port, ZN => n1935);
   U2443 : OAI221_X1 port map( B1 => n148, B2 => n1490, C1 => n404, C2 => n1491
                           , A => n1936, ZN => n1929);
   U2444 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_5_port, B1 => 
                           n1494, B2 => registers_14_5_port, ZN => n1936);
   U2445 : NAND4_X1 port map( A1 => n1937, A2 => n1938, A3 => n1939, A4 => 
                           n1940, ZN => n2955);
   U2446 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_4_port, C1 => 
                           n1449, C2 => registers_9_4_port, A => n1941, ZN => 
                           n1940);
   U2447 : OAI222_X1 port map( A1 => n469, A2 => n1451, B1 => n55, B2 => n1452,
                           C1 => n279, C2 => n1453, ZN => n1941);
   U2448 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_4_port, C1 => 
                           n1455, C2 => registers_20_4_port, A => n1942, ZN => 
                           n1939);
   U2449 : OAI22_X1 port map( A1 => n92, A2 => n1457, B1 => n317, B2 => n1458, 
                           ZN => n1942);
   U2450 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_4_port, C1 => 
                           n1460, C2 => registers_30_4_port, A => n1943, ZN => 
                           n1938);
   U2451 : OAI222_X1 port map( A1 => n470, A2 => n1462, B1 => n56, B2 => n1463,
                           C1 => n280, C2 => n1464, ZN => n1943);
   U2452 : AOI221_X1 port map( B1 => n1465, B2 => d_in(4), C1 => n1466, C2 => 
                           d_out1_4_port, A => n1944, ZN => n1937);
   U2453 : OAI22_X1 port map( A1 => n1945, A2 => n1469, B1 => n348, B2 => n1470
                           , ZN => n1944);
   U2454 : NOR4_X1 port map( A1 => n1946, A2 => n1947, A3 => n1948, A4 => n1949
                           , ZN => n1945);
   U2455 : OAI221_X1 port map( B1 => n149, B2 => n1475, C1 => n405, C2 => n1476
                           , A => n1950, ZN => n1949);
   U2456 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_4_port, B1 => 
                           n1479, B2 => registers_19_4_port, ZN => n1950);
   U2457 : OAI221_X1 port map( B1 => n215, B2 => n1480, C1 => n531, C2 => n1481
                           , A => n1951, ZN => n1948);
   U2458 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_4_port, B1 => 
                           n1484, B2 => registers_25_4_port, ZN => n1951);
   U2459 : OAI221_X1 port map( B1 => n216, B2 => n1485, C1 => n532, C2 => n1486
                           , A => n1952, ZN => n1947);
   U2460 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_4_port, B1 => 
                           n1489, B2 => registers_6_4_port, ZN => n1952);
   U2461 : OAI221_X1 port map( B1 => n150, B2 => n1490, C1 => n406, C2 => n1491
                           , A => n1953, ZN => n1946);
   U2462 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_4_port, B1 => 
                           n1494, B2 => registers_14_4_port, ZN => n1953);
   U2463 : NAND4_X1 port map( A1 => n1954, A2 => n1955, A3 => n1956, A4 => 
                           n1957, ZN => n2954);
   U2464 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_3_port, C1 => 
                           n1449, C2 => registers_9_3_port, A => n1958, ZN => 
                           n1957);
   U2465 : OAI222_X1 port map( A1 => n471, A2 => n1451, B1 => n57, B2 => n1452,
                           C1 => n281, C2 => n1453, ZN => n1958);
   U2466 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_3_port, C1 => 
                           n1455, C2 => registers_20_3_port, A => n1959, ZN => 
                           n1956);
   U2467 : OAI22_X1 port map( A1 => n93, A2 => n1457, B1 => n318, B2 => n1458, 
                           ZN => n1959);
   U2468 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_3_port, C1 => 
                           n1460, C2 => registers_30_3_port, A => n1960, ZN => 
                           n1955);
   U2469 : OAI222_X1 port map( A1 => n472, A2 => n1462, B1 => n58, B2 => n1463,
                           C1 => n282, C2 => n1464, ZN => n1960);
   U2470 : AOI221_X1 port map( B1 => n1465, B2 => d_in(3), C1 => n1466, C2 => 
                           d_out1_3_port, A => n1961, ZN => n1954);
   U2471 : OAI22_X1 port map( A1 => n1962, A2 => n1469, B1 => n349, B2 => n1470
                           , ZN => n1961);
   U2472 : NOR4_X1 port map( A1 => n1963, A2 => n1964, A3 => n1965, A4 => n1966
                           , ZN => n1962);
   U2473 : OAI221_X1 port map( B1 => n151, B2 => n1475, C1 => n407, C2 => n1476
                           , A => n1967, ZN => n1966);
   U2474 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_3_port, B1 => 
                           n1479, B2 => registers_19_3_port, ZN => n1967);
   U2475 : OAI221_X1 port map( B1 => n217, B2 => n1480, C1 => n533, C2 => n1481
                           , A => n1968, ZN => n1965);
   U2476 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_3_port, B1 => 
                           n1484, B2 => registers_25_3_port, ZN => n1968);
   U2477 : OAI221_X1 port map( B1 => n218, B2 => n1485, C1 => n534, C2 => n1486
                           , A => n1969, ZN => n1964);
   U2478 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_3_port, B1 => 
                           n1489, B2 => registers_6_3_port, ZN => n1969);
   U2479 : OAI221_X1 port map( B1 => n152, B2 => n1490, C1 => n408, C2 => n1491
                           , A => n1970, ZN => n1963);
   U2480 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_3_port, B1 => 
                           n1494, B2 => registers_14_3_port, ZN => n1970);
   U2481 : NAND4_X1 port map( A1 => n1971, A2 => n1972, A3 => n1973, A4 => 
                           n1974, ZN => n2953);
   U2482 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_2_port, C1 => 
                           n1449, C2 => registers_9_2_port, A => n1975, ZN => 
                           n1974);
   U2483 : OAI222_X1 port map( A1 => n473, A2 => n1451, B1 => n59, B2 => n1452,
                           C1 => n283, C2 => n1453, ZN => n1975);
   U2484 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_2_port, C1 => 
                           n1455, C2 => registers_20_2_port, A => n1976, ZN => 
                           n1973);
   U2485 : OAI22_X1 port map( A1 => n94, A2 => n1457, B1 => n319, B2 => n1458, 
                           ZN => n1976);
   U2486 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_2_port, C1 => 
                           n1460, C2 => registers_30_2_port, A => n1977, ZN => 
                           n1972);
   U2487 : OAI222_X1 port map( A1 => n474, A2 => n1462, B1 => n60, B2 => n1463,
                           C1 => n284, C2 => n1464, ZN => n1977);
   U2488 : AOI221_X1 port map( B1 => n1465, B2 => d_in(2), C1 => n1466, C2 => 
                           d_out1_2_port, A => n1978, ZN => n1971);
   U2489 : OAI22_X1 port map( A1 => n1979, A2 => n1469, B1 => n350, B2 => n1470
                           , ZN => n1978);
   U2490 : NOR4_X1 port map( A1 => n1980, A2 => n1981, A3 => n1982, A4 => n1983
                           , ZN => n1979);
   U2491 : OAI221_X1 port map( B1 => n153, B2 => n1475, C1 => n409, C2 => n1476
                           , A => n1984, ZN => n1983);
   U2492 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_2_port, B1 => 
                           n1479, B2 => registers_19_2_port, ZN => n1984);
   U2493 : OAI221_X1 port map( B1 => n219, B2 => n1480, C1 => n535, C2 => n1481
                           , A => n1985, ZN => n1982);
   U2494 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_2_port, B1 => 
                           n1484, B2 => registers_25_2_port, ZN => n1985);
   U2495 : OAI221_X1 port map( B1 => n220, B2 => n1485, C1 => n536, C2 => n1486
                           , A => n1986, ZN => n1981);
   U2496 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_2_port, B1 => 
                           n1489, B2 => registers_6_2_port, ZN => n1986);
   U2497 : OAI221_X1 port map( B1 => n154, B2 => n1490, C1 => n410, C2 => n1491
                           , A => n1987, ZN => n1980);
   U2498 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_2_port, B1 => 
                           n1494, B2 => registers_14_2_port, ZN => n1987);
   U2499 : NAND4_X1 port map( A1 => n1988, A2 => n1989, A3 => n1990, A4 => 
                           n1991, ZN => n2952);
   U2500 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_1_port, C1 => 
                           n1449, C2 => registers_9_1_port, A => n1992, ZN => 
                           n1991);
   U2501 : OAI222_X1 port map( A1 => n475, A2 => n1451, B1 => n61, B2 => n1452,
                           C1 => n285, C2 => n1453, ZN => n1992);
   U2502 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_1_port, C1 => 
                           n1455, C2 => registers_20_1_port, A => n1993, ZN => 
                           n1990);
   U2503 : OAI22_X1 port map( A1 => n95, A2 => n1457, B1 => n320, B2 => n1458, 
                           ZN => n1993);
   U2504 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_1_port, C1 => 
                           n1460, C2 => registers_30_1_port, A => n1994, ZN => 
                           n1989);
   U2505 : OAI222_X1 port map( A1 => n476, A2 => n1462, B1 => n62, B2 => n1463,
                           C1 => n286, C2 => n1464, ZN => n1994);
   U2506 : AOI221_X1 port map( B1 => n1465, B2 => d_in(1), C1 => n1466, C2 => 
                           d_out1_1_port, A => n1995, ZN => n1988);
   U2507 : OAI22_X1 port map( A1 => n1996, A2 => n1469, B1 => n351, B2 => n1470
                           , ZN => n1995);
   U2508 : NOR4_X1 port map( A1 => n1997, A2 => n1998, A3 => n1999, A4 => n2000
                           , ZN => n1996);
   U2509 : OAI221_X1 port map( B1 => n155, B2 => n1475, C1 => n411, C2 => n1476
                           , A => n2001, ZN => n2000);
   U2510 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_1_port, B1 => 
                           n1479, B2 => registers_19_1_port, ZN => n2001);
   U2511 : OAI221_X1 port map( B1 => n221, B2 => n1480, C1 => n537, C2 => n1481
                           , A => n2002, ZN => n1999);
   U2512 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_1_port, B1 => 
                           n1484, B2 => registers_25_1_port, ZN => n2002);
   U2513 : OAI221_X1 port map( B1 => n222, B2 => n1485, C1 => n538, C2 => n1486
                           , A => n2003, ZN => n1998);
   U2514 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_1_port, B1 => 
                           n1489, B2 => registers_6_1_port, ZN => n2003);
   U2515 : OAI221_X1 port map( B1 => n156, B2 => n1490, C1 => n412, C2 => n1491
                           , A => n2004, ZN => n1997);
   U2516 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_1_port, B1 => 
                           n1494, B2 => registers_14_1_port, ZN => n2004);
   U2517 : NAND4_X1 port map( A1 => n2005, A2 => n2006, A3 => n2007, A4 => 
                           n2008, ZN => n2951);
   U2518 : AOI221_X1 port map( B1 => n1448, B2 => registers_12_0_port, C1 => 
                           n1449, C2 => registers_9_0_port, A => n2009, ZN => 
                           n2008);
   U2519 : OAI222_X1 port map( A1 => n477, A2 => n1451, B1 => n63, B2 => n1452,
                           C1 => n287, C2 => n1453, ZN => n2009);
   U2520 : AOI221_X1 port map( B1 => n1454, B2 => registers_4_0_port, C1 => 
                           n1455, C2 => registers_20_0_port, A => n2016, ZN => 
                           n2007);
   U2521 : OAI22_X1 port map( A1 => n96, A2 => n1457, B1 => n321, B2 => n1458, 
                           ZN => n2016);
   U2522 : AND2_X1 port map( A1 => n2018, A2 => n2019, ZN => n2011);
   U2523 : AOI221_X1 port map( B1 => n1459, B2 => registers_15_0_port, C1 => 
                           n1460, C2 => registers_30_0_port, A => n2021, ZN => 
                           n2006);
   U2524 : OAI222_X1 port map( A1 => n478, A2 => n1462, B1 => n64, B2 => n1463,
                           C1 => n288, C2 => n1464, ZN => n2021);
   U2525 : AND2_X1 port map( A1 => n2022, A2 => n2019, ZN => n2014);
   U2526 : AOI221_X1 port map( B1 => n1465, B2 => d_in(0), C1 => n1466, C2 => 
                           d_out1_0_port, A => n2027, ZN => n2005);
   U2527 : OAI22_X1 port map( A1 => n2028, A2 => n1469, B1 => n352, B2 => n1470
                           , ZN => n2027);
   U2528 : INV_X1 port map( A => n1469, ZN => n2019);
   U2529 : INV_X1 port map( A => n1466, ZN => n2029);
   U2530 : NOR4_X1 port map( A1 => n2031, A2 => n2032, A3 => n2033, A4 => n2034
                           , ZN => n2028);
   U2531 : OAI221_X1 port map( B1 => n157, B2 => n1475, C1 => n413, C2 => n1476
                           , A => n2035, ZN => n2034);
   U2532 : AOI22_X1 port map( A1 => n1478, A2 => registers_22_0_port, B1 => 
                           n1479, B2 => registers_19_0_port, ZN => n2035);
   U2533 : NOR3_X1 port map( A1 => rd1_addr(0), A2 => rd1_addr(3), A3 => n2036,
                           ZN => n2010);
   U2534 : OAI221_X1 port map( B1 => n223, B2 => n1480, C1 => n539, C2 => n1481
                           , A => n2037, ZN => n2033);
   U2535 : AOI22_X1 port map( A1 => n1483, A2 => registers_28_0_port, B1 => 
                           n1484, B2 => registers_25_0_port, ZN => n2037);
   U2536 : NOR3_X1 port map( A1 => n2038, A2 => rd1_addr(3), A3 => n2036, ZN =>
                           n2012);
   U2537 : NOR2_X1 port map( A1 => rd1_addr(1), A2 => rd1_addr(2), ZN => n2018)
                           ;
   U2538 : NOR3_X1 port map( A1 => n2036, A2 => rd1_addr(0), A3 => n2039, ZN =>
                           n2023);
   U2539 : OAI221_X1 port map( B1 => n224, B2 => n1485, C1 => n540, C2 => n1486
                           , A => n2040, ZN => n2032);
   U2540 : AOI22_X1 port map( A1 => n1488, A2 => registers_3_0_port, B1 => 
                           n1489, B2 => registers_6_0_port, ZN => n2040);
   U2541 : NOR3_X1 port map( A1 => rd1_addr(3), A2 => rd1_addr(4), A3 => 
                           rd1_addr(0), ZN => n2020);
   U2542 : NOR2_X1 port map( A1 => n2041, A2 => rd1_addr(1), ZN => n2022);
   U2543 : NOR3_X1 port map( A1 => n2036, A2 => n2038, A3 => n2039, ZN => n2025
                           );
   U2544 : OAI221_X1 port map( B1 => n158, B2 => n1490, C1 => n414, C2 => n1491
                           , A => n2042, ZN => n2031);
   U2545 : AOI22_X1 port map( A1 => n1493, A2 => registers_11_0_port, B1 => 
                           n1494, B2 => registers_14_0_port, ZN => n2042);
   U2546 : NOR3_X1 port map( A1 => n2038, A2 => rd1_addr(4), A3 => n2039, ZN =>
                           n2013);
   U2547 : NOR3_X1 port map( A1 => rd1_addr(0), A2 => rd1_addr(4), A3 => n2039,
                           ZN => n2015);
   U2548 : NOR2_X1 port map( A1 => n2043, A2 => rd1_addr(2), ZN => n2024);
   U2549 : NOR3_X1 port map( A1 => rd1_addr(3), A2 => rd1_addr(4), A3 => n2038,
                           ZN => n2017);
   U2550 : INV_X1 port map( A => rd1_addr(0), ZN => n2038);
   U2551 : NOR2_X1 port map( A1 => n2041, A2 => n2043, ZN => n2026);
   U2552 : INV_X1 port map( A => rd1_addr(1), ZN => n2043);
   U2553 : NAND4_X1 port map( A1 => n2044, A2 => n2045, A3 => n2046, A4 => 
                           n2047, ZN => n2030);
   U2554 : NOR3_X1 port map( A1 => n2048, A2 => n684, A3 => n2049, ZN => n2047)
                           ;
   U2555 : XOR2_X1 port map( A => wr_addr(1), B => rd1_addr(1), Z => n2049);
   U2556 : INV_X1 port map( A => wr_en, ZN => n684);
   U2557 : XOR2_X1 port map( A => wr_addr(0), B => rd1_addr(0), Z => n2048);
   U2558 : XOR2_X1 port map( A => n2039, B => wr_addr(3), Z => n2046);
   U2559 : INV_X1 port map( A => rd1_addr(3), ZN => n2039);
   U2560 : XOR2_X1 port map( A => wr_addr(4), B => n2036, Z => n2045);
   U2561 : INV_X1 port map( A => rd1_addr(4), ZN => n2036);
   U2562 : XOR2_X1 port map( A => n2041, B => wr_addr(2), Z => n2044);
   U2563 : INV_X1 port map( A => rd1_addr(2), ZN => n2041);
   U2564 : INV_X1 port map( A => clk, ZN => N18);

end SYN_register_file_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Extender_SRC_SIZE26_DEST_SIZE32 is

   port( s : in std_logic;  i : in std_logic_vector (25 downto 0);  o : out 
         std_logic_vector (31 downto 0));

end Extender_SRC_SIZE26_DEST_SIZE32;

architecture SYN_extender_arch of Extender_SRC_SIZE26_DEST_SIZE32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal o_31 : std_logic;

begin
   o <= ( o_31, o_31, o_31, o_31, o_31, o_31, i(25), i(24), i(23), i(22), i(21)
      , i(20), i(19), i(18), i(17), i(16), i(15), i(14), i(13), i(12), i(11), 
      i(10), i(9), i(8), i(7), i(6), i(5), i(4), i(3), i(2), i(1), i(0) );
   
   U1 : AND2_X1 port map( A1 => s, A2 => i(25), ZN => o_31);

end SYN_extender_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Extender_SRC_SIZE16_DEST_SIZE32 is

   port( s : in std_logic;  i : in std_logic_vector (15 downto 0);  o : out 
         std_logic_vector (31 downto 0));

end Extender_SRC_SIZE16_DEST_SIZE32;

architecture SYN_extender_arch of Extender_SRC_SIZE16_DEST_SIZE32 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal o_31 : std_logic;

begin
   o <= ( o_31, o_31, o_31, o_31, o_31, o_31, o_31, o_31, o_31, o_31, o_31, 
      o_31, o_31, o_31, o_31, o_31, i(15), i(14), i(13), i(12), i(11), i(10), 
      i(9), i(8), i(7), i(6), i(5), i(4), i(3), i(2), i(1), i(0) );
   
   U1 : AND2_X1 port map( A1 => s, A2 => i(15), ZN => o_31);

end SYN_extender_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE5 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (4 downto 0);  
         dout : out std_logic_vector (4 downto 0));

end Mux_DATA_SIZE5;

architecture SYN_mux_arch of Mux_DATA_SIZE5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(4), B => din1(4), S => sel, Z => dout(4));
   U2 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U3 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U4 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U5 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Reg_DATA_SIZE32_0 is

   port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 0);
         dout : out std_logic_vector (31 downto 0));

end Reg_DATA_SIZE32_0;

architecture SYN_reg_arch of Reg_DATA_SIZE32_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal dout_31_port, dout_30_port, dout_29_port, dout_28_port, dout_27_port,
      dout_26_port, dout_25_port, dout_24_port, dout_23_port, dout_22_port, 
      dout_21_port, dout_20_port, dout_19_port, dout_18_port, dout_17_port, 
      dout_16_port, dout_15_port, dout_14_port, dout_13_port, dout_12_port, 
      dout_11_port, dout_10_port, dout_9_port, dout_8_port, dout_7_port, 
      dout_6_port, dout_5_port, dout_4_port, dout_3_port, dout_2_port, 
      dout_1_port, dout_0_port, n65, n66, n67, n68, n69, n70, n71, n72, n73, 
      n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88
      , n89, n90, n91, n92, n93, n94, n95, n96, net108097, net108098, net108099
      , net108100, net108101, net108102, net108103, net108104, net108105, 
      net108106, net108107, net108108, net108109, net108110, net108111, 
      net108112, net108113, net108114, net108115, net108116, net108117, 
      net108118, net108119, net108120, net108121, net108122, net108123, 
      net108124, net108125, net108126, net108127, net108128 : std_logic;

begin
   dout <= ( dout_31_port, dout_30_port, dout_29_port, dout_28_port, 
      dout_27_port, dout_26_port, dout_25_port, dout_24_port, dout_23_port, 
      dout_22_port, dout_21_port, dout_20_port, dout_19_port, dout_18_port, 
      dout_17_port, dout_16_port, dout_15_port, dout_14_port, dout_13_port, 
      dout_12_port, dout_11_port, dout_10_port, dout_9_port, dout_8_port, 
      dout_7_port, dout_6_port, dout_5_port, dout_4_port, dout_3_port, 
      dout_2_port, dout_1_port, dout_0_port );
   
   dout_reg_31_inst : DFFR_X1 port map( D => n96, CK => clk, RN => rst, Q => 
                           dout_31_port, QN => net108128);
   dout_reg_30_inst : DFFR_X1 port map( D => n95, CK => clk, RN => rst, Q => 
                           dout_30_port, QN => net108127);
   dout_reg_29_inst : DFFR_X1 port map( D => n94, CK => clk, RN => rst, Q => 
                           dout_29_port, QN => net108126);
   dout_reg_28_inst : DFFR_X1 port map( D => n93, CK => clk, RN => rst, Q => 
                           dout_28_port, QN => net108125);
   dout_reg_27_inst : DFFR_X1 port map( D => n92, CK => clk, RN => rst, Q => 
                           dout_27_port, QN => net108124);
   dout_reg_26_inst : DFFR_X1 port map( D => n91, CK => clk, RN => rst, Q => 
                           dout_26_port, QN => net108123);
   dout_reg_25_inst : DFFR_X1 port map( D => n90, CK => clk, RN => rst, Q => 
                           dout_25_port, QN => net108122);
   dout_reg_24_inst : DFFR_X1 port map( D => n89, CK => clk, RN => rst, Q => 
                           dout_24_port, QN => net108121);
   dout_reg_23_inst : DFFR_X1 port map( D => n88, CK => clk, RN => rst, Q => 
                           dout_23_port, QN => net108120);
   dout_reg_22_inst : DFFR_X1 port map( D => n87, CK => clk, RN => rst, Q => 
                           dout_22_port, QN => net108119);
   dout_reg_21_inst : DFFR_X1 port map( D => n86, CK => clk, RN => rst, Q => 
                           dout_21_port, QN => net108118);
   dout_reg_20_inst : DFFR_X1 port map( D => n85, CK => clk, RN => rst, Q => 
                           dout_20_port, QN => net108117);
   dout_reg_19_inst : DFFR_X1 port map( D => n84, CK => clk, RN => rst, Q => 
                           dout_19_port, QN => net108116);
   dout_reg_18_inst : DFFR_X1 port map( D => n83, CK => clk, RN => rst, Q => 
                           dout_18_port, QN => net108115);
   dout_reg_17_inst : DFFR_X1 port map( D => n82, CK => clk, RN => rst, Q => 
                           dout_17_port, QN => net108114);
   dout_reg_16_inst : DFFR_X1 port map( D => n81, CK => clk, RN => rst, Q => 
                           dout_16_port, QN => net108113);
   dout_reg_15_inst : DFFR_X1 port map( D => n80, CK => clk, RN => rst, Q => 
                           dout_15_port, QN => net108112);
   dout_reg_14_inst : DFFR_X1 port map( D => n79, CK => clk, RN => rst, Q => 
                           dout_14_port, QN => net108111);
   dout_reg_13_inst : DFFR_X1 port map( D => n78, CK => clk, RN => rst, Q => 
                           dout_13_port, QN => net108110);
   dout_reg_12_inst : DFFR_X1 port map( D => n77, CK => clk, RN => rst, Q => 
                           dout_12_port, QN => net108109);
   dout_reg_11_inst : DFFR_X1 port map( D => n76, CK => clk, RN => rst, Q => 
                           dout_11_port, QN => net108108);
   dout_reg_10_inst : DFFR_X1 port map( D => n75, CK => clk, RN => rst, Q => 
                           dout_10_port, QN => net108107);
   dout_reg_9_inst : DFFR_X1 port map( D => n74, CK => clk, RN => rst, Q => 
                           dout_9_port, QN => net108106);
   dout_reg_8_inst : DFFR_X1 port map( D => n73, CK => clk, RN => rst, Q => 
                           dout_8_port, QN => net108105);
   dout_reg_7_inst : DFFR_X1 port map( D => n72, CK => clk, RN => rst, Q => 
                           dout_7_port, QN => net108104);
   dout_reg_6_inst : DFFR_X1 port map( D => n71, CK => clk, RN => rst, Q => 
                           dout_6_port, QN => net108103);
   dout_reg_5_inst : DFFR_X1 port map( D => n70, CK => clk, RN => rst, Q => 
                           dout_5_port, QN => net108102);
   dout_reg_4_inst : DFFR_X1 port map( D => n69, CK => clk, RN => rst, Q => 
                           dout_4_port, QN => net108101);
   dout_reg_3_inst : DFFR_X1 port map( D => n68, CK => clk, RN => rst, Q => 
                           dout_3_port, QN => net108100);
   dout_reg_2_inst : DFFR_X1 port map( D => n67, CK => clk, RN => rst, Q => 
                           dout_2_port, QN => net108099);
   dout_reg_1_inst : DFFR_X1 port map( D => n66, CK => clk, RN => rst, Q => 
                           dout_1_port, QN => net108098);
   dout_reg_0_inst : DFFR_X1 port map( D => n65, CK => clk, RN => rst, Q => 
                           dout_0_port, QN => net108097);
   U2 : MUX2_X1 port map( A => dout_31_port, B => din(31), S => en, Z => n96);
   U3 : MUX2_X1 port map( A => dout_30_port, B => din(30), S => en, Z => n95);
   U4 : MUX2_X1 port map( A => dout_29_port, B => din(29), S => en, Z => n94);
   U5 : MUX2_X1 port map( A => dout_28_port, B => din(28), S => en, Z => n93);
   U6 : MUX2_X1 port map( A => dout_27_port, B => din(27), S => en, Z => n92);
   U7 : MUX2_X1 port map( A => dout_26_port, B => din(26), S => en, Z => n91);
   U8 : MUX2_X1 port map( A => dout_25_port, B => din(25), S => en, Z => n90);
   U9 : MUX2_X1 port map( A => dout_24_port, B => din(24), S => en, Z => n89);
   U10 : MUX2_X1 port map( A => dout_23_port, B => din(23), S => en, Z => n88);
   U11 : MUX2_X1 port map( A => dout_22_port, B => din(22), S => en, Z => n87);
   U12 : MUX2_X1 port map( A => dout_21_port, B => din(21), S => en, Z => n86);
   U13 : MUX2_X1 port map( A => dout_20_port, B => din(20), S => en, Z => n85);
   U14 : MUX2_X1 port map( A => dout_19_port, B => din(19), S => en, Z => n84);
   U15 : MUX2_X1 port map( A => dout_18_port, B => din(18), S => en, Z => n83);
   U16 : MUX2_X1 port map( A => dout_17_port, B => din(17), S => en, Z => n82);
   U17 : MUX2_X1 port map( A => dout_16_port, B => din(16), S => en, Z => n81);
   U18 : MUX2_X1 port map( A => dout_15_port, B => din(15), S => en, Z => n80);
   U19 : MUX2_X1 port map( A => dout_14_port, B => din(14), S => en, Z => n79);
   U20 : MUX2_X1 port map( A => dout_13_port, B => din(13), S => en, Z => n78);
   U21 : MUX2_X1 port map( A => dout_12_port, B => din(12), S => en, Z => n77);
   U22 : MUX2_X1 port map( A => dout_11_port, B => din(11), S => en, Z => n76);
   U23 : MUX2_X1 port map( A => dout_10_port, B => din(10), S => en, Z => n75);
   U24 : MUX2_X1 port map( A => dout_9_port, B => din(9), S => en, Z => n74);
   U25 : MUX2_X1 port map( A => dout_8_port, B => din(8), S => en, Z => n73);
   U26 : MUX2_X1 port map( A => dout_7_port, B => din(7), S => en, Z => n72);
   U27 : MUX2_X1 port map( A => dout_6_port, B => din(6), S => en, Z => n71);
   U28 : MUX2_X1 port map( A => dout_5_port, B => din(5), S => en, Z => n70);
   U29 : MUX2_X1 port map( A => dout_4_port, B => din(4), S => en, Z => n69);
   U30 : MUX2_X1 port map( A => dout_3_port, B => din(3), S => en, Z => n68);
   U31 : MUX2_X1 port map( A => dout_2_port, B => din(2), S => en, Z => n67);
   U32 : MUX2_X1 port map( A => dout_1_port, B => din(1), S => en, Z => n66);
   U33 : MUX2_X1 port map( A => dout_0_port, B => din(0), S => en, Z => n65);

end SYN_reg_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Mux_DATA_SIZE32_0 is

   port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0);  
         dout : out std_logic_vector (31 downto 0));

end Mux_DATA_SIZE32_0;

architecture SYN_mux_arch of Mux_DATA_SIZE32_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => din0(9), B => din1(9), S => sel, Z => dout(9));
   U2 : MUX2_X1 port map( A => din0(8), B => din1(8), S => sel, Z => dout(8));
   U3 : MUX2_X1 port map( A => din0(7), B => din1(7), S => sel, Z => dout(7));
   U4 : MUX2_X1 port map( A => din0(6), B => din1(6), S => sel, Z => dout(6));
   U5 : MUX2_X1 port map( A => din0(5), B => din1(5), S => sel, Z => dout(5));
   U6 : MUX2_X1 port map( A => din0(4), B => din1(4), S => sel, Z => dout(4));
   U7 : MUX2_X1 port map( A => din0(3), B => din1(3), S => sel, Z => dout(3));
   U8 : MUX2_X1 port map( A => din0(31), B => din1(31), S => sel, Z => dout(31)
                           );
   U9 : MUX2_X1 port map( A => din0(30), B => din1(30), S => sel, Z => dout(30)
                           );
   U10 : MUX2_X1 port map( A => din0(2), B => din1(2), S => sel, Z => dout(2));
   U11 : MUX2_X1 port map( A => din0(29), B => din1(29), S => sel, Z => 
                           dout(29));
   U12 : MUX2_X1 port map( A => din0(28), B => din1(28), S => sel, Z => 
                           dout(28));
   U13 : MUX2_X1 port map( A => din0(27), B => din1(27), S => sel, Z => 
                           dout(27));
   U14 : MUX2_X1 port map( A => din0(26), B => din1(26), S => sel, Z => 
                           dout(26));
   U15 : MUX2_X1 port map( A => din0(25), B => din1(25), S => sel, Z => 
                           dout(25));
   U16 : MUX2_X1 port map( A => din0(24), B => din1(24), S => sel, Z => 
                           dout(24));
   U17 : MUX2_X1 port map( A => din0(23), B => din1(23), S => sel, Z => 
                           dout(23));
   U18 : MUX2_X1 port map( A => din0(22), B => din1(22), S => sel, Z => 
                           dout(22));
   U19 : MUX2_X1 port map( A => din0(21), B => din1(21), S => sel, Z => 
                           dout(21));
   U20 : MUX2_X1 port map( A => din0(20), B => din1(20), S => sel, Z => 
                           dout(20));
   U21 : MUX2_X1 port map( A => din0(1), B => din1(1), S => sel, Z => dout(1));
   U22 : MUX2_X1 port map( A => din0(19), B => din1(19), S => sel, Z => 
                           dout(19));
   U23 : MUX2_X1 port map( A => din0(18), B => din1(18), S => sel, Z => 
                           dout(18));
   U24 : MUX2_X1 port map( A => din0(17), B => din1(17), S => sel, Z => 
                           dout(17));
   U25 : MUX2_X1 port map( A => din0(16), B => din1(16), S => sel, Z => 
                           dout(16));
   U26 : MUX2_X1 port map( A => din0(15), B => din1(15), S => sel, Z => 
                           dout(15));
   U27 : MUX2_X1 port map( A => din0(14), B => din1(14), S => sel, Z => 
                           dout(14));
   U28 : MUX2_X1 port map( A => din0(13), B => din1(13), S => sel, Z => 
                           dout(13));
   U29 : MUX2_X1 port map( A => din0(12), B => din1(12), S => sel, Z => 
                           dout(12));
   U30 : MUX2_X1 port map( A => din0(11), B => din1(11), S => sel, Z => 
                           dout(11));
   U31 : MUX2_X1 port map( A => din0(10), B => din1(10), S => sel, Z => 
                           dout(10));
   U32 : MUX2_X1 port map( A => din0(0), B => din1(0), S => sel, Z => dout(0));

end SYN_mux_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Adder_DATA_SIZE32_0 is

   port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s : 
         out std_logic_vector (31 downto 0);  cout : out std_logic);

end Adder_DATA_SIZE32_0;

architecture SYN_adder_arch of Adder_DATA_SIZE32_0 is

   component P4Adder_DATA_SIZE32_SPARSITY4_0
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;

begin
   
   ADDER0 : P4Adder_DATA_SIZE32_SPARSITY4_0 port map( cin => cin, a(31) => 
                           a(31), a(30) => a(30), a(29) => a(29), a(28) => 
                           a(28), a(27) => a(27), a(26) => a(26), a(25) => 
                           a(25), a(24) => a(24), a(23) => a(23), a(22) => 
                           a(22), a(21) => a(21), a(20) => a(20), a(19) => 
                           a(19), a(18) => a(18), a(17) => a(17), a(16) => 
                           a(16), a(15) => a(15), a(14) => a(14), a(13) => 
                           a(13), a(12) => a(12), a(11) => a(11), a(10) => 
                           a(10), a(9) => a(9), a(8) => a(8), a(7) => a(7), 
                           a(6) => a(6), a(5) => a(5), a(4) => a(4), a(3) => 
                           a(3), a(2) => a(2), a(1) => a(1), a(0) => a(0), 
                           b(31) => b(31), b(30) => b(30), b(29) => b(29), 
                           b(28) => b(28), b(27) => b(27), b(26) => b(26), 
                           b(25) => b(25), b(24) => b(24), b(23) => b(23), 
                           b(22) => b(22), b(21) => b(21), b(20) => b(20), 
                           b(19) => b(19), b(18) => b(18), b(17) => b(17), 
                           b(16) => b(16), b(15) => b(15), b(14) => b(14), 
                           b(13) => b(13), b(12) => b(12), b(11) => b(11), 
                           b(10) => b(10), b(9) => b(9), b(8) => b(8), b(7) => 
                           b(7), b(6) => b(6), b(5) => b(5), b(4) => b(4), b(3)
                           => b(3), b(2) => b(2), b(1) => b(1), b(0) => b(0), 
                           s(31) => s(31), s(30) => s(30), s(29) => s(29), 
                           s(28) => s(28), s(27) => s(27), s(26) => s(26), 
                           s(25) => s(25), s(24) => s(24), s(23) => s(23), 
                           s(22) => s(22), s(21) => s(21), s(20) => s(20), 
                           s(19) => s(19), s(18) => s(18), s(17) => s(17), 
                           s(16) => s(16), s(15) => s(15), s(14) => s(14), 
                           s(13) => s(13), s(12) => s(12), s(11) => s(11), 
                           s(10) => s(10), s(9) => s(9), s(8) => s(8), s(7) => 
                           s(7), s(6) => s(6), s(5) => s(5), s(4) => s(4), s(3)
                           => s(3), s(2) => s(2), s(1) => s(1), s(0) => s(0), 
                           cout => cout);

end SYN_adder_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Branch_DATA_SIZE32_OPCD_SIZE6_ADDR_SIZE32 is

   port( rst, clk : in std_logic;  reg_a, ld_a : in std_logic_vector (31 downto
         0);  opcd : in std_logic_vector (5 downto 0);  addr : in 
         std_logic_vector (31 downto 0);  sig_bal : in std_logic;  sig_bpw, 
         sig_brt : out std_logic);

end Branch_DATA_SIZE32_OPCD_SIZE6_ADDR_SIZE32;

architecture SYN_branch_arch of Branch_DATA_SIZE32_OPCD_SIZE6_ADDR_SIZE32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X2
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X4
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal sig_brt_tmp, bht_0_26_port, bht_0_25_port, bht_0_24_port, 
      bht_0_23_port, bht_0_22_port, bht_0_21_port, bht_0_20_port, bht_0_19_port
      , bht_0_18_port, bht_0_17_port, bht_0_16_port, bht_0_15_port, 
      bht_0_14_port, bht_0_13_port, bht_0_12_port, bht_0_11_port, bht_0_10_port
      , bht_0_9_port, bht_0_8_port, bht_0_7_port, bht_0_6_port, bht_0_5_port, 
      bht_0_4_port, bht_0_3_port, bht_0_2_port, bht_0_1_port, bht_0_0_port, 
      bht_1_26_port, bht_1_25_port, bht_1_24_port, bht_1_23_port, bht_1_22_port
      , bht_1_21_port, bht_1_20_port, bht_1_19_port, bht_1_18_port, 
      bht_1_17_port, bht_1_16_port, bht_1_15_port, bht_1_14_port, bht_1_13_port
      , bht_1_12_port, bht_1_11_port, bht_1_10_port, bht_1_9_port, bht_1_8_port
      , bht_1_7_port, bht_1_6_port, bht_1_5_port, bht_1_4_port, bht_1_3_port, 
      bht_1_2_port, bht_1_1_port, bht_1_0_port, bht_2_26_port, bht_2_25_port, 
      bht_2_24_port, bht_2_23_port, bht_2_22_port, bht_2_21_port, bht_2_20_port
      , bht_2_19_port, bht_2_18_port, bht_2_17_port, bht_2_16_port, 
      bht_2_15_port, bht_2_14_port, bht_2_13_port, bht_2_12_port, bht_2_11_port
      , bht_2_10_port, bht_2_9_port, bht_2_8_port, bht_2_7_port, bht_2_6_port, 
      bht_2_5_port, bht_2_4_port, bht_2_3_port, bht_2_2_port, bht_2_1_port, 
      bht_2_0_port, bht_3_26_port, bht_3_25_port, bht_3_24_port, bht_3_23_port,
      bht_3_22_port, bht_3_21_port, bht_3_20_port, bht_3_19_port, bht_3_18_port
      , bht_3_17_port, bht_3_16_port, bht_3_15_port, bht_3_14_port, 
      bht_3_13_port, bht_3_12_port, bht_3_11_port, bht_3_10_port, bht_3_9_port,
      bht_3_8_port, bht_3_7_port, bht_3_6_port, bht_3_5_port, bht_3_4_port, 
      bht_3_3_port, bht_3_2_port, bht_3_1_port, bht_3_0_port, bht_4_26_port, 
      bht_4_25_port, bht_4_24_port, bht_4_23_port, bht_4_22_port, bht_4_21_port
      , bht_4_20_port, bht_4_19_port, bht_4_18_port, bht_4_17_port, 
      bht_4_16_port, bht_4_15_port, bht_4_14_port, bht_4_13_port, bht_4_12_port
      , bht_4_11_port, bht_4_10_port, bht_4_9_port, bht_4_8_port, bht_4_7_port,
      bht_4_6_port, bht_4_5_port, bht_4_4_port, bht_4_3_port, bht_4_2_port, 
      bht_4_1_port, bht_4_0_port, bht_5_26_port, bht_5_25_port, bht_5_24_port, 
      bht_5_23_port, bht_5_22_port, bht_5_21_port, bht_5_20_port, bht_5_19_port
      , bht_5_18_port, bht_5_17_port, bht_5_16_port, bht_5_15_port, 
      bht_5_14_port, bht_5_13_port, bht_5_12_port, bht_5_11_port, bht_5_10_port
      , bht_5_9_port, bht_5_8_port, bht_5_7_port, bht_5_6_port, bht_5_5_port, 
      bht_5_4_port, bht_5_3_port, bht_5_2_port, bht_5_1_port, bht_5_0_port, 
      bht_6_26_port, bht_6_25_port, bht_6_24_port, bht_6_23_port, bht_6_22_port
      , bht_6_21_port, bht_6_20_port, bht_6_19_port, bht_6_18_port, 
      bht_6_17_port, bht_6_16_port, bht_6_15_port, bht_6_14_port, bht_6_13_port
      , bht_6_12_port, bht_6_11_port, bht_6_10_port, bht_6_9_port, bht_6_8_port
      , bht_6_7_port, bht_6_6_port, bht_6_5_port, bht_6_4_port, bht_6_3_port, 
      bht_6_2_port, bht_6_1_port, bht_6_0_port, bht_7_26_port, bht_7_25_port, 
      bht_7_24_port, bht_7_23_port, bht_7_22_port, bht_7_21_port, bht_7_20_port
      , bht_7_19_port, bht_7_18_port, bht_7_17_port, bht_7_16_port, 
      bht_7_15_port, bht_7_14_port, bht_7_13_port, bht_7_12_port, bht_7_11_port
      , bht_7_10_port, bht_7_9_port, bht_7_8_port, bht_7_7_port, bht_7_6_port, 
      bht_7_5_port, bht_7_4_port, bht_7_3_port, bht_7_2_port, bht_7_1_port, 
      bht_7_0_port, bht_8_26_port, bht_8_25_port, bht_8_24_port, bht_8_23_port,
      bht_8_22_port, bht_8_21_port, bht_8_20_port, bht_8_19_port, bht_8_18_port
      , bht_8_17_port, bht_8_16_port, bht_8_15_port, bht_8_14_port, 
      bht_8_13_port, bht_8_12_port, bht_8_11_port, bht_8_10_port, bht_8_9_port,
      bht_8_8_port, bht_8_7_port, bht_8_6_port, bht_8_5_port, bht_8_4_port, 
      bht_8_3_port, bht_8_2_port, bht_8_1_port, bht_8_0_port, bht_9_26_port, 
      bht_9_25_port, bht_9_24_port, bht_9_23_port, bht_9_22_port, bht_9_21_port
      , bht_9_20_port, bht_9_19_port, bht_9_18_port, bht_9_17_port, 
      bht_9_16_port, bht_9_15_port, bht_9_14_port, bht_9_13_port, bht_9_12_port
      , bht_9_11_port, bht_9_10_port, bht_9_9_port, bht_9_8_port, bht_9_7_port,
      bht_9_6_port, bht_9_5_port, bht_9_4_port, bht_9_3_port, bht_9_2_port, 
      bht_9_1_port, bht_9_0_port, bht_10_26_port, bht_10_25_port, 
      bht_10_24_port, bht_10_23_port, bht_10_22_port, bht_10_21_port, 
      bht_10_20_port, bht_10_19_port, bht_10_18_port, bht_10_17_port, 
      bht_10_16_port, bht_10_15_port, bht_10_14_port, bht_10_13_port, 
      bht_10_12_port, bht_10_11_port, bht_10_10_port, bht_10_9_port, 
      bht_10_8_port, bht_10_7_port, bht_10_6_port, bht_10_5_port, bht_10_4_port
      , bht_10_3_port, bht_10_2_port, bht_10_1_port, bht_10_0_port, 
      bht_11_26_port, bht_11_25_port, bht_11_24_port, bht_11_23_port, 
      bht_11_22_port, bht_11_21_port, bht_11_20_port, bht_11_19_port, 
      bht_11_18_port, bht_11_17_port, bht_11_16_port, bht_11_15_port, 
      bht_11_14_port, bht_11_13_port, bht_11_12_port, bht_11_11_port, 
      bht_11_10_port, bht_11_9_port, bht_11_8_port, bht_11_7_port, 
      bht_11_6_port, bht_11_5_port, bht_11_4_port, bht_11_3_port, bht_11_2_port
      , bht_11_1_port, bht_11_0_port, bht_12_26_port, bht_12_25_port, 
      bht_12_24_port, bht_12_23_port, bht_12_22_port, bht_12_21_port, 
      bht_12_20_port, bht_12_19_port, bht_12_18_port, bht_12_17_port, 
      bht_12_16_port, bht_12_15_port, bht_12_14_port, bht_12_13_port, 
      bht_12_12_port, bht_12_11_port, bht_12_10_port, bht_12_9_port, 
      bht_12_8_port, bht_12_7_port, bht_12_6_port, bht_12_5_port, bht_12_4_port
      , bht_12_3_port, bht_12_2_port, bht_12_1_port, bht_12_0_port, 
      bht_13_26_port, bht_13_25_port, bht_13_24_port, bht_13_23_port, 
      bht_13_22_port, bht_13_21_port, bht_13_20_port, bht_13_19_port, 
      bht_13_18_port, bht_13_17_port, bht_13_16_port, bht_13_15_port, 
      bht_13_14_port, bht_13_13_port, bht_13_12_port, bht_13_11_port, 
      bht_13_10_port, bht_13_9_port, bht_13_8_port, bht_13_7_port, 
      bht_13_6_port, bht_13_5_port, bht_13_4_port, bht_13_3_port, bht_13_2_port
      , bht_13_1_port, bht_13_0_port, bht_14_26_port, bht_14_25_port, 
      bht_14_24_port, bht_14_23_port, bht_14_22_port, bht_14_21_port, 
      bht_14_20_port, bht_14_19_port, bht_14_18_port, bht_14_17_port, 
      bht_14_16_port, bht_14_15_port, bht_14_14_port, bht_14_13_port, 
      bht_14_12_port, bht_14_11_port, bht_14_10_port, bht_14_9_port, 
      bht_14_8_port, bht_14_7_port, bht_14_6_port, bht_14_5_port, bht_14_4_port
      , bht_14_3_port, bht_14_2_port, bht_14_1_port, bht_14_0_port, 
      bht_15_26_port, bht_15_25_port, bht_15_24_port, bht_15_23_port, 
      bht_15_22_port, bht_15_21_port, bht_15_20_port, bht_15_19_port, 
      bht_15_18_port, bht_15_17_port, bht_15_16_port, bht_15_15_port, 
      bht_15_14_port, bht_15_13_port, bht_15_12_port, bht_15_11_port, 
      bht_15_10_port, bht_15_9_port, bht_15_8_port, bht_15_7_port, 
      bht_15_6_port, bht_15_5_port, bht_15_4_port, bht_15_3_port, bht_15_2_port
      , bht_15_1_port, bht_15_0_port, bht_16_26_port, bht_16_25_port, 
      bht_16_24_port, bht_16_23_port, bht_16_22_port, bht_16_21_port, 
      bht_16_20_port, bht_16_19_port, bht_16_18_port, bht_16_17_port, 
      bht_16_16_port, bht_16_15_port, bht_16_14_port, bht_16_13_port, 
      bht_16_12_port, bht_16_11_port, bht_16_10_port, bht_16_9_port, 
      bht_16_8_port, bht_16_7_port, bht_16_6_port, bht_16_5_port, bht_16_4_port
      , bht_16_3_port, bht_16_2_port, bht_16_1_port, bht_16_0_port, 
      bht_17_26_port, bht_17_25_port, bht_17_24_port, bht_17_23_port, 
      bht_17_22_port, bht_17_21_port, bht_17_20_port, bht_17_19_port, 
      bht_17_18_port, bht_17_17_port, bht_17_16_port, bht_17_15_port, 
      bht_17_14_port, bht_17_13_port, bht_17_12_port, bht_17_11_port, 
      bht_17_10_port, bht_17_9_port, bht_17_8_port, bht_17_7_port, 
      bht_17_6_port, bht_17_5_port, bht_17_4_port, bht_17_3_port, bht_17_2_port
      , bht_17_1_port, bht_17_0_port, bht_18_26_port, bht_18_25_port, 
      bht_18_24_port, bht_18_23_port, bht_18_22_port, bht_18_21_port, 
      bht_18_20_port, bht_18_19_port, bht_18_18_port, bht_18_17_port, 
      bht_18_16_port, bht_18_15_port, bht_18_14_port, bht_18_13_port, 
      bht_18_12_port, bht_18_11_port, bht_18_10_port, bht_18_9_port, 
      bht_18_8_port, bht_18_7_port, bht_18_6_port, bht_18_5_port, bht_18_4_port
      , bht_18_3_port, bht_18_2_port, bht_18_1_port, bht_18_0_port, 
      bht_19_26_port, bht_19_25_port, bht_19_24_port, bht_19_23_port, 
      bht_19_22_port, bht_19_21_port, bht_19_20_port, bht_19_19_port, 
      bht_19_18_port, bht_19_17_port, bht_19_16_port, bht_19_15_port, 
      bht_19_14_port, bht_19_13_port, bht_19_12_port, bht_19_11_port, 
      bht_19_10_port, bht_19_9_port, bht_19_8_port, bht_19_7_port, 
      bht_19_6_port, bht_19_5_port, bht_19_4_port, bht_19_3_port, bht_19_2_port
      , bht_19_1_port, bht_19_0_port, bht_20_26_port, bht_20_25_port, 
      bht_20_24_port, bht_20_23_port, bht_20_22_port, bht_20_21_port, 
      bht_20_20_port, bht_20_19_port, bht_20_18_port, bht_20_17_port, 
      bht_20_16_port, bht_20_15_port, bht_20_14_port, bht_20_13_port, 
      bht_20_12_port, bht_20_11_port, bht_20_10_port, bht_20_9_port, 
      bht_20_8_port, bht_20_7_port, bht_20_6_port, bht_20_5_port, bht_20_4_port
      , bht_20_3_port, bht_20_2_port, bht_20_1_port, bht_20_0_port, 
      bht_21_26_port, bht_21_25_port, bht_21_24_port, bht_21_23_port, 
      bht_21_22_port, bht_21_21_port, bht_21_20_port, bht_21_19_port, 
      bht_21_18_port, bht_21_17_port, bht_21_16_port, bht_21_15_port, 
      bht_21_14_port, bht_21_13_port, bht_21_12_port, bht_21_11_port, 
      bht_21_10_port, bht_21_9_port, bht_21_8_port, bht_21_7_port, 
      bht_21_6_port, bht_21_5_port, bht_21_4_port, bht_21_3_port, bht_21_2_port
      , bht_21_1_port, bht_21_0_port, bht_22_26_port, bht_22_25_port, 
      bht_22_24_port, bht_22_23_port, bht_22_22_port, bht_22_21_port, 
      bht_22_20_port, bht_22_19_port, bht_22_18_port, bht_22_17_port, 
      bht_22_16_port, bht_22_15_port, bht_22_14_port, bht_22_13_port, 
      bht_22_12_port, bht_22_11_port, bht_22_10_port, bht_22_9_port, 
      bht_22_8_port, bht_22_7_port, bht_22_6_port, bht_22_5_port, bht_22_4_port
      , bht_22_3_port, bht_22_2_port, bht_22_1_port, bht_22_0_port, 
      bht_23_26_port, bht_23_25_port, bht_23_24_port, bht_23_23_port, 
      bht_23_22_port, bht_23_21_port, bht_23_20_port, bht_23_19_port, 
      bht_23_18_port, bht_23_17_port, bht_23_16_port, bht_23_15_port, 
      bht_23_14_port, bht_23_13_port, bht_23_12_port, bht_23_11_port, 
      bht_23_10_port, bht_23_9_port, bht_23_8_port, bht_23_7_port, 
      bht_23_6_port, bht_23_5_port, bht_23_4_port, bht_23_3_port, bht_23_2_port
      , bht_23_1_port, bht_23_0_port, bht_24_26_port, bht_24_25_port, 
      bht_24_24_port, bht_24_23_port, bht_24_22_port, bht_24_21_port, 
      bht_24_20_port, bht_24_19_port, bht_24_18_port, bht_24_17_port, 
      bht_24_16_port, bht_24_15_port, bht_24_14_port, bht_24_13_port, 
      bht_24_12_port, bht_24_11_port, bht_24_10_port, bht_24_9_port, 
      bht_24_8_port, bht_24_7_port, bht_24_6_port, bht_24_5_port, bht_24_4_port
      , bht_24_3_port, bht_24_2_port, bht_24_1_port, bht_24_0_port, 
      bht_25_26_port, bht_25_25_port, bht_25_24_port, bht_25_23_port, 
      bht_25_22_port, bht_25_21_port, bht_25_20_port, bht_25_19_port, 
      bht_25_18_port, bht_25_17_port, bht_25_16_port, bht_25_15_port, 
      bht_25_14_port, bht_25_13_port, bht_25_12_port, bht_25_11_port, 
      bht_25_10_port, bht_25_9_port, bht_25_8_port, bht_25_7_port, 
      bht_25_6_port, bht_25_5_port, bht_25_4_port, bht_25_3_port, bht_25_2_port
      , bht_25_1_port, bht_25_0_port, bht_26_26_port, bht_26_25_port, 
      bht_26_24_port, bht_26_23_port, bht_26_22_port, bht_26_21_port, 
      bht_26_20_port, bht_26_19_port, bht_26_18_port, bht_26_17_port, 
      bht_26_16_port, bht_26_15_port, bht_26_14_port, bht_26_13_port, 
      bht_26_12_port, bht_26_11_port, bht_26_10_port, bht_26_9_port, 
      bht_26_8_port, bht_26_7_port, bht_26_6_port, bht_26_5_port, bht_26_4_port
      , bht_26_3_port, bht_26_2_port, bht_26_1_port, bht_26_0_port, 
      bht_27_26_port, bht_27_25_port, bht_27_24_port, bht_27_23_port, 
      bht_27_22_port, bht_27_21_port, bht_27_20_port, bht_27_19_port, 
      bht_27_18_port, bht_27_17_port, bht_27_16_port, bht_27_15_port, 
      bht_27_14_port, bht_27_13_port, bht_27_12_port, bht_27_11_port, 
      bht_27_10_port, bht_27_9_port, bht_27_8_port, bht_27_7_port, 
      bht_27_6_port, bht_27_5_port, bht_27_4_port, bht_27_3_port, bht_27_2_port
      , bht_27_1_port, bht_27_0_port, bht_28_26_port, bht_28_25_port, 
      bht_28_24_port, bht_28_23_port, bht_28_22_port, bht_28_21_port, 
      bht_28_20_port, bht_28_19_port, bht_28_18_port, bht_28_17_port, 
      bht_28_16_port, bht_28_15_port, bht_28_14_port, bht_28_13_port, 
      bht_28_12_port, bht_28_11_port, bht_28_10_port, bht_28_9_port, 
      bht_28_8_port, bht_28_7_port, bht_28_6_port, bht_28_5_port, bht_28_4_port
      , bht_28_3_port, bht_28_2_port, bht_28_1_port, bht_28_0_port, 
      bht_29_26_port, bht_29_25_port, bht_29_24_port, bht_29_23_port, 
      bht_29_22_port, bht_29_21_port, bht_29_20_port, bht_29_19_port, 
      bht_29_18_port, bht_29_17_port, bht_29_16_port, bht_29_15_port, 
      bht_29_14_port, bht_29_13_port, bht_29_12_port, bht_29_11_port, 
      bht_29_10_port, bht_29_9_port, bht_29_8_port, bht_29_7_port, 
      bht_29_6_port, bht_29_5_port, bht_29_4_port, bht_29_3_port, bht_29_2_port
      , bht_29_1_port, bht_29_0_port, bht_30_26_port, bht_30_25_port, 
      bht_30_24_port, bht_30_23_port, bht_30_22_port, bht_30_21_port, 
      bht_30_20_port, bht_30_19_port, bht_30_18_port, bht_30_17_port, 
      bht_30_16_port, bht_30_15_port, bht_30_14_port, bht_30_13_port, 
      bht_30_12_port, bht_30_11_port, bht_30_10_port, bht_30_9_port, 
      bht_30_8_port, bht_30_7_port, bht_30_6_port, bht_30_5_port, bht_30_4_port
      , bht_30_3_port, bht_30_2_port, bht_30_1_port, bht_30_0_port, 
      bht_31_26_port, bht_31_25_port, bht_31_24_port, bht_31_23_port, 
      bht_31_22_port, bht_31_21_port, bht_31_20_port, bht_31_19_port, 
      bht_31_18_port, bht_31_17_port, bht_31_16_port, bht_31_15_port, 
      bht_31_14_port, bht_31_13_port, bht_31_12_port, bht_31_11_port, 
      bht_31_10_port, bht_31_9_port, bht_31_8_port, bht_31_7_port, 
      bht_31_6_port, bht_31_5_port, bht_31_4_port, bht_31_3_port, bht_31_2_port
      , bht_31_1_port, bht_31_0_port, N125, N126, N127, N128, N129, N130, N131,
      N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, 
      N144, N145, N146, N147, N148, N149, N150, N151, index_r_4_port, 
      index_r_3_port, index_r_2_port, index_r_1_port, index_r_0_port, 
      entry_r_26_port, entry_r_25_port, entry_r_24_port, entry_r_23_port, 
      entry_r_22_port, entry_r_21_port, entry_r_20_port, entry_r_19_port, 
      entry_r_18_port, entry_r_17_port, entry_r_16_port, entry_r_15_port, 
      entry_r_14_port, entry_r_13_port, entry_r_12_port, entry_r_11_port, 
      entry_r_10_port, entry_r_9_port, entry_r_8_port, entry_r_7_port, 
      entry_r_6_port, entry_r_5_port, entry_r_4_port, entry_r_3_port, 
      entry_r_2_port, entry_r_1_port, entry_r_0_port, N188, sig_bal_delay, 
      opcd_delay_5_port, opcd_delay_4_port, opcd_delay_3_port, 
      opcd_delay_2_port, sig_brt_delay, N2110, N2164, N2218, N2272, N2326, 
      N2380, N2434, N2488, N2542, N2596, N2650, N2704, N2758, N2812, N2866, 
      N2920, N2974, N3028, N3082, N3136, N3190, N3244, N3298, N3352, N3406, 
      N3460, N3514, N3568, N3622, N3676, N3730, N3733, N3735, N3737, N3739, 
      N3741, N3743, N3745, N3747, N3749, N3751, N3753, N3755, N3757, N3759, 
      N3761, N3763, N3765, N3767, N3769, N3771, N3773, N3775, N3777, N3779, 
      N3781, N3783, N3784, N3785, n187, n200, n202, n207, n214, n219, n1, n2, 
      n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, 
      n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33
      , n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, 
      n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62
      , n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, 
      n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91
      , n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, 
      n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, 
      n117, n118, n119, n120, n121, n122, n123, n124, n125_port, n126_port, 
      n127_port, n128_port, n129_port, n130_port, n131_port, n132_port, 
      n133_port, n134_port, n135_port, n136_port, n137_port, n138_port, 
      n139_port, n140_port, n141_port, n142_port, n143_port, n144_port, 
      n145_port, n146_port, n147_port, n148_port, n149_port, n150_port, 
      n151_port, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n188_port, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n201, n203, n204, n205, n206, n208, n209, n210, n211, n212, 
      n213, n215, n216, n217, n218, n220, n221, n222, n223, n224, n225, n226, 
      n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, 
      n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, 
      n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, 
      n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, 
      n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, 
      n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, 
      n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, 
      n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, 
      n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, 
      n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, 
      n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, 
      n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, 
      n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, 
      n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, 
      n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, 
      n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, 
      n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, 
      n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, 
      n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, 
      n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, 
      n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, 
      n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, 
      n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, 
      n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, 
      n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, 
      n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, 
      n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, 
      n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, 
      n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, 
      n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, 
      n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, 
      n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, 
      n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, 
      n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, 
      n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, 
      n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, 
      n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, 
      n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, 
      n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, 
      n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, 
      n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, 
      n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, 
      n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742, 
      n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, 
      n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, 
      n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, 
      n779, n780, n781, n782, n783, n784, n785, net108064, net108065, net108066
      , net108067, net108068, net108069, net108070, net108071, net108072, 
      net108073, net108074, net108075, net108076, net108077, net108078, 
      net108079, net108080, net108081, net108082, net108083, net108084, 
      net108085, net108086, net108087, net108088, net108089, net108090, 
      net108091, net108092, net108093, net108094, net108095, net108096 : 
      std_logic;

begin
   sig_brt <= sig_brt_tmp;
   
   index_r_reg_4_inst : DLH_X1 port map( G => N188, D => addr(6), Q => 
                           index_r_4_port);
   index_r_reg_3_inst : DLH_X1 port map( G => N188, D => addr(5), Q => 
                           index_r_3_port);
   index_r_reg_2_inst : DLH_X1 port map( G => N188, D => addr(4), Q => 
                           index_r_2_port);
   index_r_reg_1_inst : DLH_X1 port map( G => N188, D => addr(3), Q => 
                           index_r_1_port);
   index_r_reg_0_inst : DLH_X1 port map( G => N188, D => addr(2), Q => 
                           index_r_0_port);
   sig_bal_delay_reg : DFFR_X1 port map( D => sig_bal, CK => clk, RN => rst, Q 
                           => sig_bal_delay, QN => n6);
   opcd_delay_reg_5_inst : DFFR_X1 port map( D => opcd(5), CK => clk, RN => rst
                           , Q => opcd_delay_5_port, QN => net108096);
   opcd_delay_reg_4_inst : DFFR_X1 port map( D => opcd(4), CK => clk, RN => rst
                           , Q => opcd_delay_4_port, QN => net108095);
   opcd_delay_reg_3_inst : DFFR_X1 port map( D => opcd(3), CK => clk, RN => rst
                           , Q => opcd_delay_3_port, QN => net108094);
   opcd_delay_reg_2_inst : DFFR_X1 port map( D => opcd(2), CK => clk, RN => rst
                           , Q => opcd_delay_2_port, QN => net108093);
   opcd_delay_reg_1_inst : DFFR_X1 port map( D => opcd(1), CK => clk, RN => rst
                           , Q => net108092, QN => n214);
   opcd_delay_reg_0_inst : DFFR_X1 port map( D => opcd(0), CK => clk, RN => rst
                           , Q => net108091, QN => n219);
   index_r_delay_reg_4_inst : DFFR_X1 port map( D => index_r_4_port, CK => clk,
                           RN => rst, Q => n4, QN => n35);
   index_r_delay_reg_3_inst : DFFR_X1 port map( D => index_r_3_port, CK => clk,
                           RN => rst, Q => n8, QN => n187);
   index_r_delay_reg_2_inst : DFFR_X1 port map( D => index_r_2_port, CK => clk,
                           RN => rst, Q => n1, QN => n34);
   index_r_delay_reg_1_inst : DFFR_X1 port map( D => index_r_1_port, CK => clk,
                           RN => rst, Q => n5, QN => n202);
   index_r_delay_reg_0_inst : DFFR_X1 port map( D => index_r_0_port, CK => clk,
                           RN => rst, Q => n2, QN => n200);
   bht_reg_31_25_inst : DLH_X1 port map( G => N2110, D => N3783, Q => 
                           bht_31_25_port);
   entry_r_reg_26_inst : DLH_X1 port map( G => N188, D => N151, Q => 
                           entry_r_26_port);
   entry_r_delay_reg_26_inst : DFFR_X1 port map( D => entry_r_26_port, CK => 
                           clk, RN => rst, Q => net108090, QN => n33);
   bht_reg_0_26_inst : DLH_X1 port map( G => N3784, D => N3785, Q => 
                           bht_0_26_port);
   bht_reg_2_26_inst : DLH_X1 port map( G => N3676, D => N3785, Q => 
                           bht_2_26_port);
   bht_reg_4_26_inst : DLH_X1 port map( G => N3568, D => N3785, Q => 
                           bht_4_26_port);
   bht_reg_6_26_inst : DLH_X1 port map( G => N3460, D => N3785, Q => 
                           bht_6_26_port);
   bht_reg_8_26_inst : DLH_X1 port map( G => N3352, D => N3785, Q => 
                           bht_8_26_port);
   bht_reg_10_26_inst : DLH_X1 port map( G => N3244, D => N3785, Q => 
                           bht_10_26_port);
   bht_reg_12_26_inst : DLH_X1 port map( G => N3136, D => N3785, Q => 
                           bht_12_26_port);
   bht_reg_14_26_inst : DLH_X1 port map( G => N3028, D => N3785, Q => 
                           bht_14_26_port);
   bht_reg_16_26_inst : DLH_X1 port map( G => N2920, D => N3785, Q => 
                           bht_16_26_port);
   bht_reg_18_26_inst : DLH_X1 port map( G => N2812, D => N3785, Q => 
                           bht_18_26_port);
   bht_reg_20_26_inst : DLH_X1 port map( G => N2704, D => N3785, Q => 
                           bht_20_26_port);
   bht_reg_22_26_inst : DLH_X1 port map( G => N2596, D => N3785, Q => 
                           bht_22_26_port);
   bht_reg_24_26_inst : DLH_X1 port map( G => N2488, D => N3785, Q => 
                           bht_24_26_port);
   bht_reg_26_26_inst : DLH_X1 port map( G => N2380, D => N3785, Q => 
                           bht_26_26_port);
   bht_reg_28_26_inst : DLH_X1 port map( G => N2272, D => N3785, Q => 
                           bht_28_26_port);
   bht_reg_30_26_inst : DLH_X1 port map( G => N2164, D => N3785, Q => 
                           bht_30_26_port);
   bht_reg_31_26_inst : DLH_X1 port map( G => N2110, D => N3785, Q => 
                           bht_31_26_port);
   bht_reg_29_26_inst : DLH_X1 port map( G => N2218, D => N3785, Q => 
                           bht_29_26_port);
   bht_reg_27_26_inst : DLH_X1 port map( G => N2326, D => N3785, Q => 
                           bht_27_26_port);
   bht_reg_25_26_inst : DLH_X1 port map( G => N2434, D => N3785, Q => 
                           bht_25_26_port);
   bht_reg_23_26_inst : DLH_X1 port map( G => N2542, D => N3785, Q => 
                           bht_23_26_port);
   bht_reg_21_26_inst : DLH_X1 port map( G => N2650, D => N3785, Q => 
                           bht_21_26_port);
   bht_reg_19_26_inst : DLH_X1 port map( G => N2758, D => N3785, Q => 
                           bht_19_26_port);
   bht_reg_17_26_inst : DLH_X1 port map( G => N2866, D => N3785, Q => 
                           bht_17_26_port);
   bht_reg_15_26_inst : DLH_X1 port map( G => N2974, D => N3785, Q => 
                           bht_15_26_port);
   bht_reg_13_26_inst : DLH_X1 port map( G => N3082, D => N3785, Q => 
                           bht_13_26_port);
   bht_reg_11_26_inst : DLH_X1 port map( G => N3190, D => N3785, Q => 
                           bht_11_26_port);
   bht_reg_9_26_inst : DLH_X1 port map( G => N3298, D => N3785, Q => 
                           bht_9_26_port);
   bht_reg_7_26_inst : DLH_X1 port map( G => N3406, D => N3785, Q => 
                           bht_7_26_port);
   bht_reg_5_26_inst : DLH_X1 port map( G => N3514, D => N3785, Q => 
                           bht_5_26_port);
   bht_reg_3_26_inst : DLH_X1 port map( G => N3622, D => N3785, Q => 
                           bht_3_26_port);
   bht_reg_1_26_inst : DLH_X1 port map( G => N3730, D => N3785, Q => 
                           bht_1_26_port);
   entry_r_reg_24_inst : DLH_X1 port map( G => N188, D => N149, Q => 
                           entry_r_24_port);
   entry_r_delay_reg_24_inst : DFFR_X1 port map( D => entry_r_24_port, CK => 
                           clk, RN => rst, Q => net108089, QN => n32);
   bht_reg_0_24_inst : DLH_X1 port map( G => N3784, D => N3781, Q => 
                           bht_0_24_port);
   bht_reg_2_24_inst : DLH_X1 port map( G => N3676, D => N3781, Q => 
                           bht_2_24_port);
   bht_reg_4_24_inst : DLH_X1 port map( G => N3568, D => N3781, Q => 
                           bht_4_24_port);
   bht_reg_6_24_inst : DLH_X1 port map( G => N3460, D => N3781, Q => 
                           bht_6_24_port);
   bht_reg_8_24_inst : DLH_X1 port map( G => N3352, D => N3781, Q => 
                           bht_8_24_port);
   bht_reg_10_24_inst : DLH_X1 port map( G => N3244, D => N3781, Q => 
                           bht_10_24_port);
   bht_reg_12_24_inst : DLH_X1 port map( G => N3136, D => N3781, Q => 
                           bht_12_24_port);
   bht_reg_14_24_inst : DLH_X1 port map( G => N3028, D => N3781, Q => 
                           bht_14_24_port);
   bht_reg_16_24_inst : DLH_X1 port map( G => N2920, D => N3781, Q => 
                           bht_16_24_port);
   bht_reg_18_24_inst : DLH_X1 port map( G => N2812, D => N3781, Q => 
                           bht_18_24_port);
   bht_reg_20_24_inst : DLH_X1 port map( G => N2704, D => N3781, Q => 
                           bht_20_24_port);
   bht_reg_22_24_inst : DLH_X1 port map( G => N2596, D => N3781, Q => 
                           bht_22_24_port);
   bht_reg_24_24_inst : DLH_X1 port map( G => N2488, D => N3781, Q => 
                           bht_24_24_port);
   bht_reg_26_24_inst : DLH_X1 port map( G => N2380, D => N3781, Q => 
                           bht_26_24_port);
   bht_reg_28_24_inst : DLH_X1 port map( G => N2272, D => N3781, Q => 
                           bht_28_24_port);
   bht_reg_30_24_inst : DLH_X1 port map( G => N2164, D => N3781, Q => 
                           bht_30_24_port);
   bht_reg_31_24_inst : DLH_X1 port map( G => N2110, D => N3781, Q => 
                           bht_31_24_port);
   bht_reg_29_24_inst : DLH_X1 port map( G => N2218, D => N3781, Q => 
                           bht_29_24_port);
   bht_reg_27_24_inst : DLH_X1 port map( G => N2326, D => N3781, Q => 
                           bht_27_24_port);
   bht_reg_25_24_inst : DLH_X1 port map( G => N2434, D => N3781, Q => 
                           bht_25_24_port);
   bht_reg_23_24_inst : DLH_X1 port map( G => N2542, D => N3781, Q => 
                           bht_23_24_port);
   bht_reg_21_24_inst : DLH_X1 port map( G => N2650, D => N3781, Q => 
                           bht_21_24_port);
   bht_reg_19_24_inst : DLH_X1 port map( G => N2758, D => N3781, Q => 
                           bht_19_24_port);
   bht_reg_17_24_inst : DLH_X1 port map( G => N2866, D => N3781, Q => 
                           bht_17_24_port);
   bht_reg_15_24_inst : DLH_X1 port map( G => N2974, D => N3781, Q => 
                           bht_15_24_port);
   bht_reg_13_24_inst : DLH_X1 port map( G => N3082, D => N3781, Q => 
                           bht_13_24_port);
   bht_reg_11_24_inst : DLH_X1 port map( G => N3190, D => N3781, Q => 
                           bht_11_24_port);
   bht_reg_9_24_inst : DLH_X1 port map( G => N3298, D => N3781, Q => 
                           bht_9_24_port);
   bht_reg_7_24_inst : DLH_X1 port map( G => N3406, D => N3781, Q => 
                           bht_7_24_port);
   bht_reg_5_24_inst : DLH_X1 port map( G => N3514, D => N3781, Q => 
                           bht_5_24_port);
   bht_reg_3_24_inst : DLH_X1 port map( G => N3622, D => N3781, Q => 
                           bht_3_24_port);
   bht_reg_1_24_inst : DLH_X1 port map( G => N3730, D => N3781, Q => 
                           bht_1_24_port);
   entry_r_reg_23_inst : DLH_X1 port map( G => N188, D => N148, Q => 
                           entry_r_23_port);
   entry_r_delay_reg_23_inst : DFFR_X1 port map( D => entry_r_23_port, CK => 
                           clk, RN => rst, Q => net108088, QN => n31);
   bht_reg_0_23_inst : DLH_X1 port map( G => N3784, D => N3779, Q => 
                           bht_0_23_port);
   bht_reg_2_23_inst : DLH_X1 port map( G => N3676, D => N3779, Q => 
                           bht_2_23_port);
   bht_reg_4_23_inst : DLH_X1 port map( G => N3568, D => N3779, Q => 
                           bht_4_23_port);
   bht_reg_6_23_inst : DLH_X1 port map( G => N3460, D => N3779, Q => 
                           bht_6_23_port);
   bht_reg_8_23_inst : DLH_X1 port map( G => N3352, D => N3779, Q => 
                           bht_8_23_port);
   bht_reg_10_23_inst : DLH_X1 port map( G => N3244, D => N3779, Q => 
                           bht_10_23_port);
   bht_reg_12_23_inst : DLH_X1 port map( G => N3136, D => N3779, Q => 
                           bht_12_23_port);
   bht_reg_14_23_inst : DLH_X1 port map( G => N3028, D => N3779, Q => 
                           bht_14_23_port);
   bht_reg_16_23_inst : DLH_X1 port map( G => N2920, D => N3779, Q => 
                           bht_16_23_port);
   bht_reg_18_23_inst : DLH_X1 port map( G => N2812, D => N3779, Q => 
                           bht_18_23_port);
   bht_reg_20_23_inst : DLH_X1 port map( G => N2704, D => N3779, Q => 
                           bht_20_23_port);
   bht_reg_22_23_inst : DLH_X1 port map( G => N2596, D => N3779, Q => 
                           bht_22_23_port);
   bht_reg_24_23_inst : DLH_X1 port map( G => N2488, D => N3779, Q => 
                           bht_24_23_port);
   bht_reg_26_23_inst : DLH_X1 port map( G => N2380, D => N3779, Q => 
                           bht_26_23_port);
   bht_reg_28_23_inst : DLH_X1 port map( G => N2272, D => N3779, Q => 
                           bht_28_23_port);
   bht_reg_30_23_inst : DLH_X1 port map( G => N2164, D => N3779, Q => 
                           bht_30_23_port);
   bht_reg_31_23_inst : DLH_X1 port map( G => N2110, D => N3779, Q => 
                           bht_31_23_port);
   bht_reg_29_23_inst : DLH_X1 port map( G => N2218, D => N3779, Q => 
                           bht_29_23_port);
   bht_reg_27_23_inst : DLH_X1 port map( G => N2326, D => N3779, Q => 
                           bht_27_23_port);
   bht_reg_25_23_inst : DLH_X1 port map( G => N2434, D => N3779, Q => 
                           bht_25_23_port);
   bht_reg_23_23_inst : DLH_X1 port map( G => N2542, D => N3779, Q => 
                           bht_23_23_port);
   bht_reg_21_23_inst : DLH_X1 port map( G => N2650, D => N3779, Q => 
                           bht_21_23_port);
   bht_reg_19_23_inst : DLH_X1 port map( G => N2758, D => N3779, Q => 
                           bht_19_23_port);
   bht_reg_17_23_inst : DLH_X1 port map( G => N2866, D => N3779, Q => 
                           bht_17_23_port);
   bht_reg_15_23_inst : DLH_X1 port map( G => N2974, D => N3779, Q => 
                           bht_15_23_port);
   bht_reg_13_23_inst : DLH_X1 port map( G => N3082, D => N3779, Q => 
                           bht_13_23_port);
   bht_reg_11_23_inst : DLH_X1 port map( G => N3190, D => N3779, Q => 
                           bht_11_23_port);
   bht_reg_9_23_inst : DLH_X1 port map( G => N3298, D => N3779, Q => 
                           bht_9_23_port);
   bht_reg_7_23_inst : DLH_X1 port map( G => N3406, D => N3779, Q => 
                           bht_7_23_port);
   bht_reg_5_23_inst : DLH_X1 port map( G => N3514, D => N3779, Q => 
                           bht_5_23_port);
   bht_reg_3_23_inst : DLH_X1 port map( G => N3622, D => N3779, Q => 
                           bht_3_23_port);
   bht_reg_1_23_inst : DLH_X1 port map( G => N3730, D => N3779, Q => 
                           bht_1_23_port);
   entry_r_reg_22_inst : DLH_X1 port map( G => N188, D => N147, Q => 
                           entry_r_22_port);
   entry_r_delay_reg_22_inst : DFFR_X1 port map( D => entry_r_22_port, CK => 
                           clk, RN => rst, Q => net108087, QN => n30);
   bht_reg_0_22_inst : DLH_X1 port map( G => N3784, D => N3777, Q => 
                           bht_0_22_port);
   bht_reg_2_22_inst : DLH_X1 port map( G => N3676, D => N3777, Q => 
                           bht_2_22_port);
   bht_reg_4_22_inst : DLH_X1 port map( G => N3568, D => N3777, Q => 
                           bht_4_22_port);
   bht_reg_6_22_inst : DLH_X1 port map( G => N3460, D => N3777, Q => 
                           bht_6_22_port);
   bht_reg_8_22_inst : DLH_X1 port map( G => N3352, D => N3777, Q => 
                           bht_8_22_port);
   bht_reg_10_22_inst : DLH_X1 port map( G => N3244, D => N3777, Q => 
                           bht_10_22_port);
   bht_reg_12_22_inst : DLH_X1 port map( G => N3136, D => N3777, Q => 
                           bht_12_22_port);
   bht_reg_14_22_inst : DLH_X1 port map( G => N3028, D => N3777, Q => 
                           bht_14_22_port);
   bht_reg_16_22_inst : DLH_X1 port map( G => N2920, D => N3777, Q => 
                           bht_16_22_port);
   bht_reg_18_22_inst : DLH_X1 port map( G => N2812, D => N3777, Q => 
                           bht_18_22_port);
   bht_reg_20_22_inst : DLH_X1 port map( G => N2704, D => N3777, Q => 
                           bht_20_22_port);
   bht_reg_22_22_inst : DLH_X1 port map( G => N2596, D => N3777, Q => 
                           bht_22_22_port);
   bht_reg_24_22_inst : DLH_X1 port map( G => N2488, D => N3777, Q => 
                           bht_24_22_port);
   bht_reg_26_22_inst : DLH_X1 port map( G => N2380, D => N3777, Q => 
                           bht_26_22_port);
   bht_reg_28_22_inst : DLH_X1 port map( G => N2272, D => N3777, Q => 
                           bht_28_22_port);
   bht_reg_30_22_inst : DLH_X1 port map( G => N2164, D => N3777, Q => 
                           bht_30_22_port);
   bht_reg_31_22_inst : DLH_X1 port map( G => N2110, D => N3777, Q => 
                           bht_31_22_port);
   bht_reg_29_22_inst : DLH_X1 port map( G => N2218, D => N3777, Q => 
                           bht_29_22_port);
   bht_reg_27_22_inst : DLH_X1 port map( G => N2326, D => N3777, Q => 
                           bht_27_22_port);
   bht_reg_25_22_inst : DLH_X1 port map( G => N2434, D => N3777, Q => 
                           bht_25_22_port);
   bht_reg_23_22_inst : DLH_X1 port map( G => N2542, D => N3777, Q => 
                           bht_23_22_port);
   bht_reg_21_22_inst : DLH_X1 port map( G => N2650, D => N3777, Q => 
                           bht_21_22_port);
   bht_reg_19_22_inst : DLH_X1 port map( G => N2758, D => N3777, Q => 
                           bht_19_22_port);
   bht_reg_17_22_inst : DLH_X1 port map( G => N2866, D => N3777, Q => 
                           bht_17_22_port);
   bht_reg_15_22_inst : DLH_X1 port map( G => N2974, D => N3777, Q => 
                           bht_15_22_port);
   bht_reg_13_22_inst : DLH_X1 port map( G => N3082, D => N3777, Q => 
                           bht_13_22_port);
   bht_reg_11_22_inst : DLH_X1 port map( G => N3190, D => N3777, Q => 
                           bht_11_22_port);
   bht_reg_9_22_inst : DLH_X1 port map( G => N3298, D => N3777, Q => 
                           bht_9_22_port);
   bht_reg_7_22_inst : DLH_X1 port map( G => N3406, D => N3777, Q => 
                           bht_7_22_port);
   bht_reg_5_22_inst : DLH_X1 port map( G => N3514, D => N3777, Q => 
                           bht_5_22_port);
   bht_reg_3_22_inst : DLH_X1 port map( G => N3622, D => N3777, Q => 
                           bht_3_22_port);
   bht_reg_1_22_inst : DLH_X1 port map( G => N3730, D => N3777, Q => 
                           bht_1_22_port);
   entry_r_reg_21_inst : DLH_X1 port map( G => N188, D => N146, Q => 
                           entry_r_21_port);
   entry_r_delay_reg_21_inst : DFFR_X1 port map( D => entry_r_21_port, CK => 
                           clk, RN => rst, Q => net108086, QN => n29);
   bht_reg_0_21_inst : DLH_X1 port map( G => N3784, D => N3775, Q => 
                           bht_0_21_port);
   bht_reg_2_21_inst : DLH_X1 port map( G => N3676, D => N3775, Q => 
                           bht_2_21_port);
   bht_reg_4_21_inst : DLH_X1 port map( G => N3568, D => N3775, Q => 
                           bht_4_21_port);
   bht_reg_6_21_inst : DLH_X1 port map( G => N3460, D => N3775, Q => 
                           bht_6_21_port);
   bht_reg_8_21_inst : DLH_X1 port map( G => N3352, D => N3775, Q => 
                           bht_8_21_port);
   bht_reg_10_21_inst : DLH_X1 port map( G => N3244, D => N3775, Q => 
                           bht_10_21_port);
   bht_reg_12_21_inst : DLH_X1 port map( G => N3136, D => N3775, Q => 
                           bht_12_21_port);
   bht_reg_14_21_inst : DLH_X1 port map( G => N3028, D => N3775, Q => 
                           bht_14_21_port);
   bht_reg_16_21_inst : DLH_X1 port map( G => N2920, D => N3775, Q => 
                           bht_16_21_port);
   bht_reg_18_21_inst : DLH_X1 port map( G => N2812, D => N3775, Q => 
                           bht_18_21_port);
   bht_reg_20_21_inst : DLH_X1 port map( G => N2704, D => N3775, Q => 
                           bht_20_21_port);
   bht_reg_22_21_inst : DLH_X1 port map( G => N2596, D => N3775, Q => 
                           bht_22_21_port);
   bht_reg_24_21_inst : DLH_X1 port map( G => N2488, D => N3775, Q => 
                           bht_24_21_port);
   bht_reg_26_21_inst : DLH_X1 port map( G => N2380, D => N3775, Q => 
                           bht_26_21_port);
   bht_reg_28_21_inst : DLH_X1 port map( G => N2272, D => N3775, Q => 
                           bht_28_21_port);
   bht_reg_30_21_inst : DLH_X1 port map( G => N2164, D => N3775, Q => 
                           bht_30_21_port);
   bht_reg_31_21_inst : DLH_X1 port map( G => N2110, D => N3775, Q => 
                           bht_31_21_port);
   bht_reg_29_21_inst : DLH_X1 port map( G => N2218, D => N3775, Q => 
                           bht_29_21_port);
   bht_reg_27_21_inst : DLH_X1 port map( G => N2326, D => N3775, Q => 
                           bht_27_21_port);
   bht_reg_25_21_inst : DLH_X1 port map( G => N2434, D => N3775, Q => 
                           bht_25_21_port);
   bht_reg_23_21_inst : DLH_X1 port map( G => N2542, D => N3775, Q => 
                           bht_23_21_port);
   bht_reg_21_21_inst : DLH_X1 port map( G => N2650, D => N3775, Q => 
                           bht_21_21_port);
   bht_reg_19_21_inst : DLH_X1 port map( G => N2758, D => N3775, Q => 
                           bht_19_21_port);
   bht_reg_17_21_inst : DLH_X1 port map( G => N2866, D => N3775, Q => 
                           bht_17_21_port);
   bht_reg_15_21_inst : DLH_X1 port map( G => N2974, D => N3775, Q => 
                           bht_15_21_port);
   bht_reg_13_21_inst : DLH_X1 port map( G => N3082, D => N3775, Q => 
                           bht_13_21_port);
   bht_reg_11_21_inst : DLH_X1 port map( G => N3190, D => N3775, Q => 
                           bht_11_21_port);
   bht_reg_9_21_inst : DLH_X1 port map( G => N3298, D => N3775, Q => 
                           bht_9_21_port);
   bht_reg_7_21_inst : DLH_X1 port map( G => N3406, D => N3775, Q => 
                           bht_7_21_port);
   bht_reg_5_21_inst : DLH_X1 port map( G => N3514, D => N3775, Q => 
                           bht_5_21_port);
   bht_reg_3_21_inst : DLH_X1 port map( G => N3622, D => N3775, Q => 
                           bht_3_21_port);
   bht_reg_1_21_inst : DLH_X1 port map( G => N3730, D => N3775, Q => 
                           bht_1_21_port);
   entry_r_reg_20_inst : DLH_X1 port map( G => N188, D => N145, Q => 
                           entry_r_20_port);
   entry_r_delay_reg_20_inst : DFFR_X1 port map( D => entry_r_20_port, CK => 
                           clk, RN => rst, Q => net108085, QN => n28);
   bht_reg_0_20_inst : DLH_X1 port map( G => N3784, D => N3773, Q => 
                           bht_0_20_port);
   bht_reg_2_20_inst : DLH_X1 port map( G => N3676, D => N3773, Q => 
                           bht_2_20_port);
   bht_reg_4_20_inst : DLH_X1 port map( G => N3568, D => N3773, Q => 
                           bht_4_20_port);
   bht_reg_6_20_inst : DLH_X1 port map( G => N3460, D => N3773, Q => 
                           bht_6_20_port);
   bht_reg_8_20_inst : DLH_X1 port map( G => N3352, D => N3773, Q => 
                           bht_8_20_port);
   bht_reg_10_20_inst : DLH_X1 port map( G => N3244, D => N3773, Q => 
                           bht_10_20_port);
   bht_reg_12_20_inst : DLH_X1 port map( G => N3136, D => N3773, Q => 
                           bht_12_20_port);
   bht_reg_14_20_inst : DLH_X1 port map( G => N3028, D => N3773, Q => 
                           bht_14_20_port);
   bht_reg_16_20_inst : DLH_X1 port map( G => N2920, D => N3773, Q => 
                           bht_16_20_port);
   bht_reg_18_20_inst : DLH_X1 port map( G => N2812, D => N3773, Q => 
                           bht_18_20_port);
   bht_reg_20_20_inst : DLH_X1 port map( G => N2704, D => N3773, Q => 
                           bht_20_20_port);
   bht_reg_22_20_inst : DLH_X1 port map( G => N2596, D => N3773, Q => 
                           bht_22_20_port);
   bht_reg_24_20_inst : DLH_X1 port map( G => N2488, D => N3773, Q => 
                           bht_24_20_port);
   bht_reg_26_20_inst : DLH_X1 port map( G => N2380, D => N3773, Q => 
                           bht_26_20_port);
   bht_reg_28_20_inst : DLH_X1 port map( G => N2272, D => N3773, Q => 
                           bht_28_20_port);
   bht_reg_30_20_inst : DLH_X1 port map( G => N2164, D => N3773, Q => 
                           bht_30_20_port);
   bht_reg_31_20_inst : DLH_X1 port map( G => N2110, D => N3773, Q => 
                           bht_31_20_port);
   bht_reg_29_20_inst : DLH_X1 port map( G => N2218, D => N3773, Q => 
                           bht_29_20_port);
   bht_reg_27_20_inst : DLH_X1 port map( G => N2326, D => N3773, Q => 
                           bht_27_20_port);
   bht_reg_25_20_inst : DLH_X1 port map( G => N2434, D => N3773, Q => 
                           bht_25_20_port);
   bht_reg_23_20_inst : DLH_X1 port map( G => N2542, D => N3773, Q => 
                           bht_23_20_port);
   bht_reg_21_20_inst : DLH_X1 port map( G => N2650, D => N3773, Q => 
                           bht_21_20_port);
   bht_reg_19_20_inst : DLH_X1 port map( G => N2758, D => N3773, Q => 
                           bht_19_20_port);
   bht_reg_17_20_inst : DLH_X1 port map( G => N2866, D => N3773, Q => 
                           bht_17_20_port);
   bht_reg_15_20_inst : DLH_X1 port map( G => N2974, D => N3773, Q => 
                           bht_15_20_port);
   bht_reg_13_20_inst : DLH_X1 port map( G => N3082, D => N3773, Q => 
                           bht_13_20_port);
   bht_reg_11_20_inst : DLH_X1 port map( G => N3190, D => N3773, Q => 
                           bht_11_20_port);
   bht_reg_9_20_inst : DLH_X1 port map( G => N3298, D => N3773, Q => 
                           bht_9_20_port);
   bht_reg_7_20_inst : DLH_X1 port map( G => N3406, D => N3773, Q => 
                           bht_7_20_port);
   bht_reg_5_20_inst : DLH_X1 port map( G => N3514, D => N3773, Q => 
                           bht_5_20_port);
   bht_reg_3_20_inst : DLH_X1 port map( G => N3622, D => N3773, Q => 
                           bht_3_20_port);
   bht_reg_1_20_inst : DLH_X1 port map( G => N3730, D => N3773, Q => 
                           bht_1_20_port);
   entry_r_reg_19_inst : DLH_X1 port map( G => N188, D => N144, Q => 
                           entry_r_19_port);
   entry_r_delay_reg_19_inst : DFFR_X1 port map( D => entry_r_19_port, CK => 
                           clk, RN => rst, Q => net108084, QN => n27);
   bht_reg_0_19_inst : DLH_X1 port map( G => N3784, D => N3771, Q => 
                           bht_0_19_port);
   bht_reg_2_19_inst : DLH_X1 port map( G => N3676, D => N3771, Q => 
                           bht_2_19_port);
   bht_reg_4_19_inst : DLH_X1 port map( G => N3568, D => N3771, Q => 
                           bht_4_19_port);
   bht_reg_6_19_inst : DLH_X1 port map( G => N3460, D => N3771, Q => 
                           bht_6_19_port);
   bht_reg_8_19_inst : DLH_X1 port map( G => N3352, D => N3771, Q => 
                           bht_8_19_port);
   bht_reg_10_19_inst : DLH_X1 port map( G => N3244, D => N3771, Q => 
                           bht_10_19_port);
   bht_reg_12_19_inst : DLH_X1 port map( G => N3136, D => N3771, Q => 
                           bht_12_19_port);
   bht_reg_14_19_inst : DLH_X1 port map( G => N3028, D => N3771, Q => 
                           bht_14_19_port);
   bht_reg_16_19_inst : DLH_X1 port map( G => N2920, D => N3771, Q => 
                           bht_16_19_port);
   bht_reg_18_19_inst : DLH_X1 port map( G => N2812, D => N3771, Q => 
                           bht_18_19_port);
   bht_reg_20_19_inst : DLH_X1 port map( G => N2704, D => N3771, Q => 
                           bht_20_19_port);
   bht_reg_22_19_inst : DLH_X1 port map( G => N2596, D => N3771, Q => 
                           bht_22_19_port);
   bht_reg_24_19_inst : DLH_X1 port map( G => N2488, D => N3771, Q => 
                           bht_24_19_port);
   bht_reg_26_19_inst : DLH_X1 port map( G => N2380, D => N3771, Q => 
                           bht_26_19_port);
   bht_reg_28_19_inst : DLH_X1 port map( G => N2272, D => N3771, Q => 
                           bht_28_19_port);
   bht_reg_30_19_inst : DLH_X1 port map( G => N2164, D => N3771, Q => 
                           bht_30_19_port);
   bht_reg_31_19_inst : DLH_X1 port map( G => N2110, D => N3771, Q => 
                           bht_31_19_port);
   bht_reg_29_19_inst : DLH_X1 port map( G => N2218, D => N3771, Q => 
                           bht_29_19_port);
   bht_reg_27_19_inst : DLH_X1 port map( G => N2326, D => N3771, Q => 
                           bht_27_19_port);
   bht_reg_25_19_inst : DLH_X1 port map( G => N2434, D => N3771, Q => 
                           bht_25_19_port);
   bht_reg_23_19_inst : DLH_X1 port map( G => N2542, D => N3771, Q => 
                           bht_23_19_port);
   bht_reg_21_19_inst : DLH_X1 port map( G => N2650, D => N3771, Q => 
                           bht_21_19_port);
   bht_reg_19_19_inst : DLH_X1 port map( G => N2758, D => N3771, Q => 
                           bht_19_19_port);
   bht_reg_17_19_inst : DLH_X1 port map( G => N2866, D => N3771, Q => 
                           bht_17_19_port);
   bht_reg_15_19_inst : DLH_X1 port map( G => N2974, D => N3771, Q => 
                           bht_15_19_port);
   bht_reg_13_19_inst : DLH_X1 port map( G => N3082, D => N3771, Q => 
                           bht_13_19_port);
   bht_reg_11_19_inst : DLH_X1 port map( G => N3190, D => N3771, Q => 
                           bht_11_19_port);
   bht_reg_9_19_inst : DLH_X1 port map( G => N3298, D => N3771, Q => 
                           bht_9_19_port);
   bht_reg_7_19_inst : DLH_X1 port map( G => N3406, D => N3771, Q => 
                           bht_7_19_port);
   bht_reg_5_19_inst : DLH_X1 port map( G => N3514, D => N3771, Q => 
                           bht_5_19_port);
   bht_reg_3_19_inst : DLH_X1 port map( G => N3622, D => N3771, Q => 
                           bht_3_19_port);
   bht_reg_1_19_inst : DLH_X1 port map( G => N3730, D => N3771, Q => 
                           bht_1_19_port);
   entry_r_reg_18_inst : DLH_X1 port map( G => N188, D => N143, Q => 
                           entry_r_18_port);
   entry_r_delay_reg_18_inst : DFFR_X1 port map( D => entry_r_18_port, CK => 
                           clk, RN => rst, Q => net108083, QN => n26);
   bht_reg_0_18_inst : DLH_X1 port map( G => N3784, D => N3769, Q => 
                           bht_0_18_port);
   bht_reg_2_18_inst : DLH_X1 port map( G => N3676, D => N3769, Q => 
                           bht_2_18_port);
   bht_reg_4_18_inst : DLH_X1 port map( G => N3568, D => N3769, Q => 
                           bht_4_18_port);
   bht_reg_6_18_inst : DLH_X1 port map( G => N3460, D => N3769, Q => 
                           bht_6_18_port);
   bht_reg_8_18_inst : DLH_X1 port map( G => N3352, D => N3769, Q => 
                           bht_8_18_port);
   bht_reg_10_18_inst : DLH_X1 port map( G => N3244, D => N3769, Q => 
                           bht_10_18_port);
   bht_reg_12_18_inst : DLH_X1 port map( G => N3136, D => N3769, Q => 
                           bht_12_18_port);
   bht_reg_14_18_inst : DLH_X1 port map( G => N3028, D => N3769, Q => 
                           bht_14_18_port);
   bht_reg_16_18_inst : DLH_X1 port map( G => N2920, D => N3769, Q => 
                           bht_16_18_port);
   bht_reg_18_18_inst : DLH_X1 port map( G => N2812, D => N3769, Q => 
                           bht_18_18_port);
   bht_reg_20_18_inst : DLH_X1 port map( G => N2704, D => N3769, Q => 
                           bht_20_18_port);
   bht_reg_22_18_inst : DLH_X1 port map( G => N2596, D => N3769, Q => 
                           bht_22_18_port);
   bht_reg_24_18_inst : DLH_X1 port map( G => N2488, D => N3769, Q => 
                           bht_24_18_port);
   bht_reg_26_18_inst : DLH_X1 port map( G => N2380, D => N3769, Q => 
                           bht_26_18_port);
   bht_reg_28_18_inst : DLH_X1 port map( G => N2272, D => N3769, Q => 
                           bht_28_18_port);
   bht_reg_30_18_inst : DLH_X1 port map( G => N2164, D => N3769, Q => 
                           bht_30_18_port);
   bht_reg_31_18_inst : DLH_X1 port map( G => N2110, D => N3769, Q => 
                           bht_31_18_port);
   bht_reg_29_18_inst : DLH_X1 port map( G => N2218, D => N3769, Q => 
                           bht_29_18_port);
   bht_reg_27_18_inst : DLH_X1 port map( G => N2326, D => N3769, Q => 
                           bht_27_18_port);
   bht_reg_25_18_inst : DLH_X1 port map( G => N2434, D => N3769, Q => 
                           bht_25_18_port);
   bht_reg_23_18_inst : DLH_X1 port map( G => N2542, D => N3769, Q => 
                           bht_23_18_port);
   bht_reg_21_18_inst : DLH_X1 port map( G => N2650, D => N3769, Q => 
                           bht_21_18_port);
   bht_reg_19_18_inst : DLH_X1 port map( G => N2758, D => N3769, Q => 
                           bht_19_18_port);
   bht_reg_17_18_inst : DLH_X1 port map( G => N2866, D => N3769, Q => 
                           bht_17_18_port);
   bht_reg_15_18_inst : DLH_X1 port map( G => N2974, D => N3769, Q => 
                           bht_15_18_port);
   bht_reg_13_18_inst : DLH_X1 port map( G => N3082, D => N3769, Q => 
                           bht_13_18_port);
   bht_reg_11_18_inst : DLH_X1 port map( G => N3190, D => N3769, Q => 
                           bht_11_18_port);
   bht_reg_9_18_inst : DLH_X1 port map( G => N3298, D => N3769, Q => 
                           bht_9_18_port);
   bht_reg_7_18_inst : DLH_X1 port map( G => N3406, D => N3769, Q => 
                           bht_7_18_port);
   bht_reg_5_18_inst : DLH_X1 port map( G => N3514, D => N3769, Q => 
                           bht_5_18_port);
   bht_reg_3_18_inst : DLH_X1 port map( G => N3622, D => N3769, Q => 
                           bht_3_18_port);
   bht_reg_1_18_inst : DLH_X1 port map( G => N3730, D => N3769, Q => 
                           bht_1_18_port);
   entry_r_reg_17_inst : DLH_X1 port map( G => N188, D => N142, Q => 
                           entry_r_17_port);
   entry_r_delay_reg_17_inst : DFFR_X1 port map( D => entry_r_17_port, CK => 
                           clk, RN => rst, Q => net108082, QN => n25);
   bht_reg_0_17_inst : DLH_X1 port map( G => N3784, D => N3767, Q => 
                           bht_0_17_port);
   bht_reg_2_17_inst : DLH_X1 port map( G => N3676, D => N3767, Q => 
                           bht_2_17_port);
   bht_reg_4_17_inst : DLH_X1 port map( G => N3568, D => N3767, Q => 
                           bht_4_17_port);
   bht_reg_6_17_inst : DLH_X1 port map( G => N3460, D => N3767, Q => 
                           bht_6_17_port);
   bht_reg_8_17_inst : DLH_X1 port map( G => N3352, D => N3767, Q => 
                           bht_8_17_port);
   bht_reg_10_17_inst : DLH_X1 port map( G => N3244, D => N3767, Q => 
                           bht_10_17_port);
   bht_reg_12_17_inst : DLH_X1 port map( G => N3136, D => N3767, Q => 
                           bht_12_17_port);
   bht_reg_14_17_inst : DLH_X1 port map( G => N3028, D => N3767, Q => 
                           bht_14_17_port);
   bht_reg_16_17_inst : DLH_X1 port map( G => N2920, D => N3767, Q => 
                           bht_16_17_port);
   bht_reg_18_17_inst : DLH_X1 port map( G => N2812, D => N3767, Q => 
                           bht_18_17_port);
   bht_reg_20_17_inst : DLH_X1 port map( G => N2704, D => N3767, Q => 
                           bht_20_17_port);
   bht_reg_22_17_inst : DLH_X1 port map( G => N2596, D => N3767, Q => 
                           bht_22_17_port);
   bht_reg_24_17_inst : DLH_X1 port map( G => N2488, D => N3767, Q => 
                           bht_24_17_port);
   bht_reg_26_17_inst : DLH_X1 port map( G => N2380, D => N3767, Q => 
                           bht_26_17_port);
   bht_reg_28_17_inst : DLH_X1 port map( G => N2272, D => N3767, Q => 
                           bht_28_17_port);
   bht_reg_30_17_inst : DLH_X1 port map( G => N2164, D => N3767, Q => 
                           bht_30_17_port);
   bht_reg_31_17_inst : DLH_X1 port map( G => N2110, D => N3767, Q => 
                           bht_31_17_port);
   bht_reg_29_17_inst : DLH_X1 port map( G => N2218, D => N3767, Q => 
                           bht_29_17_port);
   bht_reg_27_17_inst : DLH_X1 port map( G => N2326, D => N3767, Q => 
                           bht_27_17_port);
   bht_reg_25_17_inst : DLH_X1 port map( G => N2434, D => N3767, Q => 
                           bht_25_17_port);
   bht_reg_23_17_inst : DLH_X1 port map( G => N2542, D => N3767, Q => 
                           bht_23_17_port);
   bht_reg_21_17_inst : DLH_X1 port map( G => N2650, D => N3767, Q => 
                           bht_21_17_port);
   bht_reg_19_17_inst : DLH_X1 port map( G => N2758, D => N3767, Q => 
                           bht_19_17_port);
   bht_reg_17_17_inst : DLH_X1 port map( G => N2866, D => N3767, Q => 
                           bht_17_17_port);
   bht_reg_15_17_inst : DLH_X1 port map( G => N2974, D => N3767, Q => 
                           bht_15_17_port);
   bht_reg_13_17_inst : DLH_X1 port map( G => N3082, D => N3767, Q => 
                           bht_13_17_port);
   bht_reg_11_17_inst : DLH_X1 port map( G => N3190, D => N3767, Q => 
                           bht_11_17_port);
   bht_reg_9_17_inst : DLH_X1 port map( G => N3298, D => N3767, Q => 
                           bht_9_17_port);
   bht_reg_7_17_inst : DLH_X1 port map( G => N3406, D => N3767, Q => 
                           bht_7_17_port);
   bht_reg_5_17_inst : DLH_X1 port map( G => N3514, D => N3767, Q => 
                           bht_5_17_port);
   bht_reg_3_17_inst : DLH_X1 port map( G => N3622, D => N3767, Q => 
                           bht_3_17_port);
   bht_reg_1_17_inst : DLH_X1 port map( G => N3730, D => N3767, Q => 
                           bht_1_17_port);
   entry_r_reg_16_inst : DLH_X1 port map( G => N188, D => N141, Q => 
                           entry_r_16_port);
   entry_r_delay_reg_16_inst : DFFR_X1 port map( D => entry_r_16_port, CK => 
                           clk, RN => rst, Q => net108081, QN => n24);
   bht_reg_0_16_inst : DLH_X1 port map( G => N3784, D => N3765, Q => 
                           bht_0_16_port);
   bht_reg_2_16_inst : DLH_X1 port map( G => N3676, D => N3765, Q => 
                           bht_2_16_port);
   bht_reg_4_16_inst : DLH_X1 port map( G => N3568, D => N3765, Q => 
                           bht_4_16_port);
   bht_reg_6_16_inst : DLH_X1 port map( G => N3460, D => N3765, Q => 
                           bht_6_16_port);
   bht_reg_8_16_inst : DLH_X1 port map( G => N3352, D => N3765, Q => 
                           bht_8_16_port);
   bht_reg_10_16_inst : DLH_X1 port map( G => N3244, D => N3765, Q => 
                           bht_10_16_port);
   bht_reg_12_16_inst : DLH_X1 port map( G => N3136, D => N3765, Q => 
                           bht_12_16_port);
   bht_reg_14_16_inst : DLH_X1 port map( G => N3028, D => N3765, Q => 
                           bht_14_16_port);
   bht_reg_16_16_inst : DLH_X1 port map( G => N2920, D => N3765, Q => 
                           bht_16_16_port);
   bht_reg_18_16_inst : DLH_X1 port map( G => N2812, D => N3765, Q => 
                           bht_18_16_port);
   bht_reg_20_16_inst : DLH_X1 port map( G => N2704, D => N3765, Q => 
                           bht_20_16_port);
   bht_reg_22_16_inst : DLH_X1 port map( G => N2596, D => N3765, Q => 
                           bht_22_16_port);
   bht_reg_24_16_inst : DLH_X1 port map( G => N2488, D => N3765, Q => 
                           bht_24_16_port);
   bht_reg_26_16_inst : DLH_X1 port map( G => N2380, D => N3765, Q => 
                           bht_26_16_port);
   bht_reg_28_16_inst : DLH_X1 port map( G => N2272, D => N3765, Q => 
                           bht_28_16_port);
   bht_reg_30_16_inst : DLH_X1 port map( G => N2164, D => N3765, Q => 
                           bht_30_16_port);
   bht_reg_31_16_inst : DLH_X1 port map( G => N2110, D => N3765, Q => 
                           bht_31_16_port);
   bht_reg_29_16_inst : DLH_X1 port map( G => N2218, D => N3765, Q => 
                           bht_29_16_port);
   bht_reg_27_16_inst : DLH_X1 port map( G => N2326, D => N3765, Q => 
                           bht_27_16_port);
   bht_reg_25_16_inst : DLH_X1 port map( G => N2434, D => N3765, Q => 
                           bht_25_16_port);
   bht_reg_23_16_inst : DLH_X1 port map( G => N2542, D => N3765, Q => 
                           bht_23_16_port);
   bht_reg_21_16_inst : DLH_X1 port map( G => N2650, D => N3765, Q => 
                           bht_21_16_port);
   bht_reg_19_16_inst : DLH_X1 port map( G => N2758, D => N3765, Q => 
                           bht_19_16_port);
   bht_reg_17_16_inst : DLH_X1 port map( G => N2866, D => N3765, Q => 
                           bht_17_16_port);
   bht_reg_15_16_inst : DLH_X1 port map( G => N2974, D => N3765, Q => 
                           bht_15_16_port);
   bht_reg_13_16_inst : DLH_X1 port map( G => N3082, D => N3765, Q => 
                           bht_13_16_port);
   bht_reg_11_16_inst : DLH_X1 port map( G => N3190, D => N3765, Q => 
                           bht_11_16_port);
   bht_reg_9_16_inst : DLH_X1 port map( G => N3298, D => N3765, Q => 
                           bht_9_16_port);
   bht_reg_7_16_inst : DLH_X1 port map( G => N3406, D => N3765, Q => 
                           bht_7_16_port);
   bht_reg_5_16_inst : DLH_X1 port map( G => N3514, D => N3765, Q => 
                           bht_5_16_port);
   bht_reg_3_16_inst : DLH_X1 port map( G => N3622, D => N3765, Q => 
                           bht_3_16_port);
   bht_reg_1_16_inst : DLH_X1 port map( G => N3730, D => N3765, Q => 
                           bht_1_16_port);
   entry_r_reg_15_inst : DLH_X1 port map( G => N188, D => N140, Q => 
                           entry_r_15_port);
   entry_r_delay_reg_15_inst : DFFR_X1 port map( D => entry_r_15_port, CK => 
                           clk, RN => rst, Q => net108080, QN => n23);
   bht_reg_0_15_inst : DLH_X1 port map( G => N3784, D => N3763, Q => 
                           bht_0_15_port);
   bht_reg_2_15_inst : DLH_X1 port map( G => N3676, D => N3763, Q => 
                           bht_2_15_port);
   bht_reg_4_15_inst : DLH_X1 port map( G => N3568, D => N3763, Q => 
                           bht_4_15_port);
   bht_reg_6_15_inst : DLH_X1 port map( G => N3460, D => N3763, Q => 
                           bht_6_15_port);
   bht_reg_8_15_inst : DLH_X1 port map( G => N3352, D => N3763, Q => 
                           bht_8_15_port);
   bht_reg_10_15_inst : DLH_X1 port map( G => N3244, D => N3763, Q => 
                           bht_10_15_port);
   bht_reg_12_15_inst : DLH_X1 port map( G => N3136, D => N3763, Q => 
                           bht_12_15_port);
   bht_reg_14_15_inst : DLH_X1 port map( G => N3028, D => N3763, Q => 
                           bht_14_15_port);
   bht_reg_16_15_inst : DLH_X1 port map( G => N2920, D => N3763, Q => 
                           bht_16_15_port);
   bht_reg_18_15_inst : DLH_X1 port map( G => N2812, D => N3763, Q => 
                           bht_18_15_port);
   bht_reg_20_15_inst : DLH_X1 port map( G => N2704, D => N3763, Q => 
                           bht_20_15_port);
   bht_reg_22_15_inst : DLH_X1 port map( G => N2596, D => N3763, Q => 
                           bht_22_15_port);
   bht_reg_24_15_inst : DLH_X1 port map( G => N2488, D => N3763, Q => 
                           bht_24_15_port);
   bht_reg_26_15_inst : DLH_X1 port map( G => N2380, D => N3763, Q => 
                           bht_26_15_port);
   bht_reg_28_15_inst : DLH_X1 port map( G => N2272, D => N3763, Q => 
                           bht_28_15_port);
   bht_reg_30_15_inst : DLH_X1 port map( G => N2164, D => N3763, Q => 
                           bht_30_15_port);
   bht_reg_31_15_inst : DLH_X1 port map( G => N2110, D => N3763, Q => 
                           bht_31_15_port);
   bht_reg_29_15_inst : DLH_X1 port map( G => N2218, D => N3763, Q => 
                           bht_29_15_port);
   bht_reg_27_15_inst : DLH_X1 port map( G => N2326, D => N3763, Q => 
                           bht_27_15_port);
   bht_reg_25_15_inst : DLH_X1 port map( G => N2434, D => N3763, Q => 
                           bht_25_15_port);
   bht_reg_23_15_inst : DLH_X1 port map( G => N2542, D => N3763, Q => 
                           bht_23_15_port);
   bht_reg_21_15_inst : DLH_X1 port map( G => N2650, D => N3763, Q => 
                           bht_21_15_port);
   bht_reg_19_15_inst : DLH_X1 port map( G => N2758, D => N3763, Q => 
                           bht_19_15_port);
   bht_reg_17_15_inst : DLH_X1 port map( G => N2866, D => N3763, Q => 
                           bht_17_15_port);
   bht_reg_15_15_inst : DLH_X1 port map( G => N2974, D => N3763, Q => 
                           bht_15_15_port);
   bht_reg_13_15_inst : DLH_X1 port map( G => N3082, D => N3763, Q => 
                           bht_13_15_port);
   bht_reg_11_15_inst : DLH_X1 port map( G => N3190, D => N3763, Q => 
                           bht_11_15_port);
   bht_reg_9_15_inst : DLH_X1 port map( G => N3298, D => N3763, Q => 
                           bht_9_15_port);
   bht_reg_7_15_inst : DLH_X1 port map( G => N3406, D => N3763, Q => 
                           bht_7_15_port);
   bht_reg_5_15_inst : DLH_X1 port map( G => N3514, D => N3763, Q => 
                           bht_5_15_port);
   bht_reg_3_15_inst : DLH_X1 port map( G => N3622, D => N3763, Q => 
                           bht_3_15_port);
   bht_reg_1_15_inst : DLH_X1 port map( G => N3730, D => N3763, Q => 
                           bht_1_15_port);
   entry_r_reg_14_inst : DLH_X1 port map( G => N188, D => N139, Q => 
                           entry_r_14_port);
   entry_r_delay_reg_14_inst : DFFR_X1 port map( D => entry_r_14_port, CK => 
                           clk, RN => rst, Q => net108079, QN => n22);
   bht_reg_0_14_inst : DLH_X1 port map( G => N3784, D => N3761, Q => 
                           bht_0_14_port);
   bht_reg_2_14_inst : DLH_X1 port map( G => N3676, D => N3761, Q => 
                           bht_2_14_port);
   bht_reg_4_14_inst : DLH_X1 port map( G => N3568, D => N3761, Q => 
                           bht_4_14_port);
   bht_reg_6_14_inst : DLH_X1 port map( G => N3460, D => N3761, Q => 
                           bht_6_14_port);
   bht_reg_8_14_inst : DLH_X1 port map( G => N3352, D => N3761, Q => 
                           bht_8_14_port);
   bht_reg_10_14_inst : DLH_X1 port map( G => N3244, D => N3761, Q => 
                           bht_10_14_port);
   bht_reg_12_14_inst : DLH_X1 port map( G => N3136, D => N3761, Q => 
                           bht_12_14_port);
   bht_reg_14_14_inst : DLH_X1 port map( G => N3028, D => N3761, Q => 
                           bht_14_14_port);
   bht_reg_16_14_inst : DLH_X1 port map( G => N2920, D => N3761, Q => 
                           bht_16_14_port);
   bht_reg_18_14_inst : DLH_X1 port map( G => N2812, D => N3761, Q => 
                           bht_18_14_port);
   bht_reg_20_14_inst : DLH_X1 port map( G => N2704, D => N3761, Q => 
                           bht_20_14_port);
   bht_reg_22_14_inst : DLH_X1 port map( G => N2596, D => N3761, Q => 
                           bht_22_14_port);
   bht_reg_24_14_inst : DLH_X1 port map( G => N2488, D => N3761, Q => 
                           bht_24_14_port);
   bht_reg_26_14_inst : DLH_X1 port map( G => N2380, D => N3761, Q => 
                           bht_26_14_port);
   bht_reg_28_14_inst : DLH_X1 port map( G => N2272, D => N3761, Q => 
                           bht_28_14_port);
   bht_reg_30_14_inst : DLH_X1 port map( G => N2164, D => N3761, Q => 
                           bht_30_14_port);
   bht_reg_31_14_inst : DLH_X1 port map( G => N2110, D => N3761, Q => 
                           bht_31_14_port);
   bht_reg_29_14_inst : DLH_X1 port map( G => N2218, D => N3761, Q => 
                           bht_29_14_port);
   bht_reg_27_14_inst : DLH_X1 port map( G => N2326, D => N3761, Q => 
                           bht_27_14_port);
   bht_reg_25_14_inst : DLH_X1 port map( G => N2434, D => N3761, Q => 
                           bht_25_14_port);
   bht_reg_23_14_inst : DLH_X1 port map( G => N2542, D => N3761, Q => 
                           bht_23_14_port);
   bht_reg_21_14_inst : DLH_X1 port map( G => N2650, D => N3761, Q => 
                           bht_21_14_port);
   bht_reg_19_14_inst : DLH_X1 port map( G => N2758, D => N3761, Q => 
                           bht_19_14_port);
   bht_reg_17_14_inst : DLH_X1 port map( G => N2866, D => N3761, Q => 
                           bht_17_14_port);
   bht_reg_15_14_inst : DLH_X1 port map( G => N2974, D => N3761, Q => 
                           bht_15_14_port);
   bht_reg_13_14_inst : DLH_X1 port map( G => N3082, D => N3761, Q => 
                           bht_13_14_port);
   bht_reg_11_14_inst : DLH_X1 port map( G => N3190, D => N3761, Q => 
                           bht_11_14_port);
   bht_reg_9_14_inst : DLH_X1 port map( G => N3298, D => N3761, Q => 
                           bht_9_14_port);
   bht_reg_7_14_inst : DLH_X1 port map( G => N3406, D => N3761, Q => 
                           bht_7_14_port);
   bht_reg_5_14_inst : DLH_X1 port map( G => N3514, D => N3761, Q => 
                           bht_5_14_port);
   bht_reg_3_14_inst : DLH_X1 port map( G => N3622, D => N3761, Q => 
                           bht_3_14_port);
   bht_reg_1_14_inst : DLH_X1 port map( G => N3730, D => N3761, Q => 
                           bht_1_14_port);
   entry_r_reg_13_inst : DLH_X1 port map( G => N188, D => N138, Q => 
                           entry_r_13_port);
   entry_r_delay_reg_13_inst : DFFR_X1 port map( D => entry_r_13_port, CK => 
                           clk, RN => rst, Q => net108078, QN => n21);
   bht_reg_0_13_inst : DLH_X1 port map( G => N3784, D => N3759, Q => 
                           bht_0_13_port);
   bht_reg_2_13_inst : DLH_X1 port map( G => N3676, D => N3759, Q => 
                           bht_2_13_port);
   bht_reg_4_13_inst : DLH_X1 port map( G => N3568, D => N3759, Q => 
                           bht_4_13_port);
   bht_reg_6_13_inst : DLH_X1 port map( G => N3460, D => N3759, Q => 
                           bht_6_13_port);
   bht_reg_8_13_inst : DLH_X1 port map( G => N3352, D => N3759, Q => 
                           bht_8_13_port);
   bht_reg_10_13_inst : DLH_X1 port map( G => N3244, D => N3759, Q => 
                           bht_10_13_port);
   bht_reg_12_13_inst : DLH_X1 port map( G => N3136, D => N3759, Q => 
                           bht_12_13_port);
   bht_reg_14_13_inst : DLH_X1 port map( G => N3028, D => N3759, Q => 
                           bht_14_13_port);
   bht_reg_16_13_inst : DLH_X1 port map( G => N2920, D => N3759, Q => 
                           bht_16_13_port);
   bht_reg_18_13_inst : DLH_X1 port map( G => N2812, D => N3759, Q => 
                           bht_18_13_port);
   bht_reg_20_13_inst : DLH_X1 port map( G => N2704, D => N3759, Q => 
                           bht_20_13_port);
   bht_reg_22_13_inst : DLH_X1 port map( G => N2596, D => N3759, Q => 
                           bht_22_13_port);
   bht_reg_24_13_inst : DLH_X1 port map( G => N2488, D => N3759, Q => 
                           bht_24_13_port);
   bht_reg_26_13_inst : DLH_X1 port map( G => N2380, D => N3759, Q => 
                           bht_26_13_port);
   bht_reg_28_13_inst : DLH_X1 port map( G => N2272, D => N3759, Q => 
                           bht_28_13_port);
   bht_reg_30_13_inst : DLH_X1 port map( G => N2164, D => N3759, Q => 
                           bht_30_13_port);
   bht_reg_31_13_inst : DLH_X1 port map( G => N2110, D => N3759, Q => 
                           bht_31_13_port);
   bht_reg_29_13_inst : DLH_X1 port map( G => N2218, D => N3759, Q => 
                           bht_29_13_port);
   bht_reg_27_13_inst : DLH_X1 port map( G => N2326, D => N3759, Q => 
                           bht_27_13_port);
   bht_reg_25_13_inst : DLH_X1 port map( G => N2434, D => N3759, Q => 
                           bht_25_13_port);
   bht_reg_23_13_inst : DLH_X1 port map( G => N2542, D => N3759, Q => 
                           bht_23_13_port);
   bht_reg_21_13_inst : DLH_X1 port map( G => N2650, D => N3759, Q => 
                           bht_21_13_port);
   bht_reg_19_13_inst : DLH_X1 port map( G => N2758, D => N3759, Q => 
                           bht_19_13_port);
   bht_reg_17_13_inst : DLH_X1 port map( G => N2866, D => N3759, Q => 
                           bht_17_13_port);
   bht_reg_15_13_inst : DLH_X1 port map( G => N2974, D => N3759, Q => 
                           bht_15_13_port);
   bht_reg_13_13_inst : DLH_X1 port map( G => N3082, D => N3759, Q => 
                           bht_13_13_port);
   bht_reg_11_13_inst : DLH_X1 port map( G => N3190, D => N3759, Q => 
                           bht_11_13_port);
   bht_reg_9_13_inst : DLH_X1 port map( G => N3298, D => N3759, Q => 
                           bht_9_13_port);
   bht_reg_7_13_inst : DLH_X1 port map( G => N3406, D => N3759, Q => 
                           bht_7_13_port);
   bht_reg_5_13_inst : DLH_X1 port map( G => N3514, D => N3759, Q => 
                           bht_5_13_port);
   bht_reg_3_13_inst : DLH_X1 port map( G => N3622, D => N3759, Q => 
                           bht_3_13_port);
   bht_reg_1_13_inst : DLH_X1 port map( G => N3730, D => N3759, Q => 
                           bht_1_13_port);
   entry_r_reg_12_inst : DLH_X1 port map( G => N188, D => N137, Q => 
                           entry_r_12_port);
   entry_r_delay_reg_12_inst : DFFR_X1 port map( D => entry_r_12_port, CK => 
                           clk, RN => rst, Q => net108077, QN => n20);
   bht_reg_0_12_inst : DLH_X1 port map( G => N3784, D => N3757, Q => 
                           bht_0_12_port);
   bht_reg_2_12_inst : DLH_X1 port map( G => N3676, D => N3757, Q => 
                           bht_2_12_port);
   bht_reg_4_12_inst : DLH_X1 port map( G => N3568, D => N3757, Q => 
                           bht_4_12_port);
   bht_reg_6_12_inst : DLH_X1 port map( G => N3460, D => N3757, Q => 
                           bht_6_12_port);
   bht_reg_8_12_inst : DLH_X1 port map( G => N3352, D => N3757, Q => 
                           bht_8_12_port);
   bht_reg_10_12_inst : DLH_X1 port map( G => N3244, D => N3757, Q => 
                           bht_10_12_port);
   bht_reg_12_12_inst : DLH_X1 port map( G => N3136, D => N3757, Q => 
                           bht_12_12_port);
   bht_reg_14_12_inst : DLH_X1 port map( G => N3028, D => N3757, Q => 
                           bht_14_12_port);
   bht_reg_16_12_inst : DLH_X1 port map( G => N2920, D => N3757, Q => 
                           bht_16_12_port);
   bht_reg_18_12_inst : DLH_X1 port map( G => N2812, D => N3757, Q => 
                           bht_18_12_port);
   bht_reg_20_12_inst : DLH_X1 port map( G => N2704, D => N3757, Q => 
                           bht_20_12_port);
   bht_reg_22_12_inst : DLH_X1 port map( G => N2596, D => N3757, Q => 
                           bht_22_12_port);
   bht_reg_24_12_inst : DLH_X1 port map( G => N2488, D => N3757, Q => 
                           bht_24_12_port);
   bht_reg_26_12_inst : DLH_X1 port map( G => N2380, D => N3757, Q => 
                           bht_26_12_port);
   bht_reg_28_12_inst : DLH_X1 port map( G => N2272, D => N3757, Q => 
                           bht_28_12_port);
   bht_reg_30_12_inst : DLH_X1 port map( G => N2164, D => N3757, Q => 
                           bht_30_12_port);
   bht_reg_31_12_inst : DLH_X1 port map( G => N2110, D => N3757, Q => 
                           bht_31_12_port);
   bht_reg_29_12_inst : DLH_X1 port map( G => N2218, D => N3757, Q => 
                           bht_29_12_port);
   bht_reg_27_12_inst : DLH_X1 port map( G => N2326, D => N3757, Q => 
                           bht_27_12_port);
   bht_reg_25_12_inst : DLH_X1 port map( G => N2434, D => N3757, Q => 
                           bht_25_12_port);
   bht_reg_23_12_inst : DLH_X1 port map( G => N2542, D => N3757, Q => 
                           bht_23_12_port);
   bht_reg_21_12_inst : DLH_X1 port map( G => N2650, D => N3757, Q => 
                           bht_21_12_port);
   bht_reg_19_12_inst : DLH_X1 port map( G => N2758, D => N3757, Q => 
                           bht_19_12_port);
   bht_reg_17_12_inst : DLH_X1 port map( G => N2866, D => N3757, Q => 
                           bht_17_12_port);
   bht_reg_15_12_inst : DLH_X1 port map( G => N2974, D => N3757, Q => 
                           bht_15_12_port);
   bht_reg_13_12_inst : DLH_X1 port map( G => N3082, D => N3757, Q => 
                           bht_13_12_port);
   bht_reg_11_12_inst : DLH_X1 port map( G => N3190, D => N3757, Q => 
                           bht_11_12_port);
   bht_reg_9_12_inst : DLH_X1 port map( G => N3298, D => N3757, Q => 
                           bht_9_12_port);
   bht_reg_7_12_inst : DLH_X1 port map( G => N3406, D => N3757, Q => 
                           bht_7_12_port);
   bht_reg_5_12_inst : DLH_X1 port map( G => N3514, D => N3757, Q => 
                           bht_5_12_port);
   bht_reg_3_12_inst : DLH_X1 port map( G => N3622, D => N3757, Q => 
                           bht_3_12_port);
   bht_reg_1_12_inst : DLH_X1 port map( G => N3730, D => N3757, Q => 
                           bht_1_12_port);
   entry_r_reg_11_inst : DLH_X1 port map( G => N188, D => N136, Q => 
                           entry_r_11_port);
   entry_r_delay_reg_11_inst : DFFR_X1 port map( D => entry_r_11_port, CK => 
                           clk, RN => rst, Q => net108076, QN => n19);
   bht_reg_0_11_inst : DLH_X1 port map( G => N3784, D => N3755, Q => 
                           bht_0_11_port);
   bht_reg_2_11_inst : DLH_X1 port map( G => N3676, D => N3755, Q => 
                           bht_2_11_port);
   bht_reg_4_11_inst : DLH_X1 port map( G => N3568, D => N3755, Q => 
                           bht_4_11_port);
   bht_reg_6_11_inst : DLH_X1 port map( G => N3460, D => N3755, Q => 
                           bht_6_11_port);
   bht_reg_8_11_inst : DLH_X1 port map( G => N3352, D => N3755, Q => 
                           bht_8_11_port);
   bht_reg_10_11_inst : DLH_X1 port map( G => N3244, D => N3755, Q => 
                           bht_10_11_port);
   bht_reg_12_11_inst : DLH_X1 port map( G => N3136, D => N3755, Q => 
                           bht_12_11_port);
   bht_reg_14_11_inst : DLH_X1 port map( G => N3028, D => N3755, Q => 
                           bht_14_11_port);
   bht_reg_16_11_inst : DLH_X1 port map( G => N2920, D => N3755, Q => 
                           bht_16_11_port);
   bht_reg_18_11_inst : DLH_X1 port map( G => N2812, D => N3755, Q => 
                           bht_18_11_port);
   bht_reg_20_11_inst : DLH_X1 port map( G => N2704, D => N3755, Q => 
                           bht_20_11_port);
   bht_reg_22_11_inst : DLH_X1 port map( G => N2596, D => N3755, Q => 
                           bht_22_11_port);
   bht_reg_24_11_inst : DLH_X1 port map( G => N2488, D => N3755, Q => 
                           bht_24_11_port);
   bht_reg_26_11_inst : DLH_X1 port map( G => N2380, D => N3755, Q => 
                           bht_26_11_port);
   bht_reg_28_11_inst : DLH_X1 port map( G => N2272, D => N3755, Q => 
                           bht_28_11_port);
   bht_reg_30_11_inst : DLH_X1 port map( G => N2164, D => N3755, Q => 
                           bht_30_11_port);
   bht_reg_31_11_inst : DLH_X1 port map( G => N2110, D => N3755, Q => 
                           bht_31_11_port);
   bht_reg_29_11_inst : DLH_X1 port map( G => N2218, D => N3755, Q => 
                           bht_29_11_port);
   bht_reg_27_11_inst : DLH_X1 port map( G => N2326, D => N3755, Q => 
                           bht_27_11_port);
   bht_reg_25_11_inst : DLH_X1 port map( G => N2434, D => N3755, Q => 
                           bht_25_11_port);
   bht_reg_23_11_inst : DLH_X1 port map( G => N2542, D => N3755, Q => 
                           bht_23_11_port);
   bht_reg_21_11_inst : DLH_X1 port map( G => N2650, D => N3755, Q => 
                           bht_21_11_port);
   bht_reg_19_11_inst : DLH_X1 port map( G => N2758, D => N3755, Q => 
                           bht_19_11_port);
   bht_reg_17_11_inst : DLH_X1 port map( G => N2866, D => N3755, Q => 
                           bht_17_11_port);
   bht_reg_15_11_inst : DLH_X1 port map( G => N2974, D => N3755, Q => 
                           bht_15_11_port);
   bht_reg_13_11_inst : DLH_X1 port map( G => N3082, D => N3755, Q => 
                           bht_13_11_port);
   bht_reg_11_11_inst : DLH_X1 port map( G => N3190, D => N3755, Q => 
                           bht_11_11_port);
   bht_reg_9_11_inst : DLH_X1 port map( G => N3298, D => N3755, Q => 
                           bht_9_11_port);
   bht_reg_7_11_inst : DLH_X1 port map( G => N3406, D => N3755, Q => 
                           bht_7_11_port);
   bht_reg_5_11_inst : DLH_X1 port map( G => N3514, D => N3755, Q => 
                           bht_5_11_port);
   bht_reg_3_11_inst : DLH_X1 port map( G => N3622, D => N3755, Q => 
                           bht_3_11_port);
   bht_reg_1_11_inst : DLH_X1 port map( G => N3730, D => N3755, Q => 
                           bht_1_11_port);
   entry_r_reg_10_inst : DLH_X1 port map( G => N188, D => N135, Q => 
                           entry_r_10_port);
   entry_r_delay_reg_10_inst : DFFR_X1 port map( D => entry_r_10_port, CK => 
                           clk, RN => rst, Q => net108075, QN => n18);
   bht_reg_0_10_inst : DLH_X1 port map( G => N3784, D => N3753, Q => 
                           bht_0_10_port);
   bht_reg_2_10_inst : DLH_X1 port map( G => N3676, D => N3753, Q => 
                           bht_2_10_port);
   bht_reg_4_10_inst : DLH_X1 port map( G => N3568, D => N3753, Q => 
                           bht_4_10_port);
   bht_reg_6_10_inst : DLH_X1 port map( G => N3460, D => N3753, Q => 
                           bht_6_10_port);
   bht_reg_8_10_inst : DLH_X1 port map( G => N3352, D => N3753, Q => 
                           bht_8_10_port);
   bht_reg_10_10_inst : DLH_X1 port map( G => N3244, D => N3753, Q => 
                           bht_10_10_port);
   bht_reg_12_10_inst : DLH_X1 port map( G => N3136, D => N3753, Q => 
                           bht_12_10_port);
   bht_reg_14_10_inst : DLH_X1 port map( G => N3028, D => N3753, Q => 
                           bht_14_10_port);
   bht_reg_16_10_inst : DLH_X1 port map( G => N2920, D => N3753, Q => 
                           bht_16_10_port);
   bht_reg_18_10_inst : DLH_X1 port map( G => N2812, D => N3753, Q => 
                           bht_18_10_port);
   bht_reg_20_10_inst : DLH_X1 port map( G => N2704, D => N3753, Q => 
                           bht_20_10_port);
   bht_reg_22_10_inst : DLH_X1 port map( G => N2596, D => N3753, Q => 
                           bht_22_10_port);
   bht_reg_24_10_inst : DLH_X1 port map( G => N2488, D => N3753, Q => 
                           bht_24_10_port);
   bht_reg_26_10_inst : DLH_X1 port map( G => N2380, D => N3753, Q => 
                           bht_26_10_port);
   bht_reg_28_10_inst : DLH_X1 port map( G => N2272, D => N3753, Q => 
                           bht_28_10_port);
   bht_reg_30_10_inst : DLH_X1 port map( G => N2164, D => N3753, Q => 
                           bht_30_10_port);
   bht_reg_31_10_inst : DLH_X1 port map( G => N2110, D => N3753, Q => 
                           bht_31_10_port);
   bht_reg_29_10_inst : DLH_X1 port map( G => N2218, D => N3753, Q => 
                           bht_29_10_port);
   bht_reg_27_10_inst : DLH_X1 port map( G => N2326, D => N3753, Q => 
                           bht_27_10_port);
   bht_reg_25_10_inst : DLH_X1 port map( G => N2434, D => N3753, Q => 
                           bht_25_10_port);
   bht_reg_23_10_inst : DLH_X1 port map( G => N2542, D => N3753, Q => 
                           bht_23_10_port);
   bht_reg_21_10_inst : DLH_X1 port map( G => N2650, D => N3753, Q => 
                           bht_21_10_port);
   bht_reg_19_10_inst : DLH_X1 port map( G => N2758, D => N3753, Q => 
                           bht_19_10_port);
   bht_reg_17_10_inst : DLH_X1 port map( G => N2866, D => N3753, Q => 
                           bht_17_10_port);
   bht_reg_15_10_inst : DLH_X1 port map( G => N2974, D => N3753, Q => 
                           bht_15_10_port);
   bht_reg_13_10_inst : DLH_X1 port map( G => N3082, D => N3753, Q => 
                           bht_13_10_port);
   bht_reg_11_10_inst : DLH_X1 port map( G => N3190, D => N3753, Q => 
                           bht_11_10_port);
   bht_reg_9_10_inst : DLH_X1 port map( G => N3298, D => N3753, Q => 
                           bht_9_10_port);
   bht_reg_7_10_inst : DLH_X1 port map( G => N3406, D => N3753, Q => 
                           bht_7_10_port);
   bht_reg_5_10_inst : DLH_X1 port map( G => N3514, D => N3753, Q => 
                           bht_5_10_port);
   bht_reg_3_10_inst : DLH_X1 port map( G => N3622, D => N3753, Q => 
                           bht_3_10_port);
   bht_reg_1_10_inst : DLH_X1 port map( G => N3730, D => N3753, Q => 
                           bht_1_10_port);
   entry_r_reg_9_inst : DLH_X1 port map( G => N188, D => N134, Q => 
                           entry_r_9_port);
   entry_r_delay_reg_9_inst : DFFR_X1 port map( D => entry_r_9_port, CK => clk,
                           RN => rst, Q => net108074, QN => n17);
   bht_reg_0_9_inst : DLH_X1 port map( G => N3784, D => N3751, Q => 
                           bht_0_9_port);
   bht_reg_2_9_inst : DLH_X1 port map( G => N3676, D => N3751, Q => 
                           bht_2_9_port);
   bht_reg_4_9_inst : DLH_X1 port map( G => N3568, D => N3751, Q => 
                           bht_4_9_port);
   bht_reg_6_9_inst : DLH_X1 port map( G => N3460, D => N3751, Q => 
                           bht_6_9_port);
   bht_reg_8_9_inst : DLH_X1 port map( G => N3352, D => N3751, Q => 
                           bht_8_9_port);
   bht_reg_10_9_inst : DLH_X1 port map( G => N3244, D => N3751, Q => 
                           bht_10_9_port);
   bht_reg_12_9_inst : DLH_X1 port map( G => N3136, D => N3751, Q => 
                           bht_12_9_port);
   bht_reg_14_9_inst : DLH_X1 port map( G => N3028, D => N3751, Q => 
                           bht_14_9_port);
   bht_reg_16_9_inst : DLH_X1 port map( G => N2920, D => N3751, Q => 
                           bht_16_9_port);
   bht_reg_18_9_inst : DLH_X1 port map( G => N2812, D => N3751, Q => 
                           bht_18_9_port);
   bht_reg_20_9_inst : DLH_X1 port map( G => N2704, D => N3751, Q => 
                           bht_20_9_port);
   bht_reg_22_9_inst : DLH_X1 port map( G => N2596, D => N3751, Q => 
                           bht_22_9_port);
   bht_reg_24_9_inst : DLH_X1 port map( G => N2488, D => N3751, Q => 
                           bht_24_9_port);
   bht_reg_26_9_inst : DLH_X1 port map( G => N2380, D => N3751, Q => 
                           bht_26_9_port);
   bht_reg_28_9_inst : DLH_X1 port map( G => N2272, D => N3751, Q => 
                           bht_28_9_port);
   bht_reg_30_9_inst : DLH_X1 port map( G => N2164, D => N3751, Q => 
                           bht_30_9_port);
   bht_reg_31_9_inst : DLH_X1 port map( G => N2110, D => N3751, Q => 
                           bht_31_9_port);
   bht_reg_29_9_inst : DLH_X1 port map( G => N2218, D => N3751, Q => 
                           bht_29_9_port);
   bht_reg_27_9_inst : DLH_X1 port map( G => N2326, D => N3751, Q => 
                           bht_27_9_port);
   bht_reg_25_9_inst : DLH_X1 port map( G => N2434, D => N3751, Q => 
                           bht_25_9_port);
   bht_reg_23_9_inst : DLH_X1 port map( G => N2542, D => N3751, Q => 
                           bht_23_9_port);
   bht_reg_21_9_inst : DLH_X1 port map( G => N2650, D => N3751, Q => 
                           bht_21_9_port);
   bht_reg_19_9_inst : DLH_X1 port map( G => N2758, D => N3751, Q => 
                           bht_19_9_port);
   bht_reg_17_9_inst : DLH_X1 port map( G => N2866, D => N3751, Q => 
                           bht_17_9_port);
   bht_reg_15_9_inst : DLH_X1 port map( G => N2974, D => N3751, Q => 
                           bht_15_9_port);
   bht_reg_13_9_inst : DLH_X1 port map( G => N3082, D => N3751, Q => 
                           bht_13_9_port);
   bht_reg_11_9_inst : DLH_X1 port map( G => N3190, D => N3751, Q => 
                           bht_11_9_port);
   bht_reg_9_9_inst : DLH_X1 port map( G => N3298, D => N3751, Q => 
                           bht_9_9_port);
   bht_reg_7_9_inst : DLH_X1 port map( G => N3406, D => N3751, Q => 
                           bht_7_9_port);
   bht_reg_5_9_inst : DLH_X1 port map( G => N3514, D => N3751, Q => 
                           bht_5_9_port);
   bht_reg_3_9_inst : DLH_X1 port map( G => N3622, D => N3751, Q => 
                           bht_3_9_port);
   bht_reg_1_9_inst : DLH_X1 port map( G => N3730, D => N3751, Q => 
                           bht_1_9_port);
   entry_r_reg_8_inst : DLH_X1 port map( G => N188, D => N133, Q => 
                           entry_r_8_port);
   entry_r_delay_reg_8_inst : DFFR_X1 port map( D => entry_r_8_port, CK => clk,
                           RN => rst, Q => net108073, QN => n16);
   bht_reg_0_8_inst : DLH_X1 port map( G => N3784, D => N3749, Q => 
                           bht_0_8_port);
   bht_reg_2_8_inst : DLH_X1 port map( G => N3676, D => N3749, Q => 
                           bht_2_8_port);
   bht_reg_4_8_inst : DLH_X1 port map( G => N3568, D => N3749, Q => 
                           bht_4_8_port);
   bht_reg_6_8_inst : DLH_X1 port map( G => N3460, D => N3749, Q => 
                           bht_6_8_port);
   bht_reg_8_8_inst : DLH_X1 port map( G => N3352, D => N3749, Q => 
                           bht_8_8_port);
   bht_reg_10_8_inst : DLH_X1 port map( G => N3244, D => N3749, Q => 
                           bht_10_8_port);
   bht_reg_12_8_inst : DLH_X1 port map( G => N3136, D => N3749, Q => 
                           bht_12_8_port);
   bht_reg_14_8_inst : DLH_X1 port map( G => N3028, D => N3749, Q => 
                           bht_14_8_port);
   bht_reg_16_8_inst : DLH_X1 port map( G => N2920, D => N3749, Q => 
                           bht_16_8_port);
   bht_reg_18_8_inst : DLH_X1 port map( G => N2812, D => N3749, Q => 
                           bht_18_8_port);
   bht_reg_20_8_inst : DLH_X1 port map( G => N2704, D => N3749, Q => 
                           bht_20_8_port);
   bht_reg_22_8_inst : DLH_X1 port map( G => N2596, D => N3749, Q => 
                           bht_22_8_port);
   bht_reg_24_8_inst : DLH_X1 port map( G => N2488, D => N3749, Q => 
                           bht_24_8_port);
   bht_reg_26_8_inst : DLH_X1 port map( G => N2380, D => N3749, Q => 
                           bht_26_8_port);
   bht_reg_28_8_inst : DLH_X1 port map( G => N2272, D => N3749, Q => 
                           bht_28_8_port);
   bht_reg_30_8_inst : DLH_X1 port map( G => N2164, D => N3749, Q => 
                           bht_30_8_port);
   bht_reg_31_8_inst : DLH_X1 port map( G => N2110, D => N3749, Q => 
                           bht_31_8_port);
   bht_reg_29_8_inst : DLH_X1 port map( G => N2218, D => N3749, Q => 
                           bht_29_8_port);
   bht_reg_27_8_inst : DLH_X1 port map( G => N2326, D => N3749, Q => 
                           bht_27_8_port);
   bht_reg_25_8_inst : DLH_X1 port map( G => N2434, D => N3749, Q => 
                           bht_25_8_port);
   bht_reg_23_8_inst : DLH_X1 port map( G => N2542, D => N3749, Q => 
                           bht_23_8_port);
   bht_reg_21_8_inst : DLH_X1 port map( G => N2650, D => N3749, Q => 
                           bht_21_8_port);
   bht_reg_19_8_inst : DLH_X1 port map( G => N2758, D => N3749, Q => 
                           bht_19_8_port);
   bht_reg_17_8_inst : DLH_X1 port map( G => N2866, D => N3749, Q => 
                           bht_17_8_port);
   bht_reg_15_8_inst : DLH_X1 port map( G => N2974, D => N3749, Q => 
                           bht_15_8_port);
   bht_reg_13_8_inst : DLH_X1 port map( G => N3082, D => N3749, Q => 
                           bht_13_8_port);
   bht_reg_11_8_inst : DLH_X1 port map( G => N3190, D => N3749, Q => 
                           bht_11_8_port);
   bht_reg_9_8_inst : DLH_X1 port map( G => N3298, D => N3749, Q => 
                           bht_9_8_port);
   bht_reg_7_8_inst : DLH_X1 port map( G => N3406, D => N3749, Q => 
                           bht_7_8_port);
   bht_reg_5_8_inst : DLH_X1 port map( G => N3514, D => N3749, Q => 
                           bht_5_8_port);
   bht_reg_3_8_inst : DLH_X1 port map( G => N3622, D => N3749, Q => 
                           bht_3_8_port);
   bht_reg_1_8_inst : DLH_X1 port map( G => N3730, D => N3749, Q => 
                           bht_1_8_port);
   entry_r_reg_7_inst : DLH_X1 port map( G => N188, D => N132, Q => 
                           entry_r_7_port);
   entry_r_delay_reg_7_inst : DFFR_X1 port map( D => entry_r_7_port, CK => clk,
                           RN => rst, Q => net108072, QN => n15);
   bht_reg_0_7_inst : DLH_X1 port map( G => N3784, D => N3747, Q => 
                           bht_0_7_port);
   bht_reg_2_7_inst : DLH_X1 port map( G => N3676, D => N3747, Q => 
                           bht_2_7_port);
   bht_reg_4_7_inst : DLH_X1 port map( G => N3568, D => N3747, Q => 
                           bht_4_7_port);
   bht_reg_6_7_inst : DLH_X1 port map( G => N3460, D => N3747, Q => 
                           bht_6_7_port);
   bht_reg_8_7_inst : DLH_X1 port map( G => N3352, D => N3747, Q => 
                           bht_8_7_port);
   bht_reg_10_7_inst : DLH_X1 port map( G => N3244, D => N3747, Q => 
                           bht_10_7_port);
   bht_reg_12_7_inst : DLH_X1 port map( G => N3136, D => N3747, Q => 
                           bht_12_7_port);
   bht_reg_14_7_inst : DLH_X1 port map( G => N3028, D => N3747, Q => 
                           bht_14_7_port);
   bht_reg_16_7_inst : DLH_X1 port map( G => N2920, D => N3747, Q => 
                           bht_16_7_port);
   bht_reg_18_7_inst : DLH_X1 port map( G => N2812, D => N3747, Q => 
                           bht_18_7_port);
   bht_reg_20_7_inst : DLH_X1 port map( G => N2704, D => N3747, Q => 
                           bht_20_7_port);
   bht_reg_22_7_inst : DLH_X1 port map( G => N2596, D => N3747, Q => 
                           bht_22_7_port);
   bht_reg_24_7_inst : DLH_X1 port map( G => N2488, D => N3747, Q => 
                           bht_24_7_port);
   bht_reg_26_7_inst : DLH_X1 port map( G => N2380, D => N3747, Q => 
                           bht_26_7_port);
   bht_reg_28_7_inst : DLH_X1 port map( G => N2272, D => N3747, Q => 
                           bht_28_7_port);
   bht_reg_30_7_inst : DLH_X1 port map( G => N2164, D => N3747, Q => 
                           bht_30_7_port);
   bht_reg_31_7_inst : DLH_X1 port map( G => N2110, D => N3747, Q => 
                           bht_31_7_port);
   bht_reg_29_7_inst : DLH_X1 port map( G => N2218, D => N3747, Q => 
                           bht_29_7_port);
   bht_reg_27_7_inst : DLH_X1 port map( G => N2326, D => N3747, Q => 
                           bht_27_7_port);
   bht_reg_25_7_inst : DLH_X1 port map( G => N2434, D => N3747, Q => 
                           bht_25_7_port);
   bht_reg_23_7_inst : DLH_X1 port map( G => N2542, D => N3747, Q => 
                           bht_23_7_port);
   bht_reg_21_7_inst : DLH_X1 port map( G => N2650, D => N3747, Q => 
                           bht_21_7_port);
   bht_reg_19_7_inst : DLH_X1 port map( G => N2758, D => N3747, Q => 
                           bht_19_7_port);
   bht_reg_17_7_inst : DLH_X1 port map( G => N2866, D => N3747, Q => 
                           bht_17_7_port);
   bht_reg_15_7_inst : DLH_X1 port map( G => N2974, D => N3747, Q => 
                           bht_15_7_port);
   bht_reg_13_7_inst : DLH_X1 port map( G => N3082, D => N3747, Q => 
                           bht_13_7_port);
   bht_reg_11_7_inst : DLH_X1 port map( G => N3190, D => N3747, Q => 
                           bht_11_7_port);
   bht_reg_9_7_inst : DLH_X1 port map( G => N3298, D => N3747, Q => 
                           bht_9_7_port);
   bht_reg_7_7_inst : DLH_X1 port map( G => N3406, D => N3747, Q => 
                           bht_7_7_port);
   bht_reg_5_7_inst : DLH_X1 port map( G => N3514, D => N3747, Q => 
                           bht_5_7_port);
   bht_reg_3_7_inst : DLH_X1 port map( G => N3622, D => N3747, Q => 
                           bht_3_7_port);
   bht_reg_1_7_inst : DLH_X1 port map( G => N3730, D => N3747, Q => 
                           bht_1_7_port);
   entry_r_reg_6_inst : DLH_X1 port map( G => N188, D => N131, Q => 
                           entry_r_6_port);
   entry_r_delay_reg_6_inst : DFFR_X1 port map( D => entry_r_6_port, CK => clk,
                           RN => rst, Q => net108071, QN => n14);
   bht_reg_0_6_inst : DLH_X1 port map( G => N3784, D => N3745, Q => 
                           bht_0_6_port);
   bht_reg_2_6_inst : DLH_X1 port map( G => N3676, D => N3745, Q => 
                           bht_2_6_port);
   bht_reg_4_6_inst : DLH_X1 port map( G => N3568, D => N3745, Q => 
                           bht_4_6_port);
   bht_reg_6_6_inst : DLH_X1 port map( G => N3460, D => N3745, Q => 
                           bht_6_6_port);
   bht_reg_8_6_inst : DLH_X1 port map( G => N3352, D => N3745, Q => 
                           bht_8_6_port);
   bht_reg_10_6_inst : DLH_X1 port map( G => N3244, D => N3745, Q => 
                           bht_10_6_port);
   bht_reg_12_6_inst : DLH_X1 port map( G => N3136, D => N3745, Q => 
                           bht_12_6_port);
   bht_reg_14_6_inst : DLH_X1 port map( G => N3028, D => N3745, Q => 
                           bht_14_6_port);
   bht_reg_16_6_inst : DLH_X1 port map( G => N2920, D => N3745, Q => 
                           bht_16_6_port);
   bht_reg_18_6_inst : DLH_X1 port map( G => N2812, D => N3745, Q => 
                           bht_18_6_port);
   bht_reg_20_6_inst : DLH_X1 port map( G => N2704, D => N3745, Q => 
                           bht_20_6_port);
   bht_reg_22_6_inst : DLH_X1 port map( G => N2596, D => N3745, Q => 
                           bht_22_6_port);
   bht_reg_24_6_inst : DLH_X1 port map( G => N2488, D => N3745, Q => 
                           bht_24_6_port);
   bht_reg_26_6_inst : DLH_X1 port map( G => N2380, D => N3745, Q => 
                           bht_26_6_port);
   bht_reg_28_6_inst : DLH_X1 port map( G => N2272, D => N3745, Q => 
                           bht_28_6_port);
   bht_reg_30_6_inst : DLH_X1 port map( G => N2164, D => N3745, Q => 
                           bht_30_6_port);
   bht_reg_31_6_inst : DLH_X1 port map( G => N2110, D => N3745, Q => 
                           bht_31_6_port);
   bht_reg_29_6_inst : DLH_X1 port map( G => N2218, D => N3745, Q => 
                           bht_29_6_port);
   bht_reg_27_6_inst : DLH_X1 port map( G => N2326, D => N3745, Q => 
                           bht_27_6_port);
   bht_reg_25_6_inst : DLH_X1 port map( G => N2434, D => N3745, Q => 
                           bht_25_6_port);
   bht_reg_23_6_inst : DLH_X1 port map( G => N2542, D => N3745, Q => 
                           bht_23_6_port);
   bht_reg_21_6_inst : DLH_X1 port map( G => N2650, D => N3745, Q => 
                           bht_21_6_port);
   bht_reg_19_6_inst : DLH_X1 port map( G => N2758, D => N3745, Q => 
                           bht_19_6_port);
   bht_reg_17_6_inst : DLH_X1 port map( G => N2866, D => N3745, Q => 
                           bht_17_6_port);
   bht_reg_15_6_inst : DLH_X1 port map( G => N2974, D => N3745, Q => 
                           bht_15_6_port);
   bht_reg_13_6_inst : DLH_X1 port map( G => N3082, D => N3745, Q => 
                           bht_13_6_port);
   bht_reg_11_6_inst : DLH_X1 port map( G => N3190, D => N3745, Q => 
                           bht_11_6_port);
   bht_reg_9_6_inst : DLH_X1 port map( G => N3298, D => N3745, Q => 
                           bht_9_6_port);
   bht_reg_7_6_inst : DLH_X1 port map( G => N3406, D => N3745, Q => 
                           bht_7_6_port);
   bht_reg_5_6_inst : DLH_X1 port map( G => N3514, D => N3745, Q => 
                           bht_5_6_port);
   bht_reg_3_6_inst : DLH_X1 port map( G => N3622, D => N3745, Q => 
                           bht_3_6_port);
   bht_reg_1_6_inst : DLH_X1 port map( G => N3730, D => N3745, Q => 
                           bht_1_6_port);
   entry_r_reg_5_inst : DLH_X1 port map( G => N188, D => N130, Q => 
                           entry_r_5_port);
   entry_r_delay_reg_5_inst : DFFR_X1 port map( D => entry_r_5_port, CK => clk,
                           RN => rst, Q => net108070, QN => n13);
   bht_reg_0_5_inst : DLH_X1 port map( G => N3784, D => N3743, Q => 
                           bht_0_5_port);
   bht_reg_2_5_inst : DLH_X1 port map( G => N3676, D => N3743, Q => 
                           bht_2_5_port);
   bht_reg_4_5_inst : DLH_X1 port map( G => N3568, D => N3743, Q => 
                           bht_4_5_port);
   bht_reg_6_5_inst : DLH_X1 port map( G => N3460, D => N3743, Q => 
                           bht_6_5_port);
   bht_reg_8_5_inst : DLH_X1 port map( G => N3352, D => N3743, Q => 
                           bht_8_5_port);
   bht_reg_10_5_inst : DLH_X1 port map( G => N3244, D => N3743, Q => 
                           bht_10_5_port);
   bht_reg_12_5_inst : DLH_X1 port map( G => N3136, D => N3743, Q => 
                           bht_12_5_port);
   bht_reg_14_5_inst : DLH_X1 port map( G => N3028, D => N3743, Q => 
                           bht_14_5_port);
   bht_reg_16_5_inst : DLH_X1 port map( G => N2920, D => N3743, Q => 
                           bht_16_5_port);
   bht_reg_18_5_inst : DLH_X1 port map( G => N2812, D => N3743, Q => 
                           bht_18_5_port);
   bht_reg_20_5_inst : DLH_X1 port map( G => N2704, D => N3743, Q => 
                           bht_20_5_port);
   bht_reg_22_5_inst : DLH_X1 port map( G => N2596, D => N3743, Q => 
                           bht_22_5_port);
   bht_reg_24_5_inst : DLH_X1 port map( G => N2488, D => N3743, Q => 
                           bht_24_5_port);
   bht_reg_26_5_inst : DLH_X1 port map( G => N2380, D => N3743, Q => 
                           bht_26_5_port);
   bht_reg_28_5_inst : DLH_X1 port map( G => N2272, D => N3743, Q => 
                           bht_28_5_port);
   bht_reg_30_5_inst : DLH_X1 port map( G => N2164, D => N3743, Q => 
                           bht_30_5_port);
   bht_reg_31_5_inst : DLH_X1 port map( G => N2110, D => N3743, Q => 
                           bht_31_5_port);
   bht_reg_29_5_inst : DLH_X1 port map( G => N2218, D => N3743, Q => 
                           bht_29_5_port);
   bht_reg_27_5_inst : DLH_X1 port map( G => N2326, D => N3743, Q => 
                           bht_27_5_port);
   bht_reg_25_5_inst : DLH_X1 port map( G => N2434, D => N3743, Q => 
                           bht_25_5_port);
   bht_reg_23_5_inst : DLH_X1 port map( G => N2542, D => N3743, Q => 
                           bht_23_5_port);
   bht_reg_21_5_inst : DLH_X1 port map( G => N2650, D => N3743, Q => 
                           bht_21_5_port);
   bht_reg_19_5_inst : DLH_X1 port map( G => N2758, D => N3743, Q => 
                           bht_19_5_port);
   bht_reg_17_5_inst : DLH_X1 port map( G => N2866, D => N3743, Q => 
                           bht_17_5_port);
   bht_reg_15_5_inst : DLH_X1 port map( G => N2974, D => N3743, Q => 
                           bht_15_5_port);
   bht_reg_13_5_inst : DLH_X1 port map( G => N3082, D => N3743, Q => 
                           bht_13_5_port);
   bht_reg_11_5_inst : DLH_X1 port map( G => N3190, D => N3743, Q => 
                           bht_11_5_port);
   bht_reg_9_5_inst : DLH_X1 port map( G => N3298, D => N3743, Q => 
                           bht_9_5_port);
   bht_reg_7_5_inst : DLH_X1 port map( G => N3406, D => N3743, Q => 
                           bht_7_5_port);
   bht_reg_5_5_inst : DLH_X1 port map( G => N3514, D => N3743, Q => 
                           bht_5_5_port);
   bht_reg_3_5_inst : DLH_X1 port map( G => N3622, D => N3743, Q => 
                           bht_3_5_port);
   bht_reg_1_5_inst : DLH_X1 port map( G => N3730, D => N3743, Q => 
                           bht_1_5_port);
   entry_r_reg_4_inst : DLH_X1 port map( G => N188, D => N129, Q => 
                           entry_r_4_port);
   entry_r_delay_reg_4_inst : DFFR_X1 port map( D => entry_r_4_port, CK => clk,
                           RN => rst, Q => net108069, QN => n12);
   bht_reg_0_4_inst : DLH_X1 port map( G => N3784, D => N3741, Q => 
                           bht_0_4_port);
   bht_reg_2_4_inst : DLH_X1 port map( G => N3676, D => N3741, Q => 
                           bht_2_4_port);
   bht_reg_4_4_inst : DLH_X1 port map( G => N3568, D => N3741, Q => 
                           bht_4_4_port);
   bht_reg_6_4_inst : DLH_X1 port map( G => N3460, D => N3741, Q => 
                           bht_6_4_port);
   bht_reg_8_4_inst : DLH_X1 port map( G => N3352, D => N3741, Q => 
                           bht_8_4_port);
   bht_reg_10_4_inst : DLH_X1 port map( G => N3244, D => N3741, Q => 
                           bht_10_4_port);
   bht_reg_12_4_inst : DLH_X1 port map( G => N3136, D => N3741, Q => 
                           bht_12_4_port);
   bht_reg_14_4_inst : DLH_X1 port map( G => N3028, D => N3741, Q => 
                           bht_14_4_port);
   bht_reg_16_4_inst : DLH_X1 port map( G => N2920, D => N3741, Q => 
                           bht_16_4_port);
   bht_reg_18_4_inst : DLH_X1 port map( G => N2812, D => N3741, Q => 
                           bht_18_4_port);
   bht_reg_20_4_inst : DLH_X1 port map( G => N2704, D => N3741, Q => 
                           bht_20_4_port);
   bht_reg_22_4_inst : DLH_X1 port map( G => N2596, D => N3741, Q => 
                           bht_22_4_port);
   bht_reg_24_4_inst : DLH_X1 port map( G => N2488, D => N3741, Q => 
                           bht_24_4_port);
   bht_reg_26_4_inst : DLH_X1 port map( G => N2380, D => N3741, Q => 
                           bht_26_4_port);
   bht_reg_28_4_inst : DLH_X1 port map( G => N2272, D => N3741, Q => 
                           bht_28_4_port);
   bht_reg_30_4_inst : DLH_X1 port map( G => N2164, D => N3741, Q => 
                           bht_30_4_port);
   bht_reg_31_4_inst : DLH_X1 port map( G => N2110, D => N3741, Q => 
                           bht_31_4_port);
   bht_reg_29_4_inst : DLH_X1 port map( G => N2218, D => N3741, Q => 
                           bht_29_4_port);
   bht_reg_27_4_inst : DLH_X1 port map( G => N2326, D => N3741, Q => 
                           bht_27_4_port);
   bht_reg_25_4_inst : DLH_X1 port map( G => N2434, D => N3741, Q => 
                           bht_25_4_port);
   bht_reg_23_4_inst : DLH_X1 port map( G => N2542, D => N3741, Q => 
                           bht_23_4_port);
   bht_reg_21_4_inst : DLH_X1 port map( G => N2650, D => N3741, Q => 
                           bht_21_4_port);
   bht_reg_19_4_inst : DLH_X1 port map( G => N2758, D => N3741, Q => 
                           bht_19_4_port);
   bht_reg_17_4_inst : DLH_X1 port map( G => N2866, D => N3741, Q => 
                           bht_17_4_port);
   bht_reg_15_4_inst : DLH_X1 port map( G => N2974, D => N3741, Q => 
                           bht_15_4_port);
   bht_reg_13_4_inst : DLH_X1 port map( G => N3082, D => N3741, Q => 
                           bht_13_4_port);
   bht_reg_11_4_inst : DLH_X1 port map( G => N3190, D => N3741, Q => 
                           bht_11_4_port);
   bht_reg_9_4_inst : DLH_X1 port map( G => N3298, D => N3741, Q => 
                           bht_9_4_port);
   bht_reg_7_4_inst : DLH_X1 port map( G => N3406, D => N3741, Q => 
                           bht_7_4_port);
   bht_reg_5_4_inst : DLH_X1 port map( G => N3514, D => N3741, Q => 
                           bht_5_4_port);
   bht_reg_3_4_inst : DLH_X1 port map( G => N3622, D => N3741, Q => 
                           bht_3_4_port);
   bht_reg_1_4_inst : DLH_X1 port map( G => N3730, D => N3741, Q => 
                           bht_1_4_port);
   entry_r_reg_3_inst : DLH_X1 port map( G => N188, D => N128, Q => 
                           entry_r_3_port);
   entry_r_delay_reg_3_inst : DFFR_X1 port map( D => entry_r_3_port, CK => clk,
                           RN => rst, Q => net108068, QN => n11);
   bht_reg_0_3_inst : DLH_X1 port map( G => N3784, D => N3739, Q => 
                           bht_0_3_port);
   bht_reg_2_3_inst : DLH_X1 port map( G => N3676, D => N3739, Q => 
                           bht_2_3_port);
   bht_reg_4_3_inst : DLH_X1 port map( G => N3568, D => N3739, Q => 
                           bht_4_3_port);
   bht_reg_6_3_inst : DLH_X1 port map( G => N3460, D => N3739, Q => 
                           bht_6_3_port);
   bht_reg_8_3_inst : DLH_X1 port map( G => N3352, D => N3739, Q => 
                           bht_8_3_port);
   bht_reg_10_3_inst : DLH_X1 port map( G => N3244, D => N3739, Q => 
                           bht_10_3_port);
   bht_reg_12_3_inst : DLH_X1 port map( G => N3136, D => N3739, Q => 
                           bht_12_3_port);
   bht_reg_14_3_inst : DLH_X1 port map( G => N3028, D => N3739, Q => 
                           bht_14_3_port);
   bht_reg_16_3_inst : DLH_X1 port map( G => N2920, D => N3739, Q => 
                           bht_16_3_port);
   bht_reg_18_3_inst : DLH_X1 port map( G => N2812, D => N3739, Q => 
                           bht_18_3_port);
   bht_reg_20_3_inst : DLH_X1 port map( G => N2704, D => N3739, Q => 
                           bht_20_3_port);
   bht_reg_22_3_inst : DLH_X1 port map( G => N2596, D => N3739, Q => 
                           bht_22_3_port);
   bht_reg_24_3_inst : DLH_X1 port map( G => N2488, D => N3739, Q => 
                           bht_24_3_port);
   bht_reg_26_3_inst : DLH_X1 port map( G => N2380, D => N3739, Q => 
                           bht_26_3_port);
   bht_reg_28_3_inst : DLH_X1 port map( G => N2272, D => N3739, Q => 
                           bht_28_3_port);
   bht_reg_30_3_inst : DLH_X1 port map( G => N2164, D => N3739, Q => 
                           bht_30_3_port);
   bht_reg_31_3_inst : DLH_X1 port map( G => N2110, D => N3739, Q => 
                           bht_31_3_port);
   bht_reg_29_3_inst : DLH_X1 port map( G => N2218, D => N3739, Q => 
                           bht_29_3_port);
   bht_reg_27_3_inst : DLH_X1 port map( G => N2326, D => N3739, Q => 
                           bht_27_3_port);
   bht_reg_25_3_inst : DLH_X1 port map( G => N2434, D => N3739, Q => 
                           bht_25_3_port);
   bht_reg_23_3_inst : DLH_X1 port map( G => N2542, D => N3739, Q => 
                           bht_23_3_port);
   bht_reg_21_3_inst : DLH_X1 port map( G => N2650, D => N3739, Q => 
                           bht_21_3_port);
   bht_reg_19_3_inst : DLH_X1 port map( G => N2758, D => N3739, Q => 
                           bht_19_3_port);
   bht_reg_17_3_inst : DLH_X1 port map( G => N2866, D => N3739, Q => 
                           bht_17_3_port);
   bht_reg_15_3_inst : DLH_X1 port map( G => N2974, D => N3739, Q => 
                           bht_15_3_port);
   bht_reg_13_3_inst : DLH_X1 port map( G => N3082, D => N3739, Q => 
                           bht_13_3_port);
   bht_reg_11_3_inst : DLH_X1 port map( G => N3190, D => N3739, Q => 
                           bht_11_3_port);
   bht_reg_9_3_inst : DLH_X1 port map( G => N3298, D => N3739, Q => 
                           bht_9_3_port);
   bht_reg_7_3_inst : DLH_X1 port map( G => N3406, D => N3739, Q => 
                           bht_7_3_port);
   bht_reg_5_3_inst : DLH_X1 port map( G => N3514, D => N3739, Q => 
                           bht_5_3_port);
   bht_reg_3_3_inst : DLH_X1 port map( G => N3622, D => N3739, Q => 
                           bht_3_3_port);
   bht_reg_1_3_inst : DLH_X1 port map( G => N3730, D => N3739, Q => 
                           bht_1_3_port);
   entry_r_reg_2_inst : DLH_X1 port map( G => N188, D => N127, Q => 
                           entry_r_2_port);
   entry_r_delay_reg_2_inst : DFFR_X1 port map( D => entry_r_2_port, CK => clk,
                           RN => rst, Q => net108067, QN => n10);
   bht_reg_0_2_inst : DLH_X1 port map( G => N3784, D => N3737, Q => 
                           bht_0_2_port);
   bht_reg_2_2_inst : DLH_X1 port map( G => N3676, D => N3737, Q => 
                           bht_2_2_port);
   bht_reg_4_2_inst : DLH_X1 port map( G => N3568, D => N3737, Q => 
                           bht_4_2_port);
   bht_reg_6_2_inst : DLH_X1 port map( G => N3460, D => N3737, Q => 
                           bht_6_2_port);
   bht_reg_8_2_inst : DLH_X1 port map( G => N3352, D => N3737, Q => 
                           bht_8_2_port);
   bht_reg_10_2_inst : DLH_X1 port map( G => N3244, D => N3737, Q => 
                           bht_10_2_port);
   bht_reg_12_2_inst : DLH_X1 port map( G => N3136, D => N3737, Q => 
                           bht_12_2_port);
   bht_reg_14_2_inst : DLH_X1 port map( G => N3028, D => N3737, Q => 
                           bht_14_2_port);
   bht_reg_16_2_inst : DLH_X1 port map( G => N2920, D => N3737, Q => 
                           bht_16_2_port);
   bht_reg_18_2_inst : DLH_X1 port map( G => N2812, D => N3737, Q => 
                           bht_18_2_port);
   bht_reg_20_2_inst : DLH_X1 port map( G => N2704, D => N3737, Q => 
                           bht_20_2_port);
   bht_reg_22_2_inst : DLH_X1 port map( G => N2596, D => N3737, Q => 
                           bht_22_2_port);
   bht_reg_24_2_inst : DLH_X1 port map( G => N2488, D => N3737, Q => 
                           bht_24_2_port);
   bht_reg_26_2_inst : DLH_X1 port map( G => N2380, D => N3737, Q => 
                           bht_26_2_port);
   bht_reg_28_2_inst : DLH_X1 port map( G => N2272, D => N3737, Q => 
                           bht_28_2_port);
   bht_reg_30_2_inst : DLH_X1 port map( G => N2164, D => N3737, Q => 
                           bht_30_2_port);
   bht_reg_31_2_inst : DLH_X1 port map( G => N2110, D => N3737, Q => 
                           bht_31_2_port);
   bht_reg_29_2_inst : DLH_X1 port map( G => N2218, D => N3737, Q => 
                           bht_29_2_port);
   bht_reg_27_2_inst : DLH_X1 port map( G => N2326, D => N3737, Q => 
                           bht_27_2_port);
   bht_reg_25_2_inst : DLH_X1 port map( G => N2434, D => N3737, Q => 
                           bht_25_2_port);
   bht_reg_23_2_inst : DLH_X1 port map( G => N2542, D => N3737, Q => 
                           bht_23_2_port);
   bht_reg_21_2_inst : DLH_X1 port map( G => N2650, D => N3737, Q => 
                           bht_21_2_port);
   bht_reg_19_2_inst : DLH_X1 port map( G => N2758, D => N3737, Q => 
                           bht_19_2_port);
   bht_reg_17_2_inst : DLH_X1 port map( G => N2866, D => N3737, Q => 
                           bht_17_2_port);
   bht_reg_15_2_inst : DLH_X1 port map( G => N2974, D => N3737, Q => 
                           bht_15_2_port);
   bht_reg_13_2_inst : DLH_X1 port map( G => N3082, D => N3737, Q => 
                           bht_13_2_port);
   bht_reg_11_2_inst : DLH_X1 port map( G => N3190, D => N3737, Q => 
                           bht_11_2_port);
   bht_reg_9_2_inst : DLH_X1 port map( G => N3298, D => N3737, Q => 
                           bht_9_2_port);
   bht_reg_7_2_inst : DLH_X1 port map( G => N3406, D => N3737, Q => 
                           bht_7_2_port);
   bht_reg_5_2_inst : DLH_X1 port map( G => N3514, D => N3737, Q => 
                           bht_5_2_port);
   bht_reg_3_2_inst : DLH_X1 port map( G => N3622, D => N3737, Q => 
                           bht_3_2_port);
   bht_reg_1_2_inst : DLH_X1 port map( G => N3730, D => N3737, Q => 
                           bht_1_2_port);
   sig_brt_delay_reg : DFFR_X1 port map( D => sig_brt_tmp, CK => clk, RN => rst
                           , Q => sig_brt_delay, QN => n7);
   bht_reg_0_0_inst : DLH_X1 port map( G => N3784, D => N3733, Q => 
                           bht_0_0_port);
   bht_reg_2_0_inst : DLH_X1 port map( G => N3676, D => N3733, Q => 
                           bht_2_0_port);
   bht_reg_4_0_inst : DLH_X1 port map( G => N3568, D => N3733, Q => 
                           bht_4_0_port);
   bht_reg_6_0_inst : DLH_X1 port map( G => N3460, D => N3733, Q => 
                           bht_6_0_port);
   bht_reg_8_0_inst : DLH_X1 port map( G => N3352, D => N3733, Q => 
                           bht_8_0_port);
   bht_reg_10_0_inst : DLH_X1 port map( G => N3244, D => N3733, Q => 
                           bht_10_0_port);
   bht_reg_12_0_inst : DLH_X1 port map( G => N3136, D => N3733, Q => 
                           bht_12_0_port);
   bht_reg_14_0_inst : DLH_X1 port map( G => N3028, D => N3733, Q => 
                           bht_14_0_port);
   bht_reg_16_0_inst : DLH_X1 port map( G => N2920, D => N3733, Q => 
                           bht_16_0_port);
   bht_reg_18_0_inst : DLH_X1 port map( G => N2812, D => N3733, Q => 
                           bht_18_0_port);
   bht_reg_20_0_inst : DLH_X1 port map( G => N2704, D => N3733, Q => 
                           bht_20_0_port);
   bht_reg_22_0_inst : DLH_X1 port map( G => N2596, D => N3733, Q => 
                           bht_22_0_port);
   bht_reg_24_0_inst : DLH_X1 port map( G => N2488, D => N3733, Q => 
                           bht_24_0_port);
   bht_reg_26_0_inst : DLH_X1 port map( G => N2380, D => N3733, Q => 
                           bht_26_0_port);
   bht_reg_28_0_inst : DLH_X1 port map( G => N2272, D => N3733, Q => 
                           bht_28_0_port);
   bht_reg_30_0_inst : DLH_X1 port map( G => N2164, D => N3733, Q => 
                           bht_30_0_port);
   bht_reg_31_0_inst : DLH_X1 port map( G => N2110, D => N3733, Q => 
                           bht_31_0_port);
   bht_reg_29_0_inst : DLH_X1 port map( G => N2218, D => N3733, Q => 
                           bht_29_0_port);
   bht_reg_27_0_inst : DLH_X1 port map( G => N2326, D => N3733, Q => 
                           bht_27_0_port);
   bht_reg_25_0_inst : DLH_X1 port map( G => N2434, D => N3733, Q => 
                           bht_25_0_port);
   bht_reg_23_0_inst : DLH_X1 port map( G => N2542, D => N3733, Q => 
                           bht_23_0_port);
   bht_reg_21_0_inst : DLH_X1 port map( G => N2650, D => N3733, Q => 
                           bht_21_0_port);
   bht_reg_19_0_inst : DLH_X1 port map( G => N2758, D => N3733, Q => 
                           bht_19_0_port);
   bht_reg_17_0_inst : DLH_X1 port map( G => N2866, D => N3733, Q => 
                           bht_17_0_port);
   bht_reg_15_0_inst : DLH_X1 port map( G => N2974, D => N3733, Q => 
                           bht_15_0_port);
   bht_reg_13_0_inst : DLH_X1 port map( G => N3082, D => N3733, Q => 
                           bht_13_0_port);
   bht_reg_11_0_inst : DLH_X1 port map( G => N3190, D => N3733, Q => 
                           bht_11_0_port);
   bht_reg_9_0_inst : DLH_X1 port map( G => N3298, D => N3733, Q => 
                           bht_9_0_port);
   bht_reg_7_0_inst : DLH_X1 port map( G => N3406, D => N3733, Q => 
                           bht_7_0_port);
   bht_reg_5_0_inst : DLH_X1 port map( G => N3514, D => N3733, Q => 
                           bht_5_0_port);
   bht_reg_3_0_inst : DLH_X1 port map( G => N3622, D => N3733, Q => 
                           bht_3_0_port);
   bht_reg_1_0_inst : DLH_X1 port map( G => N3730, D => N3733, Q => 
                           bht_1_0_port);
   entry_r_reg_0_inst : DLH_X1 port map( G => N188, D => N125, Q => 
                           entry_r_0_port);
   entry_r_delay_reg_0_inst : DFFR_X1 port map( D => entry_r_0_port, CK => clk,
                           RN => rst, Q => net108066, QN => n207);
   bht_reg_0_1_inst : DLH_X1 port map( G => N3784, D => N3735, Q => 
                           bht_0_1_port);
   bht_reg_2_1_inst : DLH_X1 port map( G => N3676, D => N3735, Q => 
                           bht_2_1_port);
   bht_reg_4_1_inst : DLH_X1 port map( G => N3568, D => N3735, Q => 
                           bht_4_1_port);
   bht_reg_6_1_inst : DLH_X1 port map( G => N3460, D => N3735, Q => 
                           bht_6_1_port);
   bht_reg_8_1_inst : DLH_X1 port map( G => N3352, D => N3735, Q => 
                           bht_8_1_port);
   bht_reg_10_1_inst : DLH_X1 port map( G => N3244, D => N3735, Q => 
                           bht_10_1_port);
   bht_reg_12_1_inst : DLH_X1 port map( G => N3136, D => N3735, Q => 
                           bht_12_1_port);
   bht_reg_14_1_inst : DLH_X1 port map( G => N3028, D => N3735, Q => 
                           bht_14_1_port);
   bht_reg_16_1_inst : DLH_X1 port map( G => N2920, D => N3735, Q => 
                           bht_16_1_port);
   bht_reg_18_1_inst : DLH_X1 port map( G => N2812, D => N3735, Q => 
                           bht_18_1_port);
   bht_reg_20_1_inst : DLH_X1 port map( G => N2704, D => N3735, Q => 
                           bht_20_1_port);
   bht_reg_22_1_inst : DLH_X1 port map( G => N2596, D => N3735, Q => 
                           bht_22_1_port);
   bht_reg_24_1_inst : DLH_X1 port map( G => N2488, D => N3735, Q => 
                           bht_24_1_port);
   bht_reg_26_1_inst : DLH_X1 port map( G => N2380, D => N3735, Q => 
                           bht_26_1_port);
   bht_reg_28_1_inst : DLH_X1 port map( G => N2272, D => N3735, Q => 
                           bht_28_1_port);
   bht_reg_30_1_inst : DLH_X1 port map( G => N2164, D => N3735, Q => 
                           bht_30_1_port);
   bht_reg_31_1_inst : DLH_X1 port map( G => N2110, D => N3735, Q => 
                           bht_31_1_port);
   bht_reg_29_1_inst : DLH_X1 port map( G => N2218, D => N3735, Q => 
                           bht_29_1_port);
   bht_reg_27_1_inst : DLH_X1 port map( G => N2326, D => N3735, Q => 
                           bht_27_1_port);
   bht_reg_25_1_inst : DLH_X1 port map( G => N2434, D => N3735, Q => 
                           bht_25_1_port);
   bht_reg_23_1_inst : DLH_X1 port map( G => N2542, D => N3735, Q => 
                           bht_23_1_port);
   bht_reg_21_1_inst : DLH_X1 port map( G => N2650, D => N3735, Q => 
                           bht_21_1_port);
   bht_reg_19_1_inst : DLH_X1 port map( G => N2758, D => N3735, Q => 
                           bht_19_1_port);
   bht_reg_17_1_inst : DLH_X1 port map( G => N2866, D => N3735, Q => 
                           bht_17_1_port);
   bht_reg_15_1_inst : DLH_X1 port map( G => N2974, D => N3735, Q => 
                           bht_15_1_port);
   bht_reg_13_1_inst : DLH_X1 port map( G => N3082, D => N3735, Q => 
                           bht_13_1_port);
   bht_reg_11_1_inst : DLH_X1 port map( G => N3190, D => N3735, Q => 
                           bht_11_1_port);
   bht_reg_9_1_inst : DLH_X1 port map( G => N3298, D => N3735, Q => 
                           bht_9_1_port);
   bht_reg_7_1_inst : DLH_X1 port map( G => N3406, D => N3735, Q => 
                           bht_7_1_port);
   bht_reg_5_1_inst : DLH_X1 port map( G => N3514, D => N3735, Q => 
                           bht_5_1_port);
   bht_reg_3_1_inst : DLH_X1 port map( G => N3622, D => N3735, Q => 
                           bht_3_1_port);
   bht_reg_1_1_inst : DLH_X1 port map( G => N3730, D => N3735, Q => 
                           bht_1_1_port);
   entry_r_reg_1_inst : DLH_X1 port map( G => N188, D => N126, Q => 
                           entry_r_1_port);
   entry_r_delay_reg_1_inst : DFFR_X1 port map( D => entry_r_1_port, CK => clk,
                           RN => rst, Q => n3, QN => net108065);
   entry_r_reg_25_inst : DLH_X1 port map( G => N188, D => N150, Q => 
                           entry_r_25_port);
   entry_r_delay_reg_25_inst : DFFR_X1 port map( D => entry_r_25_port, CK => 
                           clk, RN => rst, Q => net108064, QN => n9);
   bht_reg_0_25_inst : DLH_X1 port map( G => N3784, D => N3783, Q => 
                           bht_0_25_port);
   bht_reg_2_25_inst : DLH_X1 port map( G => N3676, D => N3783, Q => 
                           bht_2_25_port);
   bht_reg_4_25_inst : DLH_X1 port map( G => N3568, D => N3783, Q => 
                           bht_4_25_port);
   bht_reg_6_25_inst : DLH_X1 port map( G => N3460, D => N3783, Q => 
                           bht_6_25_port);
   bht_reg_8_25_inst : DLH_X1 port map( G => N3352, D => N3783, Q => 
                           bht_8_25_port);
   bht_reg_10_25_inst : DLH_X1 port map( G => N3244, D => N3783, Q => 
                           bht_10_25_port);
   bht_reg_12_25_inst : DLH_X1 port map( G => N3136, D => N3783, Q => 
                           bht_12_25_port);
   bht_reg_14_25_inst : DLH_X1 port map( G => N3028, D => N3783, Q => 
                           bht_14_25_port);
   bht_reg_16_25_inst : DLH_X1 port map( G => N2920, D => N3783, Q => 
                           bht_16_25_port);
   bht_reg_18_25_inst : DLH_X1 port map( G => N2812, D => N3783, Q => 
                           bht_18_25_port);
   bht_reg_20_25_inst : DLH_X1 port map( G => N2704, D => N3783, Q => 
                           bht_20_25_port);
   bht_reg_22_25_inst : DLH_X1 port map( G => N2596, D => N3783, Q => 
                           bht_22_25_port);
   bht_reg_24_25_inst : DLH_X1 port map( G => N2488, D => N3783, Q => 
                           bht_24_25_port);
   bht_reg_26_25_inst : DLH_X1 port map( G => N2380, D => N3783, Q => 
                           bht_26_25_port);
   bht_reg_28_25_inst : DLH_X1 port map( G => N2272, D => N3783, Q => 
                           bht_28_25_port);
   bht_reg_30_25_inst : DLH_X1 port map( G => N2164, D => N3783, Q => 
                           bht_30_25_port);
   bht_reg_29_25_inst : DLH_X1 port map( G => N2218, D => N3783, Q => 
                           bht_29_25_port);
   bht_reg_27_25_inst : DLH_X1 port map( G => N2326, D => N3783, Q => 
                           bht_27_25_port);
   bht_reg_25_25_inst : DLH_X1 port map( G => N2434, D => N3783, Q => 
                           bht_25_25_port);
   bht_reg_23_25_inst : DLH_X1 port map( G => N2542, D => N3783, Q => 
                           bht_23_25_port);
   bht_reg_21_25_inst : DLH_X1 port map( G => N2650, D => N3783, Q => 
                           bht_21_25_port);
   bht_reg_19_25_inst : DLH_X1 port map( G => N2758, D => N3783, Q => 
                           bht_19_25_port);
   bht_reg_17_25_inst : DLH_X1 port map( G => N2866, D => N3783, Q => 
                           bht_17_25_port);
   bht_reg_15_25_inst : DLH_X1 port map( G => N2974, D => N3783, Q => 
                           bht_15_25_port);
   bht_reg_13_25_inst : DLH_X1 port map( G => N3082, D => N3783, Q => 
                           bht_13_25_port);
   bht_reg_11_25_inst : DLH_X1 port map( G => N3190, D => N3783, Q => 
                           bht_11_25_port);
   bht_reg_9_25_inst : DLH_X1 port map( G => N3298, D => N3783, Q => 
                           bht_9_25_port);
   bht_reg_7_25_inst : DLH_X1 port map( G => N3406, D => N3783, Q => 
                           bht_7_25_port);
   bht_reg_5_25_inst : DLH_X1 port map( G => N3514, D => N3783, Q => 
                           bht_5_25_port);
   bht_reg_3_25_inst : DLH_X1 port map( G => N3622, D => N3783, Q => 
                           bht_3_25_port);
   bht_reg_1_25_inst : DLH_X1 port map( G => N3730, D => N3783, Q => 
                           bht_1_25_port);
   U3 : AND2_X2 port map( A1 => n761, A2 => n758, ZN => n121);
   U4 : AND2_X2 port map( A1 => n770, A2 => n762, ZN => n135_port);
   U5 : AND2_X2 port map( A1 => n776, A2 => n759, ZN => n143_port);
   U6 : AND2_X2 port map( A1 => n783, A2 => n763, ZN => n161);
   U7 : OAI21_X2 port map( B1 => n72, B2 => n75, A => rst, ZN => N2110);
   U8 : OAI21_X2 port map( B1 => n69, B2 => n73, A => rst, ZN => N3136);
   U9 : OAI21_X2 port map( B1 => n71, B2 => n74, A => rst, ZN => N2596);
   U10 : OAI21_X2 port map( B1 => n45, B2 => n46, A => rst, ZN => N3784);
   U11 : AND2_X2 port map( A1 => n762, A2 => n758, ZN => n123);
   U12 : AND2_X2 port map( A1 => n770, A2 => n761, ZN => n133_port);
   U13 : AND2_X2 port map( A1 => n783, A2 => n759, ZN => n155);
   U14 : AND2_X2 port map( A1 => n776, A2 => n763, ZN => n149_port);
   U15 : OAI21_X2 port map( B1 => n68, B2 => n75, A => rst, ZN => N2326);
   U16 : OAI21_X2 port map( B1 => n66, B2 => n74, A => rst, ZN => N2866);
   U17 : OAI21_X2 port map( B1 => n70, B2 => n73, A => rst, ZN => N3082);
   U18 : OAI21_X2 port map( B1 => n45, B2 => n67, A => rst, ZN => N3676);
   U19 : AND2_X2 port map( A1 => n758, A2 => n759, ZN => n119);
   U20 : AND2_X2 port map( A1 => n770, A2 => n763, ZN => n137_port);
   U21 : AND2_X2 port map( A1 => n783, A2 => n761, ZN => n157);
   U22 : AND2_X2 port map( A1 => n776, A2 => n762, ZN => n147_port);
   U23 : OAI21_X2 port map( B1 => n66, B2 => n75, A => rst, ZN => N2434);
   U24 : OAI21_X2 port map( B1 => n67, B2 => n73, A => rst, ZN => N3244);
   U25 : OAI21_X2 port map( B1 => n46, B2 => n74, A => rst, ZN => N2920);
   U26 : OAI21_X2 port map( B1 => n45, B2 => n69, A => rst, ZN => N3568);
   U27 : AND2_X2 port map( A1 => n763, A2 => n758, ZN => n125_port);
   U28 : AND2_X2 port map( A1 => n770, A2 => n759, ZN => n131_port);
   U29 : AND2_X2 port map( A1 => n783, A2 => n762, ZN => n159);
   U30 : AND2_X2 port map( A1 => n776, A2 => n761, ZN => n145_port);
   U31 : OAI21_X2 port map( B1 => n70, B2 => n75, A => rst, ZN => N2218);
   U32 : OAI21_X2 port map( B1 => n68, B2 => n74, A => rst, ZN => N2758);
   U33 : OAI21_X2 port map( B1 => n66, B2 => n73, A => rst, ZN => N3298);
   U34 : OAI21_X2 port map( B1 => n45, B2 => n71, A => rst, ZN => N3460);
   U35 : AND2_X2 port map( A1 => n761, A2 => n760, ZN => n120);
   U36 : AND2_X2 port map( A1 => n771, A2 => n762, ZN => n134_port);
   U37 : AND2_X2 port map( A1 => n777, A2 => n759, ZN => n142_port);
   U38 : AND2_X2 port map( A1 => n784, A2 => n763, ZN => n160);
   U39 : OAI21_X2 port map( B1 => n46, B2 => n73, A => rst, ZN => N3352);
   U40 : OAI21_X2 port map( B1 => n69, B2 => n74, A => rst, ZN => N2704);
   U41 : OAI21_X2 port map( B1 => n67, B2 => n75, A => rst, ZN => N2380);
   U42 : OAI21_X2 port map( B1 => n45, B2 => n72, A => rst, ZN => N3406);
   U43 : AND2_X2 port map( A1 => n762, A2 => n760, ZN => n122);
   U44 : AND2_X2 port map( A1 => n771, A2 => n761, ZN => n132_port);
   U45 : AND2_X2 port map( A1 => n784, A2 => n759, ZN => n154);
   U46 : AND2_X2 port map( A1 => n777, A2 => n763, ZN => n148_port);
   U47 : OAI21_X2 port map( B1 => n71, B2 => n73, A => rst, ZN => N3028);
   U48 : OAI21_X2 port map( B1 => n72, B2 => n74, A => rst, ZN => N2542);
   U49 : OAI21_X2 port map( B1 => n46, B2 => n75, A => rst, ZN => N2488);
   U50 : OAI21_X2 port map( B1 => n45, B2 => n70, A => rst, ZN => N3514);
   U51 : OAI22_X4 port map( A1 => n49, A2 => n43, B1 => n47, B2 => n50, ZN => 
                           N3733);
   U52 : AND2_X2 port map( A1 => n760, A2 => n759, ZN => n118);
   U53 : AND2_X2 port map( A1 => n771, A2 => n763, ZN => n136_port);
   U54 : AND2_X2 port map( A1 => n784, A2 => n761, ZN => n156);
   U55 : AND2_X2 port map( A1 => n777, A2 => n762, ZN => n146_port);
   U56 : OAI21_X2 port map( B1 => n67, B2 => n74, A => rst, ZN => N2812);
   U57 : OAI21_X2 port map( B1 => n69, B2 => n75, A => rst, ZN => N2272);
   U58 : OAI21_X2 port map( B1 => n72, B2 => n73, A => rst, ZN => N2974);
   U59 : OAI21_X2 port map( B1 => n45, B2 => n68, A => rst, ZN => N3622);
   U60 : INV_X2 port map( A => rst, ZN => n44);
   U61 : OAI22_X4 port map( A1 => n207, A2 => n43, B1 => n47, B2 => n48, ZN => 
                           N3735);
   U62 : AND2_X2 port map( A1 => n763, A2 => n760, ZN => n124);
   U63 : AND2_X2 port map( A1 => n771, A2 => n759, ZN => n130_port);
   U64 : AND2_X2 port map( A1 => n784, A2 => n762, ZN => n158);
   U65 : AND2_X2 port map( A1 => n777, A2 => n761, ZN => n144_port);
   U66 : OAI21_X2 port map( B1 => n71, B2 => n75, A => rst, ZN => N2164);
   U67 : OAI21_X2 port map( B1 => n70, B2 => n74, A => rst, ZN => N2650);
   U68 : OAI21_X2 port map( B1 => n68, B2 => n73, A => rst, ZN => N3190);
   U69 : OAI21_X2 port map( B1 => n45, B2 => n66, A => rst, ZN => N3730);
   U70 : NAND4_X2 port map( A1 => n163, A2 => n164, A3 => n165, A4 => n166, ZN 
                           => n42);
   U71 : NOR2_X2 port map( A1 => n9, A2 => n44, ZN => N3783);
   U72 : NOR2_X2 port map( A1 => n33, A2 => n44, ZN => N3785);
   U73 : NOR2_X2 port map( A1 => n32, A2 => n44, ZN => N3781);
   U74 : NOR2_X2 port map( A1 => n31, A2 => n44, ZN => N3779);
   U75 : NOR2_X2 port map( A1 => n30, A2 => n44, ZN => N3777);
   U76 : NOR2_X2 port map( A1 => n29, A2 => n44, ZN => N3775);
   U77 : NOR2_X2 port map( A1 => n28, A2 => n44, ZN => N3773);
   U78 : NOR2_X2 port map( A1 => n27, A2 => n44, ZN => N3771);
   U79 : NOR2_X2 port map( A1 => n26, A2 => n44, ZN => N3769);
   U80 : NOR2_X2 port map( A1 => n25, A2 => n44, ZN => N3767);
   U81 : NOR2_X2 port map( A1 => n24, A2 => n44, ZN => N3765);
   U82 : NOR2_X2 port map( A1 => n23, A2 => n44, ZN => N3763);
   U83 : NOR2_X2 port map( A1 => n22, A2 => n44, ZN => N3761);
   U84 : NOR2_X2 port map( A1 => n21, A2 => n44, ZN => N3759);
   U85 : NOR2_X2 port map( A1 => n20, A2 => n44, ZN => N3757);
   U86 : NOR2_X2 port map( A1 => n19, A2 => n44, ZN => N3755);
   U87 : NOR2_X2 port map( A1 => n18, A2 => n44, ZN => N3753);
   U88 : NOR2_X2 port map( A1 => n17, A2 => n44, ZN => N3751);
   U89 : NOR2_X2 port map( A1 => n16, A2 => n44, ZN => N3749);
   U90 : NOR2_X2 port map( A1 => n15, A2 => n44, ZN => N3747);
   U91 : NOR2_X2 port map( A1 => n14, A2 => n44, ZN => N3745);
   U92 : NOR2_X2 port map( A1 => n13, A2 => n44, ZN => N3743);
   U93 : NOR2_X2 port map( A1 => n12, A2 => n44, ZN => N3741);
   U94 : NOR2_X2 port map( A1 => n11, A2 => n44, ZN => N3739);
   U95 : NOR2_X2 port map( A1 => n10, A2 => n44, ZN => N3737);
   U96 : NOR2_X4 port map( A1 => n43, A2 => n6, ZN => sig_bpw);
   U97 : OAI21_X1 port map( B1 => n36, B2 => n37, A => n38, ZN => sig_brt_tmp);
   U98 : NAND4_X1 port map( A1 => rst, A2 => opcd(2), A3 => n39, A4 => n40, ZN 
                           => n38);
   U99 : NOR4_X1 port map( A1 => sig_bal, A2 => opcd(5), A3 => opcd(4), A4 => 
                           opcd(3), ZN => n40);
   U100 : NOR2_X1 port map( A1 => opcd(1), A2 => n41, ZN => n39);
   U101 : XOR2_X1 port map( A => n42, B => opcd(0), Z => n41);
   U102 : INV_X1 port map( A => N126, ZN => n36);
   U103 : NAND2_X1 port map( A1 => rst, A2 => n3, ZN => n48);
   U104 : NAND2_X1 port map( A1 => sig_brt_delay, A2 => rst, ZN => n50);
   U105 : NAND2_X1 port map( A1 => rst, A2 => n47, ZN => n43);
   U106 : NAND4_X1 port map( A1 => opcd_delay_2_port, A2 => n214, A3 => n51, A4
                           => n52, ZN => n47);
   U107 : NOR3_X1 port map( A1 => opcd_delay_3_port, A2 => opcd_delay_5_port, 
                           A3 => opcd_delay_4_port, ZN => n52);
   U108 : XOR2_X1 port map( A => n53, B => n54, Z => n51);
   U109 : NOR2_X1 port map( A1 => n55, A2 => n56, ZN => n54);
   U110 : NAND4_X1 port map( A1 => n57, A2 => n58, A3 => n59, A4 => n60, ZN => 
                           n56);
   U111 : NOR4_X1 port map( A1 => ld_a(23), A2 => ld_a(22), A3 => ld_a(21), A4 
                           => ld_a(20), ZN => n60);
   U112 : NOR4_X1 port map( A1 => ld_a(1), A2 => ld_a(19), A3 => ld_a(18), A4 
                           => ld_a(17), ZN => n59);
   U113 : NOR4_X1 port map( A1 => ld_a(16), A2 => ld_a(15), A3 => ld_a(14), A4 
                           => ld_a(13), ZN => n58);
   U114 : NOR4_X1 port map( A1 => ld_a(12), A2 => ld_a(11), A3 => ld_a(10), A4 
                           => ld_a(0), ZN => n57);
   U115 : NAND4_X1 port map( A1 => n61, A2 => n62, A3 => n63, A4 => n64, ZN => 
                           n55);
   U116 : NOR4_X1 port map( A1 => ld_a(9), A2 => ld_a(8), A3 => ld_a(7), A4 => 
                           ld_a(6), ZN => n64);
   U117 : NOR4_X1 port map( A1 => ld_a(5), A2 => ld_a(4), A3 => ld_a(3), A4 => 
                           ld_a(31), ZN => n63);
   U118 : NOR4_X1 port map( A1 => ld_a(30), A2 => ld_a(2), A3 => ld_a(29), A4 
                           => ld_a(28), ZN => n62);
   U119 : NOR4_X1 port map( A1 => ld_a(27), A2 => ld_a(26), A3 => ld_a(25), A4 
                           => ld_a(24), ZN => n61);
   U120 : XNOR2_X1 port map( A => n219, B => n7, ZN => n53);
   U121 : AOI22_X1 port map( A1 => n65, A2 => n7, B1 => n207, B2 => n3, ZN => 
                           n49);
   U122 : OR2_X1 port map( A1 => n3, A2 => n207, ZN => n65);
   U123 : NAND3_X1 port map( A1 => n187, A2 => sig_bal_delay, A3 => n35, ZN => 
                           n45);
   U124 : NAND3_X1 port map( A1 => sig_bal_delay, A2 => n8, A3 => n35, ZN => 
                           n73);
   U125 : NAND3_X1 port map( A1 => sig_bal_delay, A2 => n4, A3 => n187, ZN => 
                           n74);
   U126 : NAND3_X1 port map( A1 => n202, A2 => n200, A3 => n34, ZN => n46);
   U127 : NAND3_X1 port map( A1 => n202, A2 => n2, A3 => n34, ZN => n66);
   U128 : NAND3_X1 port map( A1 => n200, A2 => n5, A3 => n34, ZN => n67);
   U129 : NAND3_X1 port map( A1 => n2, A2 => n5, A3 => n34, ZN => n68);
   U130 : NAND3_X1 port map( A1 => n200, A2 => n1, A3 => n202, ZN => n69);
   U131 : NAND3_X1 port map( A1 => n2, A2 => n1, A3 => n202, ZN => n70);
   U132 : NAND3_X1 port map( A1 => n5, A2 => n1, A3 => n200, ZN => n71);
   U133 : NAND3_X1 port map( A1 => n8, A2 => n4, A3 => sig_bal_delay, ZN => n75
                           );
   U134 : NAND3_X1 port map( A1 => n5, A2 => n1, A3 => n2, ZN => n72);
   U135 : INV_X1 port map( A => n37, ZN => N188);
   U136 : NAND2_X1 port map( A1 => rst, A2 => sig_bal, ZN => n37);
   U137 : MUX2_X1 port map( A => n76, B => addr(31), S => n42, Z => N151);
   U138 : MUX2_X1 port map( A => n77, B => addr(30), S => n42, Z => N150);
   U139 : MUX2_X1 port map( A => n78, B => addr(29), S => n42, Z => N149);
   U140 : INV_X1 port map( A => n79, ZN => n78);
   U141 : MUX2_X1 port map( A => n80, B => addr(28), S => n42, Z => N148);
   U142 : INV_X1 port map( A => n81, ZN => n80);
   U143 : MUX2_X1 port map( A => n82, B => addr(27), S => n42, Z => N147);
   U144 : MUX2_X1 port map( A => n83, B => addr(26), S => n42, Z => N146);
   U145 : MUX2_X1 port map( A => n84, B => addr(25), S => n42, Z => N145);
   U146 : MUX2_X1 port map( A => n85, B => addr(24), S => n42, Z => N144);
   U147 : MUX2_X1 port map( A => n86, B => addr(23), S => n42, Z => N143);
   U148 : MUX2_X1 port map( A => n87, B => addr(22), S => n42, Z => N142);
   U149 : MUX2_X1 port map( A => n88, B => addr(21), S => n42, Z => N141);
   U150 : MUX2_X1 port map( A => n89, B => addr(20), S => n42, Z => N140);
   U151 : MUX2_X1 port map( A => n90, B => addr(19), S => n42, Z => N139);
   U152 : INV_X1 port map( A => n91, ZN => n90);
   U153 : MUX2_X1 port map( A => n92, B => addr(18), S => n42, Z => N138);
   U154 : INV_X1 port map( A => n93, ZN => n92);
   U155 : MUX2_X1 port map( A => n94, B => addr(17), S => n42, Z => N137);
   U156 : INV_X1 port map( A => n95, ZN => n94);
   U157 : MUX2_X1 port map( A => n96, B => addr(16), S => n42, Z => N136);
   U158 : MUX2_X1 port map( A => n97, B => addr(15), S => n42, Z => N135);
   U159 : MUX2_X1 port map( A => n98, B => addr(14), S => n42, Z => N134);
   U160 : MUX2_X1 port map( A => n99, B => addr(13), S => n42, Z => N133);
   U161 : INV_X1 port map( A => n100, ZN => n99);
   U162 : MUX2_X1 port map( A => n101, B => addr(12), S => n42, Z => N132);
   U163 : INV_X1 port map( A => n102, ZN => n101);
   U164 : MUX2_X1 port map( A => n103, B => addr(11), S => n42, Z => N131);
   U165 : MUX2_X1 port map( A => n104, B => addr(10), S => n42, Z => N130);
   U166 : MUX2_X1 port map( A => n105, B => addr(9), S => n42, Z => N129);
   U167 : INV_X1 port map( A => n106, ZN => n105);
   U168 : MUX2_X1 port map( A => n107, B => addr(8), S => n42, Z => N128);
   U169 : MUX2_X1 port map( A => n108, B => addr(7), S => n42, Z => N127);
   U170 : NOR2_X1 port map( A1 => n109, A2 => n42, ZN => N126);
   U171 : NOR4_X1 port map( A1 => n110, A2 => n111, A3 => n112, A4 => n113, ZN 
                           => n109);
   U172 : NAND4_X1 port map( A1 => n114, A2 => n115, A3 => n116, A4 => n117, ZN
                           => n113);
   U173 : AOI22_X1 port map( A1 => bht_14_1_port, A2 => n118, B1 => 
                           bht_15_1_port, B2 => n119, ZN => n117);
   U174 : AOI22_X1 port map( A1 => bht_12_1_port, A2 => n120, B1 => 
                           bht_13_1_port, B2 => n121, ZN => n116);
   U175 : AOI22_X1 port map( A1 => bht_10_1_port, A2 => n122, B1 => 
                           bht_11_1_port, B2 => n123, ZN => n115);
   U176 : AOI22_X1 port map( A1 => bht_8_1_port, A2 => n124, B1 => bht_9_1_port
                           , B2 => n125_port, ZN => n114);
   U177 : NAND4_X1 port map( A1 => n126_port, A2 => n127_port, A3 => n128_port,
                           A4 => n129_port, ZN => n112);
   U178 : AOI22_X1 port map( A1 => bht_6_1_port, A2 => n130_port, B1 => 
                           bht_7_1_port, B2 => n131_port, ZN => n129_port);
   U179 : AOI22_X1 port map( A1 => bht_4_1_port, A2 => n132_port, B1 => 
                           bht_5_1_port, B2 => n133_port, ZN => n128_port);
   U180 : AOI22_X1 port map( A1 => bht_2_1_port, A2 => n134_port, B1 => 
                           bht_3_1_port, B2 => n135_port, ZN => n127_port);
   U181 : AOI22_X1 port map( A1 => bht_0_1_port, A2 => n136_port, B1 => 
                           bht_1_1_port, B2 => n137_port, ZN => n126_port);
   U182 : NAND4_X1 port map( A1 => n138_port, A2 => n139_port, A3 => n140_port,
                           A4 => n141_port, ZN => n111);
   U183 : AOI22_X1 port map( A1 => bht_30_1_port, A2 => n142_port, B1 => 
                           bht_31_1_port, B2 => n143_port, ZN => n141_port);
   U184 : AOI22_X1 port map( A1 => bht_28_1_port, A2 => n144_port, B1 => 
                           bht_29_1_port, B2 => n145_port, ZN => n140_port);
   U185 : AOI22_X1 port map( A1 => bht_26_1_port, A2 => n146_port, B1 => 
                           bht_27_1_port, B2 => n147_port, ZN => n139_port);
   U186 : AOI22_X1 port map( A1 => bht_24_1_port, A2 => n148_port, B1 => 
                           bht_25_1_port, B2 => n149_port, ZN => n138_port);
   U187 : NAND4_X1 port map( A1 => n150_port, A2 => n151_port, A3 => n152, A4 
                           => n153, ZN => n110);
   U188 : AOI22_X1 port map( A1 => bht_22_1_port, A2 => n154, B1 => 
                           bht_23_1_port, B2 => n155, ZN => n153);
   U189 : AOI22_X1 port map( A1 => bht_20_1_port, A2 => n156, B1 => 
                           bht_21_1_port, B2 => n157, ZN => n152);
   U190 : AOI22_X1 port map( A1 => bht_18_1_port, A2 => n158, B1 => 
                           bht_19_1_port, B2 => n159, ZN => n151_port);
   U191 : AOI22_X1 port map( A1 => bht_16_1_port, A2 => n160, B1 => 
                           bht_17_1_port, B2 => n161, ZN => n150_port);
   U192 : NOR2_X1 port map( A1 => n162, A2 => n42, ZN => N125);
   U193 : NOR4_X1 port map( A1 => n167, A2 => n168, A3 => n169, A4 => n170, ZN 
                           => n166);
   U194 : OAI222_X1 port map( A1 => n171, A2 => n87, B1 => n172, B2 => n88, C1 
                           => n173, C2 => n86, ZN => n170);
   U195 : OAI222_X1 port map( A1 => n174, A2 => n82, B1 => n175, B2 => n83, C1 
                           => n176, C2 => n89, ZN => n169);
   U196 : OAI222_X1 port map( A1 => n177, A2 => n85, B1 => n178, B2 => n76, C1 
                           => n179, C2 => n84, ZN => n168);
   U197 : INV_X1 port map( A => n180, ZN => n167);
   U198 : AOI222_X1 port map( A1 => n181, A2 => n79, B1 => n182, B2 => n81, C1 
                           => n183, C2 => n184, ZN => n180);
   U199 : AOI211_X1 port map( C1 => n106, C2 => n185, A => n186, B => n188_port
                           , ZN => n165);
   U200 : OAI22_X1 port map( A1 => n189, A2 => n97, B1 => n190, B2 => n98, ZN 
                           => n188_port);
   U201 : INV_X1 port map( A => n191, ZN => n97);
   U202 : INV_X1 port map( A => n192, ZN => n189);
   U203 : OAI221_X1 port map( B1 => n193, B2 => n104, C1 => n194, C2 => n103, A
                           => n195, ZN => n186);
   U204 : MUX2_X1 port map( A => n196, B => n197, S => sig_bal, Z => n195);
   U205 : NOR4_X1 port map( A1 => n198, A2 => n199, A3 => n201, A4 => n203, ZN 
                           => n197);
   U206 : OAI211_X1 port map( C1 => n204, C2 => n205, A => n206, B => n208, ZN 
                           => n203);
   U207 : XNOR2_X1 port map( A => addr(8), B => n107, ZN => n208);
   U208 : OR4_X1 port map( A1 => n209, A2 => n210, A3 => n211, A4 => n212, ZN 
                           => n107);
   U209 : NAND4_X1 port map( A1 => n213, A2 => n215, A3 => n216, A4 => n217, ZN
                           => n212);
   U210 : AOI22_X1 port map( A1 => bht_6_3_port, A2 => n130_port, B1 => 
                           bht_7_3_port, B2 => n131_port, ZN => n217);
   U211 : AOI22_X1 port map( A1 => bht_4_3_port, A2 => n132_port, B1 => 
                           bht_5_3_port, B2 => n133_port, ZN => n216);
   U212 : AOI22_X1 port map( A1 => bht_2_3_port, A2 => n134_port, B1 => 
                           bht_3_3_port, B2 => n135_port, ZN => n215);
   U213 : AOI22_X1 port map( A1 => bht_0_3_port, A2 => n136_port, B1 => 
                           bht_1_3_port, B2 => n137_port, ZN => n213);
   U214 : NAND4_X1 port map( A1 => n218, A2 => n220, A3 => n221, A4 => n222, ZN
                           => n211);
   U215 : AOI22_X1 port map( A1 => bht_14_3_port, A2 => n118, B1 => 
                           bht_15_3_port, B2 => n119, ZN => n222);
   U216 : AOI22_X1 port map( A1 => bht_12_3_port, A2 => n120, B1 => 
                           bht_13_3_port, B2 => n121, ZN => n221);
   U217 : AOI22_X1 port map( A1 => bht_10_3_port, A2 => n122, B1 => 
                           bht_11_3_port, B2 => n123, ZN => n220);
   U218 : AOI22_X1 port map( A1 => bht_8_3_port, A2 => n124, B1 => bht_9_3_port
                           , B2 => n125_port, ZN => n218);
   U219 : NAND4_X1 port map( A1 => n223, A2 => n224, A3 => n225, A4 => n226, ZN
                           => n210);
   U220 : AOI22_X1 port map( A1 => bht_22_3_port, A2 => n154, B1 => 
                           bht_23_3_port, B2 => n155, ZN => n226);
   U221 : AOI22_X1 port map( A1 => bht_20_3_port, A2 => n156, B1 => 
                           bht_21_3_port, B2 => n157, ZN => n225);
   U222 : AOI22_X1 port map( A1 => bht_18_3_port, A2 => n158, B1 => 
                           bht_19_3_port, B2 => n159, ZN => n224);
   U223 : AOI22_X1 port map( A1 => bht_16_3_port, A2 => n160, B1 => 
                           bht_17_3_port, B2 => n161, ZN => n223);
   U224 : NAND4_X1 port map( A1 => n227, A2 => n228, A3 => n229, A4 => n230, ZN
                           => n209);
   U225 : AOI22_X1 port map( A1 => bht_30_3_port, A2 => n142_port, B1 => 
                           bht_31_3_port, B2 => n143_port, ZN => n230);
   U226 : AOI22_X1 port map( A1 => bht_28_3_port, A2 => n144_port, B1 => 
                           bht_29_3_port, B2 => n145_port, ZN => n229);
   U227 : AOI22_X1 port map( A1 => bht_26_3_port, A2 => n146_port, B1 => 
                           bht_27_3_port, B2 => n147_port, ZN => n228);
   U228 : AOI22_X1 port map( A1 => bht_24_3_port, A2 => n148_port, B1 => 
                           bht_25_3_port, B2 => n149_port, ZN => n227);
   U229 : XNOR2_X1 port map( A => addr(7), B => n108, ZN => n206);
   U230 : OR4_X1 port map( A1 => n231, A2 => n232, A3 => n233, A4 => n234, ZN 
                           => n108);
   U231 : NAND4_X1 port map( A1 => n235, A2 => n236, A3 => n237, A4 => n238, ZN
                           => n234);
   U232 : AOI22_X1 port map( A1 => bht_6_2_port, A2 => n130_port, B1 => 
                           bht_7_2_port, B2 => n131_port, ZN => n238);
   U233 : AOI22_X1 port map( A1 => bht_4_2_port, A2 => n132_port, B1 => 
                           bht_5_2_port, B2 => n133_port, ZN => n237);
   U234 : AOI22_X1 port map( A1 => bht_2_2_port, A2 => n134_port, B1 => 
                           bht_3_2_port, B2 => n135_port, ZN => n236);
   U235 : AOI22_X1 port map( A1 => bht_0_2_port, A2 => n136_port, B1 => 
                           bht_1_2_port, B2 => n137_port, ZN => n235);
   U236 : NAND4_X1 port map( A1 => n239, A2 => n240, A3 => n241, A4 => n242, ZN
                           => n233);
   U237 : AOI22_X1 port map( A1 => bht_14_2_port, A2 => n118, B1 => 
                           bht_15_2_port, B2 => n119, ZN => n242);
   U238 : AOI22_X1 port map( A1 => bht_12_2_port, A2 => n120, B1 => 
                           bht_13_2_port, B2 => n121, ZN => n241);
   U239 : AOI22_X1 port map( A1 => bht_10_2_port, A2 => n122, B1 => 
                           bht_11_2_port, B2 => n123, ZN => n240);
   U240 : AOI22_X1 port map( A1 => bht_8_2_port, A2 => n124, B1 => bht_9_2_port
                           , B2 => n125_port, ZN => n239);
   U241 : NAND4_X1 port map( A1 => n243, A2 => n244, A3 => n245, A4 => n246, ZN
                           => n232);
   U242 : AOI22_X1 port map( A1 => bht_22_2_port, A2 => n154, B1 => 
                           bht_23_2_port, B2 => n155, ZN => n246);
   U243 : AOI22_X1 port map( A1 => bht_20_2_port, A2 => n156, B1 => 
                           bht_21_2_port, B2 => n157, ZN => n245);
   U244 : AOI22_X1 port map( A1 => bht_18_2_port, A2 => n158, B1 => 
                           bht_19_2_port, B2 => n159, ZN => n244);
   U245 : AOI22_X1 port map( A1 => bht_16_2_port, A2 => n160, B1 => 
                           bht_17_2_port, B2 => n161, ZN => n243);
   U246 : NAND4_X1 port map( A1 => n247, A2 => n248, A3 => n249, A4 => n250, ZN
                           => n231);
   U247 : AOI22_X1 port map( A1 => bht_30_2_port, A2 => n142_port, B1 => 
                           bht_31_2_port, B2 => n143_port, ZN => n250);
   U248 : AOI22_X1 port map( A1 => bht_28_2_port, A2 => n144_port, B1 => 
                           bht_29_2_port, B2 => n145_port, ZN => n249);
   U249 : AOI22_X1 port map( A1 => bht_26_2_port, A2 => n146_port, B1 => 
                           bht_27_2_port, B2 => n147_port, ZN => n248);
   U250 : AOI22_X1 port map( A1 => bht_24_2_port, A2 => n148_port, B1 => 
                           bht_25_2_port, B2 => n149_port, ZN => n247);
   U251 : OAI222_X1 port map( A1 => n106, A2 => n185, B1 => n191, B2 => n192, 
                           C1 => n251, C2 => n252, ZN => n201);
   U252 : NOR4_X1 port map( A1 => n253, A2 => n254, A3 => n255, A4 => n256, ZN 
                           => n191);
   U253 : NAND4_X1 port map( A1 => n257, A2 => n258, A3 => n259, A4 => n260, ZN
                           => n256);
   U254 : AOI22_X1 port map( A1 => bht_6_10_port, A2 => n130_port, B1 => 
                           bht_7_10_port, B2 => n131_port, ZN => n260);
   U255 : AOI22_X1 port map( A1 => bht_4_10_port, A2 => n132_port, B1 => 
                           bht_5_10_port, B2 => n133_port, ZN => n259);
   U256 : AOI22_X1 port map( A1 => bht_2_10_port, A2 => n134_port, B1 => 
                           bht_3_10_port, B2 => n135_port, ZN => n258);
   U257 : AOI22_X1 port map( A1 => bht_0_10_port, A2 => n136_port, B1 => 
                           bht_1_10_port, B2 => n137_port, ZN => n257);
   U258 : NAND4_X1 port map( A1 => n261, A2 => n262, A3 => n263, A4 => n264, ZN
                           => n255);
   U259 : AOI22_X1 port map( A1 => bht_14_10_port, A2 => n118, B1 => 
                           bht_15_10_port, B2 => n119, ZN => n264);
   U260 : AOI22_X1 port map( A1 => bht_12_10_port, A2 => n120, B1 => 
                           bht_13_10_port, B2 => n121, ZN => n263);
   U261 : AOI22_X1 port map( A1 => bht_10_10_port, A2 => n122, B1 => 
                           bht_11_10_port, B2 => n123, ZN => n262);
   U262 : AOI22_X1 port map( A1 => bht_8_10_port, A2 => n124, B1 => 
                           bht_9_10_port, B2 => n125_port, ZN => n261);
   U263 : NAND4_X1 port map( A1 => n265, A2 => n266, A3 => n267, A4 => n268, ZN
                           => n254);
   U264 : AOI22_X1 port map( A1 => bht_22_10_port, A2 => n154, B1 => 
                           bht_23_10_port, B2 => n155, ZN => n268);
   U265 : AOI22_X1 port map( A1 => bht_20_10_port, A2 => n156, B1 => 
                           bht_21_10_port, B2 => n157, ZN => n267);
   U266 : AOI22_X1 port map( A1 => bht_18_10_port, A2 => n158, B1 => 
                           bht_19_10_port, B2 => n159, ZN => n266);
   U267 : AOI22_X1 port map( A1 => bht_16_10_port, A2 => n160, B1 => 
                           bht_17_10_port, B2 => n161, ZN => n265);
   U268 : NAND4_X1 port map( A1 => n269, A2 => n270, A3 => n271, A4 => n272, ZN
                           => n253);
   U269 : AOI22_X1 port map( A1 => bht_30_10_port, A2 => n142_port, B1 => 
                           bht_31_10_port, B2 => n143_port, ZN => n272);
   U270 : AOI22_X1 port map( A1 => bht_28_10_port, A2 => n144_port, B1 => 
                           bht_29_10_port, B2 => n145_port, ZN => n271);
   U271 : AOI22_X1 port map( A1 => bht_26_10_port, A2 => n146_port, B1 => 
                           bht_27_10_port, B2 => n147_port, ZN => n270);
   U272 : AOI22_X1 port map( A1 => bht_24_10_port, A2 => n148_port, B1 => 
                           bht_25_10_port, B2 => n149_port, ZN => n269);
   U273 : INV_X1 port map( A => n273, ZN => n199);
   U274 : AOI211_X1 port map( C1 => n98, C2 => n190, A => n274, B => n275, ZN 
                           => n273);
   U275 : OAI222_X1 port map( A1 => n276, A2 => n91, B1 => n277, B2 => n95, C1 
                           => n278, C2 => n93, ZN => n275);
   U276 : OAI22_X1 port map( A1 => n279, A2 => n102, B1 => n280, B2 => n100, ZN
                           => n274);
   U277 : INV_X1 port map( A => n281, ZN => n190);
   U278 : OR4_X1 port map( A1 => n282, A2 => n283, A3 => n284, A4 => n285, ZN 
                           => n98);
   U279 : NAND4_X1 port map( A1 => n286, A2 => n287, A3 => n288, A4 => n289, ZN
                           => n285);
   U280 : AOI22_X1 port map( A1 => bht_6_9_port, A2 => n130_port, B1 => 
                           bht_7_9_port, B2 => n131_port, ZN => n289);
   U281 : AOI22_X1 port map( A1 => bht_4_9_port, A2 => n132_port, B1 => 
                           bht_5_9_port, B2 => n133_port, ZN => n288);
   U282 : AOI22_X1 port map( A1 => bht_2_9_port, A2 => n134_port, B1 => 
                           bht_3_9_port, B2 => n135_port, ZN => n287);
   U283 : AOI22_X1 port map( A1 => bht_0_9_port, A2 => n136_port, B1 => 
                           bht_1_9_port, B2 => n137_port, ZN => n286);
   U284 : NAND4_X1 port map( A1 => n290, A2 => n291, A3 => n292, A4 => n293, ZN
                           => n284);
   U285 : AOI22_X1 port map( A1 => bht_14_9_port, A2 => n118, B1 => 
                           bht_15_9_port, B2 => n119, ZN => n293);
   U286 : AOI22_X1 port map( A1 => bht_12_9_port, A2 => n120, B1 => 
                           bht_13_9_port, B2 => n121, ZN => n292);
   U287 : AOI22_X1 port map( A1 => bht_10_9_port, A2 => n122, B1 => 
                           bht_11_9_port, B2 => n123, ZN => n291);
   U288 : AOI22_X1 port map( A1 => bht_8_9_port, A2 => n124, B1 => bht_9_9_port
                           , B2 => n125_port, ZN => n290);
   U289 : NAND4_X1 port map( A1 => n294, A2 => n295, A3 => n296, A4 => n297, ZN
                           => n283);
   U290 : AOI22_X1 port map( A1 => bht_22_9_port, A2 => n154, B1 => 
                           bht_23_9_port, B2 => n155, ZN => n297);
   U291 : AOI22_X1 port map( A1 => bht_20_9_port, A2 => n156, B1 => 
                           bht_21_9_port, B2 => n157, ZN => n296);
   U292 : AOI22_X1 port map( A1 => bht_18_9_port, A2 => n158, B1 => 
                           bht_19_9_port, B2 => n159, ZN => n295);
   U293 : AOI22_X1 port map( A1 => bht_16_9_port, A2 => n160, B1 => 
                           bht_17_9_port, B2 => n161, ZN => n294);
   U294 : NAND4_X1 port map( A1 => n298, A2 => n299, A3 => n300, A4 => n301, ZN
                           => n282);
   U295 : AOI22_X1 port map( A1 => bht_30_9_port, A2 => n142_port, B1 => 
                           bht_31_9_port, B2 => n143_port, ZN => n301);
   U296 : AOI22_X1 port map( A1 => bht_28_9_port, A2 => n144_port, B1 => 
                           bht_29_9_port, B2 => n145_port, ZN => n300);
   U297 : AOI22_X1 port map( A1 => bht_26_9_port, A2 => n146_port, B1 => 
                           bht_27_9_port, B2 => n147_port, ZN => n299);
   U298 : AOI22_X1 port map( A1 => bht_24_9_port, A2 => n148_port, B1 => 
                           bht_25_9_port, B2 => n149_port, ZN => n298);
   U299 : NAND4_X1 port map( A1 => n302, A2 => n303, A3 => n304, A4 => n305, ZN
                           => n198);
   U300 : AOI221_X1 port map( B1 => n306, B2 => n77, C1 => n178, C2 => n76, A 
                           => n307, ZN => n305);
   U301 : OAI22_X1 port map( A1 => n79, A2 => n181, B1 => n81, B2 => n182, ZN 
                           => n307);
   U302 : NOR4_X1 port map( A1 => n308, A2 => n309, A3 => n310, A4 => n311, ZN 
                           => n81);
   U303 : NAND4_X1 port map( A1 => n312, A2 => n313, A3 => n314, A4 => n315, ZN
                           => n311);
   U304 : AOI22_X1 port map( A1 => bht_6_23_port, A2 => n130_port, B1 => 
                           bht_7_23_port, B2 => n131_port, ZN => n315);
   U305 : AOI22_X1 port map( A1 => bht_4_23_port, A2 => n132_port, B1 => 
                           bht_5_23_port, B2 => n133_port, ZN => n314);
   U306 : AOI22_X1 port map( A1 => bht_2_23_port, A2 => n134_port, B1 => 
                           bht_3_23_port, B2 => n135_port, ZN => n313);
   U307 : AOI22_X1 port map( A1 => bht_0_23_port, A2 => n136_port, B1 => 
                           bht_1_23_port, B2 => n137_port, ZN => n312);
   U308 : NAND4_X1 port map( A1 => n316, A2 => n317, A3 => n318, A4 => n319, ZN
                           => n310);
   U309 : AOI22_X1 port map( A1 => bht_14_23_port, A2 => n118, B1 => 
                           bht_15_23_port, B2 => n119, ZN => n319);
   U310 : AOI22_X1 port map( A1 => bht_12_23_port, A2 => n120, B1 => 
                           bht_13_23_port, B2 => n121, ZN => n318);
   U311 : AOI22_X1 port map( A1 => bht_10_23_port, A2 => n122, B1 => 
                           bht_11_23_port, B2 => n123, ZN => n317);
   U312 : AOI22_X1 port map( A1 => bht_8_23_port, A2 => n124, B1 => 
                           bht_9_23_port, B2 => n125_port, ZN => n316);
   U313 : NAND4_X1 port map( A1 => n320, A2 => n321, A3 => n322, A4 => n323, ZN
                           => n309);
   U314 : AOI22_X1 port map( A1 => bht_22_23_port, A2 => n154, B1 => 
                           bht_23_23_port, B2 => n155, ZN => n323);
   U315 : AOI22_X1 port map( A1 => bht_20_23_port, A2 => n156, B1 => 
                           bht_21_23_port, B2 => n157, ZN => n322);
   U316 : AOI22_X1 port map( A1 => bht_18_23_port, A2 => n158, B1 => 
                           bht_19_23_port, B2 => n159, ZN => n321);
   U317 : AOI22_X1 port map( A1 => bht_16_23_port, A2 => n160, B1 => 
                           bht_17_23_port, B2 => n161, ZN => n320);
   U318 : NAND4_X1 port map( A1 => n324, A2 => n325, A3 => n326, A4 => n327, ZN
                           => n308);
   U319 : AOI22_X1 port map( A1 => bht_30_23_port, A2 => n142_port, B1 => 
                           bht_31_23_port, B2 => n143_port, ZN => n327);
   U320 : AOI22_X1 port map( A1 => bht_28_23_port, A2 => n144_port, B1 => 
                           bht_29_23_port, B2 => n145_port, ZN => n326);
   U321 : AOI22_X1 port map( A1 => bht_26_23_port, A2 => n146_port, B1 => 
                           bht_27_23_port, B2 => n147_port, ZN => n325);
   U322 : AOI22_X1 port map( A1 => bht_24_23_port, A2 => n148_port, B1 => 
                           bht_25_23_port, B2 => n149_port, ZN => n324);
   U323 : NOR4_X1 port map( A1 => n328, A2 => n329, A3 => n330, A4 => n331, ZN 
                           => n79);
   U324 : NAND4_X1 port map( A1 => n332, A2 => n333, A3 => n334, A4 => n335, ZN
                           => n331);
   U325 : AOI22_X1 port map( A1 => bht_6_24_port, A2 => n130_port, B1 => 
                           bht_7_24_port, B2 => n131_port, ZN => n335);
   U326 : AOI22_X1 port map( A1 => bht_4_24_port, A2 => n132_port, B1 => 
                           bht_5_24_port, B2 => n133_port, ZN => n334);
   U327 : AOI22_X1 port map( A1 => bht_2_24_port, A2 => n134_port, B1 => 
                           bht_3_24_port, B2 => n135_port, ZN => n333);
   U328 : AOI22_X1 port map( A1 => bht_0_24_port, A2 => n136_port, B1 => 
                           bht_1_24_port, B2 => n137_port, ZN => n332);
   U329 : NAND4_X1 port map( A1 => n336, A2 => n337, A3 => n338, A4 => n339, ZN
                           => n330);
   U330 : AOI22_X1 port map( A1 => bht_14_24_port, A2 => n118, B1 => 
                           bht_15_24_port, B2 => n119, ZN => n339);
   U331 : AOI22_X1 port map( A1 => bht_12_24_port, A2 => n120, B1 => 
                           bht_13_24_port, B2 => n121, ZN => n338);
   U332 : AOI22_X1 port map( A1 => bht_10_24_port, A2 => n122, B1 => 
                           bht_11_24_port, B2 => n123, ZN => n337);
   U333 : AOI22_X1 port map( A1 => bht_8_24_port, A2 => n124, B1 => 
                           bht_9_24_port, B2 => n125_port, ZN => n336);
   U334 : NAND4_X1 port map( A1 => n340, A2 => n341, A3 => n342, A4 => n343, ZN
                           => n329);
   U335 : AOI22_X1 port map( A1 => bht_22_24_port, A2 => n154, B1 => 
                           bht_23_24_port, B2 => n155, ZN => n343);
   U336 : AOI22_X1 port map( A1 => bht_20_24_port, A2 => n156, B1 => 
                           bht_21_24_port, B2 => n157, ZN => n342);
   U337 : AOI22_X1 port map( A1 => bht_18_24_port, A2 => n158, B1 => 
                           bht_19_24_port, B2 => n159, ZN => n341);
   U338 : AOI22_X1 port map( A1 => bht_16_24_port, A2 => n160, B1 => 
                           bht_17_24_port, B2 => n161, ZN => n340);
   U339 : NAND4_X1 port map( A1 => n344, A2 => n345, A3 => n346, A4 => n347, ZN
                           => n328);
   U340 : AOI22_X1 port map( A1 => bht_30_24_port, A2 => n142_port, B1 => 
                           bht_31_24_port, B2 => n143_port, ZN => n347);
   U341 : AOI22_X1 port map( A1 => bht_28_24_port, A2 => n144_port, B1 => 
                           bht_29_24_port, B2 => n145_port, ZN => n346);
   U342 : AOI22_X1 port map( A1 => bht_26_24_port, A2 => n146_port, B1 => 
                           bht_27_24_port, B2 => n147_port, ZN => n345);
   U343 : AOI22_X1 port map( A1 => bht_24_24_port, A2 => n148_port, B1 => 
                           bht_25_24_port, B2 => n149_port, ZN => n344);
   U344 : OR4_X1 port map( A1 => n348, A2 => n349, A3 => n350, A4 => n351, ZN 
                           => n76);
   U345 : NAND4_X1 port map( A1 => n352, A2 => n353, A3 => n354, A4 => n355, ZN
                           => n351);
   U346 : AOI22_X1 port map( A1 => bht_6_26_port, A2 => n130_port, B1 => 
                           bht_7_26_port, B2 => n131_port, ZN => n355);
   U347 : AOI22_X1 port map( A1 => bht_4_26_port, A2 => n132_port, B1 => 
                           bht_5_26_port, B2 => n133_port, ZN => n354);
   U348 : AOI22_X1 port map( A1 => bht_2_26_port, A2 => n134_port, B1 => 
                           bht_3_26_port, B2 => n135_port, ZN => n353);
   U349 : AOI22_X1 port map( A1 => bht_0_26_port, A2 => n136_port, B1 => 
                           bht_1_26_port, B2 => n137_port, ZN => n352);
   U350 : NAND4_X1 port map( A1 => n356, A2 => n357, A3 => n358, A4 => n359, ZN
                           => n350);
   U351 : AOI22_X1 port map( A1 => bht_14_26_port, A2 => n118, B1 => 
                           bht_15_26_port, B2 => n119, ZN => n359);
   U352 : AOI22_X1 port map( A1 => bht_12_26_port, A2 => n120, B1 => 
                           bht_13_26_port, B2 => n121, ZN => n358);
   U353 : AOI22_X1 port map( A1 => bht_10_26_port, A2 => n122, B1 => 
                           bht_11_26_port, B2 => n123, ZN => n357);
   U354 : AOI22_X1 port map( A1 => bht_8_26_port, A2 => n124, B1 => 
                           bht_9_26_port, B2 => n125_port, ZN => n356);
   U355 : NAND4_X1 port map( A1 => n360, A2 => n361, A3 => n362, A4 => n363, ZN
                           => n349);
   U356 : AOI22_X1 port map( A1 => bht_22_26_port, A2 => n154, B1 => 
                           bht_23_26_port, B2 => n155, ZN => n363);
   U357 : AOI22_X1 port map( A1 => bht_20_26_port, A2 => n156, B1 => 
                           bht_21_26_port, B2 => n157, ZN => n362);
   U358 : AOI22_X1 port map( A1 => bht_18_26_port, A2 => n158, B1 => 
                           bht_19_26_port, B2 => n159, ZN => n361);
   U359 : AOI22_X1 port map( A1 => bht_16_26_port, A2 => n160, B1 => 
                           bht_17_26_port, B2 => n161, ZN => n360);
   U360 : NAND4_X1 port map( A1 => n364, A2 => n365, A3 => n366, A4 => n367, ZN
                           => n348);
   U361 : AOI22_X1 port map( A1 => bht_30_26_port, A2 => n142_port, B1 => 
                           bht_31_26_port, B2 => n143_port, ZN => n367);
   U362 : AOI22_X1 port map( A1 => bht_28_26_port, A2 => n144_port, B1 => 
                           bht_29_26_port, B2 => n145_port, ZN => n366);
   U363 : AOI22_X1 port map( A1 => bht_26_26_port, A2 => n146_port, B1 => 
                           bht_27_26_port, B2 => n147_port, ZN => n365);
   U364 : AOI22_X1 port map( A1 => bht_24_26_port, A2 => n148_port, B1 => 
                           bht_25_26_port, B2 => n149_port, ZN => n364);
   U365 : INV_X1 port map( A => n368, ZN => n178);
   U366 : INV_X1 port map( A => n184, ZN => n77);
   U367 : NOR4_X1 port map( A1 => n369, A2 => n370, A3 => n371, A4 => n372, ZN 
                           => n184);
   U368 : NAND4_X1 port map( A1 => n373, A2 => n374, A3 => n375, A4 => n376, ZN
                           => n372);
   U369 : AOI22_X1 port map( A1 => bht_6_25_port, A2 => n130_port, B1 => 
                           bht_7_25_port, B2 => n131_port, ZN => n376);
   U370 : AOI22_X1 port map( A1 => bht_4_25_port, A2 => n132_port, B1 => 
                           bht_5_25_port, B2 => n133_port, ZN => n375);
   U371 : AOI22_X1 port map( A1 => bht_2_25_port, A2 => n134_port, B1 => 
                           bht_3_25_port, B2 => n135_port, ZN => n374);
   U372 : AOI22_X1 port map( A1 => bht_0_25_port, A2 => n136_port, B1 => 
                           bht_1_25_port, B2 => n137_port, ZN => n373);
   U373 : NAND4_X1 port map( A1 => n377, A2 => n378, A3 => n379, A4 => n380, ZN
                           => n371);
   U374 : AOI22_X1 port map( A1 => bht_14_25_port, A2 => n118, B1 => 
                           bht_15_25_port, B2 => n119, ZN => n380);
   U375 : AOI22_X1 port map( A1 => bht_12_25_port, A2 => n120, B1 => 
                           bht_13_25_port, B2 => n121, ZN => n379);
   U376 : AOI22_X1 port map( A1 => bht_10_25_port, A2 => n122, B1 => 
                           bht_11_25_port, B2 => n123, ZN => n378);
   U377 : AOI22_X1 port map( A1 => bht_8_25_port, A2 => n124, B1 => 
                           bht_9_25_port, B2 => n125_port, ZN => n377);
   U378 : NAND4_X1 port map( A1 => n381, A2 => n382, A3 => n383, A4 => n384, ZN
                           => n370);
   U379 : AOI22_X1 port map( A1 => bht_22_25_port, A2 => n154, B1 => 
                           bht_23_25_port, B2 => n155, ZN => n384);
   U380 : AOI22_X1 port map( A1 => bht_20_25_port, A2 => n156, B1 => 
                           bht_21_25_port, B2 => n157, ZN => n383);
   U381 : AOI22_X1 port map( A1 => bht_18_25_port, A2 => n158, B1 => 
                           bht_19_25_port, B2 => n159, ZN => n382);
   U382 : AOI22_X1 port map( A1 => bht_16_25_port, A2 => n160, B1 => 
                           bht_17_25_port, B2 => n161, ZN => n381);
   U383 : NAND4_X1 port map( A1 => n385, A2 => n386, A3 => n387, A4 => n388, ZN
                           => n369);
   U384 : AOI22_X1 port map( A1 => bht_30_25_port, A2 => n142_port, B1 => 
                           bht_31_25_port, B2 => n143_port, ZN => n388);
   U385 : AOI22_X1 port map( A1 => bht_28_25_port, A2 => n144_port, B1 => 
                           bht_29_25_port, B2 => n145_port, ZN => n387);
   U386 : AOI22_X1 port map( A1 => bht_26_25_port, A2 => n146_port, B1 => 
                           bht_27_25_port, B2 => n147_port, ZN => n386);
   U387 : AOI22_X1 port map( A1 => bht_24_25_port, A2 => n148_port, B1 => 
                           bht_25_25_port, B2 => n149_port, ZN => n385);
   U388 : INV_X1 port map( A => n183, ZN => n306);
   U389 : AOI222_X1 port map( A1 => n175, A2 => n83, B1 => n177, B2 => n85, C1 
                           => n179, C2 => n84, ZN => n304);
   U390 : OR4_X1 port map( A1 => n389, A2 => n390, A3 => n391, A4 => n392, ZN 
                           => n84);
   U391 : NAND4_X1 port map( A1 => n393, A2 => n394, A3 => n395, A4 => n396, ZN
                           => n392);
   U392 : AOI22_X1 port map( A1 => bht_6_20_port, A2 => n130_port, B1 => 
                           bht_7_20_port, B2 => n131_port, ZN => n396);
   U393 : AOI22_X1 port map( A1 => bht_4_20_port, A2 => n132_port, B1 => 
                           bht_5_20_port, B2 => n133_port, ZN => n395);
   U394 : AOI22_X1 port map( A1 => bht_2_20_port, A2 => n134_port, B1 => 
                           bht_3_20_port, B2 => n135_port, ZN => n394);
   U395 : AOI22_X1 port map( A1 => bht_0_20_port, A2 => n136_port, B1 => 
                           bht_1_20_port, B2 => n137_port, ZN => n393);
   U396 : NAND4_X1 port map( A1 => n397, A2 => n398, A3 => n399, A4 => n400, ZN
                           => n391);
   U397 : AOI22_X1 port map( A1 => bht_14_20_port, A2 => n118, B1 => 
                           bht_15_20_port, B2 => n119, ZN => n400);
   U398 : AOI22_X1 port map( A1 => bht_12_20_port, A2 => n120, B1 => 
                           bht_13_20_port, B2 => n121, ZN => n399);
   U399 : AOI22_X1 port map( A1 => bht_10_20_port, A2 => n122, B1 => 
                           bht_11_20_port, B2 => n123, ZN => n398);
   U400 : AOI22_X1 port map( A1 => bht_8_20_port, A2 => n124, B1 => 
                           bht_9_20_port, B2 => n125_port, ZN => n397);
   U401 : NAND4_X1 port map( A1 => n401, A2 => n402, A3 => n403, A4 => n404, ZN
                           => n390);
   U402 : AOI22_X1 port map( A1 => bht_22_20_port, A2 => n154, B1 => 
                           bht_23_20_port, B2 => n155, ZN => n404);
   U403 : AOI22_X1 port map( A1 => bht_20_20_port, A2 => n156, B1 => 
                           bht_21_20_port, B2 => n157, ZN => n403);
   U404 : AOI22_X1 port map( A1 => bht_18_20_port, A2 => n158, B1 => 
                           bht_19_20_port, B2 => n159, ZN => n402);
   U405 : AOI22_X1 port map( A1 => bht_16_20_port, A2 => n160, B1 => 
                           bht_17_20_port, B2 => n161, ZN => n401);
   U406 : NAND4_X1 port map( A1 => n405, A2 => n406, A3 => n407, A4 => n408, ZN
                           => n389);
   U407 : AOI22_X1 port map( A1 => bht_30_20_port, A2 => n142_port, B1 => 
                           bht_31_20_port, B2 => n143_port, ZN => n408);
   U408 : AOI22_X1 port map( A1 => bht_28_20_port, A2 => n144_port, B1 => 
                           bht_29_20_port, B2 => n145_port, ZN => n407);
   U409 : AOI22_X1 port map( A1 => bht_26_20_port, A2 => n146_port, B1 => 
                           bht_27_20_port, B2 => n147_port, ZN => n406);
   U410 : AOI22_X1 port map( A1 => bht_24_20_port, A2 => n148_port, B1 => 
                           bht_25_20_port, B2 => n149_port, ZN => n405);
   U411 : INV_X1 port map( A => n409, ZN => n179);
   U412 : OR4_X1 port map( A1 => n410, A2 => n411, A3 => n412, A4 => n413, ZN 
                           => n85);
   U413 : NAND4_X1 port map( A1 => n414, A2 => n415, A3 => n416, A4 => n417, ZN
                           => n413);
   U414 : AOI22_X1 port map( A1 => bht_6_19_port, A2 => n130_port, B1 => 
                           bht_7_19_port, B2 => n131_port, ZN => n417);
   U415 : AOI22_X1 port map( A1 => bht_4_19_port, A2 => n132_port, B1 => 
                           bht_5_19_port, B2 => n133_port, ZN => n416);
   U416 : AOI22_X1 port map( A1 => bht_2_19_port, A2 => n134_port, B1 => 
                           bht_3_19_port, B2 => n135_port, ZN => n415);
   U417 : AOI22_X1 port map( A1 => bht_0_19_port, A2 => n136_port, B1 => 
                           bht_1_19_port, B2 => n137_port, ZN => n414);
   U418 : NAND4_X1 port map( A1 => n418, A2 => n419, A3 => n420, A4 => n421, ZN
                           => n412);
   U419 : AOI22_X1 port map( A1 => bht_14_19_port, A2 => n118, B1 => 
                           bht_15_19_port, B2 => n119, ZN => n421);
   U420 : AOI22_X1 port map( A1 => bht_12_19_port, A2 => n120, B1 => 
                           bht_13_19_port, B2 => n121, ZN => n420);
   U421 : AOI22_X1 port map( A1 => bht_10_19_port, A2 => n122, B1 => 
                           bht_11_19_port, B2 => n123, ZN => n419);
   U422 : AOI22_X1 port map( A1 => bht_8_19_port, A2 => n124, B1 => 
                           bht_9_19_port, B2 => n125_port, ZN => n418);
   U423 : NAND4_X1 port map( A1 => n422, A2 => n423, A3 => n424, A4 => n425, ZN
                           => n411);
   U424 : AOI22_X1 port map( A1 => bht_22_19_port, A2 => n154, B1 => 
                           bht_23_19_port, B2 => n155, ZN => n425);
   U425 : AOI22_X1 port map( A1 => bht_20_19_port, A2 => n156, B1 => 
                           bht_21_19_port, B2 => n157, ZN => n424);
   U426 : AOI22_X1 port map( A1 => bht_18_19_port, A2 => n158, B1 => 
                           bht_19_19_port, B2 => n159, ZN => n423);
   U427 : AOI22_X1 port map( A1 => bht_16_19_port, A2 => n160, B1 => 
                           bht_17_19_port, B2 => n161, ZN => n422);
   U428 : NAND4_X1 port map( A1 => n426, A2 => n427, A3 => n428, A4 => n429, ZN
                           => n410);
   U429 : AOI22_X1 port map( A1 => bht_30_19_port, A2 => n142_port, B1 => 
                           bht_31_19_port, B2 => n143_port, ZN => n429);
   U430 : AOI22_X1 port map( A1 => bht_28_19_port, A2 => n144_port, B1 => 
                           bht_29_19_port, B2 => n145_port, ZN => n428);
   U431 : AOI22_X1 port map( A1 => bht_26_19_port, A2 => n146_port, B1 => 
                           bht_27_19_port, B2 => n147_port, ZN => n427);
   U432 : AOI22_X1 port map( A1 => bht_24_19_port, A2 => n148_port, B1 => 
                           bht_25_19_port, B2 => n149_port, ZN => n426);
   U433 : INV_X1 port map( A => n430, ZN => n177);
   U434 : OR4_X1 port map( A1 => n431, A2 => n432, A3 => n433, A4 => n434, ZN 
                           => n83);
   U435 : NAND4_X1 port map( A1 => n435, A2 => n436, A3 => n437, A4 => n438, ZN
                           => n434);
   U436 : AOI22_X1 port map( A1 => bht_6_21_port, A2 => n130_port, B1 => 
                           bht_7_21_port, B2 => n131_port, ZN => n438);
   U437 : AOI22_X1 port map( A1 => bht_4_21_port, A2 => n132_port, B1 => 
                           bht_5_21_port, B2 => n133_port, ZN => n437);
   U438 : AOI22_X1 port map( A1 => bht_2_21_port, A2 => n134_port, B1 => 
                           bht_3_21_port, B2 => n135_port, ZN => n436);
   U439 : AOI22_X1 port map( A1 => bht_0_21_port, A2 => n136_port, B1 => 
                           bht_1_21_port, B2 => n137_port, ZN => n435);
   U440 : NAND4_X1 port map( A1 => n439, A2 => n440, A3 => n441, A4 => n442, ZN
                           => n433);
   U441 : AOI22_X1 port map( A1 => bht_14_21_port, A2 => n118, B1 => 
                           bht_15_21_port, B2 => n119, ZN => n442);
   U442 : AOI22_X1 port map( A1 => bht_12_21_port, A2 => n120, B1 => 
                           bht_13_21_port, B2 => n121, ZN => n441);
   U443 : AOI22_X1 port map( A1 => bht_10_21_port, A2 => n122, B1 => 
                           bht_11_21_port, B2 => n123, ZN => n440);
   U444 : AOI22_X1 port map( A1 => bht_8_21_port, A2 => n124, B1 => 
                           bht_9_21_port, B2 => n125_port, ZN => n439);
   U445 : NAND4_X1 port map( A1 => n443, A2 => n444, A3 => n445, A4 => n446, ZN
                           => n432);
   U446 : AOI22_X1 port map( A1 => bht_22_21_port, A2 => n154, B1 => 
                           bht_23_21_port, B2 => n155, ZN => n446);
   U447 : AOI22_X1 port map( A1 => bht_20_21_port, A2 => n156, B1 => 
                           bht_21_21_port, B2 => n157, ZN => n445);
   U448 : AOI22_X1 port map( A1 => bht_18_21_port, A2 => n158, B1 => 
                           bht_19_21_port, B2 => n159, ZN => n444);
   U449 : AOI22_X1 port map( A1 => bht_16_21_port, A2 => n160, B1 => 
                           bht_17_21_port, B2 => n161, ZN => n443);
   U450 : NAND4_X1 port map( A1 => n447, A2 => n448, A3 => n449, A4 => n450, ZN
                           => n431);
   U451 : AOI22_X1 port map( A1 => bht_30_21_port, A2 => n142_port, B1 => 
                           bht_31_21_port, B2 => n143_port, ZN => n450);
   U452 : AOI22_X1 port map( A1 => bht_28_21_port, A2 => n144_port, B1 => 
                           bht_29_21_port, B2 => n145_port, ZN => n449);
   U453 : AOI22_X1 port map( A1 => bht_26_21_port, A2 => n146_port, B1 => 
                           bht_27_21_port, B2 => n147_port, ZN => n448);
   U454 : AOI22_X1 port map( A1 => bht_24_21_port, A2 => n148_port, B1 => 
                           bht_25_21_port, B2 => n149_port, ZN => n447);
   U455 : INV_X1 port map( A => n451, ZN => n175);
   U456 : AOI222_X1 port map( A1 => n172, A2 => n88, B1 => n174, B2 => n82, C1 
                           => n176, C2 => n89, ZN => n303);
   U457 : OR4_X1 port map( A1 => n452, A2 => n453, A3 => n454, A4 => n455, ZN 
                           => n89);
   U458 : NAND4_X1 port map( A1 => n456, A2 => n457, A3 => n458, A4 => n459, ZN
                           => n455);
   U459 : AOI22_X1 port map( A1 => bht_6_15_port, A2 => n130_port, B1 => 
                           bht_7_15_port, B2 => n131_port, ZN => n459);
   U460 : AOI22_X1 port map( A1 => bht_4_15_port, A2 => n132_port, B1 => 
                           bht_5_15_port, B2 => n133_port, ZN => n458);
   U461 : AOI22_X1 port map( A1 => bht_2_15_port, A2 => n134_port, B1 => 
                           bht_3_15_port, B2 => n135_port, ZN => n457);
   U462 : AOI22_X1 port map( A1 => bht_0_15_port, A2 => n136_port, B1 => 
                           bht_1_15_port, B2 => n137_port, ZN => n456);
   U463 : NAND4_X1 port map( A1 => n460, A2 => n461, A3 => n462, A4 => n463, ZN
                           => n454);
   U464 : AOI22_X1 port map( A1 => bht_14_15_port, A2 => n118, B1 => 
                           bht_15_15_port, B2 => n119, ZN => n463);
   U465 : AOI22_X1 port map( A1 => bht_12_15_port, A2 => n120, B1 => 
                           bht_13_15_port, B2 => n121, ZN => n462);
   U466 : AOI22_X1 port map( A1 => bht_10_15_port, A2 => n122, B1 => 
                           bht_11_15_port, B2 => n123, ZN => n461);
   U467 : AOI22_X1 port map( A1 => bht_8_15_port, A2 => n124, B1 => 
                           bht_9_15_port, B2 => n125_port, ZN => n460);
   U468 : NAND4_X1 port map( A1 => n464, A2 => n465, A3 => n466, A4 => n467, ZN
                           => n453);
   U469 : AOI22_X1 port map( A1 => bht_22_15_port, A2 => n154, B1 => 
                           bht_23_15_port, B2 => n155, ZN => n467);
   U470 : AOI22_X1 port map( A1 => bht_20_15_port, A2 => n156, B1 => 
                           bht_21_15_port, B2 => n157, ZN => n466);
   U471 : AOI22_X1 port map( A1 => bht_18_15_port, A2 => n158, B1 => 
                           bht_19_15_port, B2 => n159, ZN => n465);
   U472 : AOI22_X1 port map( A1 => bht_16_15_port, A2 => n160, B1 => 
                           bht_17_15_port, B2 => n161, ZN => n464);
   U473 : NAND4_X1 port map( A1 => n468, A2 => n469, A3 => n470, A4 => n471, ZN
                           => n452);
   U474 : AOI22_X1 port map( A1 => bht_30_15_port, A2 => n142_port, B1 => 
                           bht_31_15_port, B2 => n143_port, ZN => n471);
   U475 : AOI22_X1 port map( A1 => bht_28_15_port, A2 => n144_port, B1 => 
                           bht_29_15_port, B2 => n145_port, ZN => n470);
   U476 : AOI22_X1 port map( A1 => bht_26_15_port, A2 => n146_port, B1 => 
                           bht_27_15_port, B2 => n147_port, ZN => n469);
   U477 : AOI22_X1 port map( A1 => bht_24_15_port, A2 => n148_port, B1 => 
                           bht_25_15_port, B2 => n149_port, ZN => n468);
   U478 : INV_X1 port map( A => n472, ZN => n176);
   U479 : OR4_X1 port map( A1 => n473, A2 => n474, A3 => n475, A4 => n476, ZN 
                           => n82);
   U480 : NAND4_X1 port map( A1 => n477, A2 => n478, A3 => n479, A4 => n480, ZN
                           => n476);
   U481 : AOI22_X1 port map( A1 => bht_6_22_port, A2 => n130_port, B1 => 
                           bht_7_22_port, B2 => n131_port, ZN => n480);
   U482 : AOI22_X1 port map( A1 => bht_4_22_port, A2 => n132_port, B1 => 
                           bht_5_22_port, B2 => n133_port, ZN => n479);
   U483 : AOI22_X1 port map( A1 => bht_2_22_port, A2 => n134_port, B1 => 
                           bht_3_22_port, B2 => n135_port, ZN => n478);
   U484 : AOI22_X1 port map( A1 => bht_0_22_port, A2 => n136_port, B1 => 
                           bht_1_22_port, B2 => n137_port, ZN => n477);
   U485 : NAND4_X1 port map( A1 => n481, A2 => n482, A3 => n483, A4 => n484, ZN
                           => n475);
   U486 : AOI22_X1 port map( A1 => bht_14_22_port, A2 => n118, B1 => 
                           bht_15_22_port, B2 => n119, ZN => n484);
   U487 : AOI22_X1 port map( A1 => bht_12_22_port, A2 => n120, B1 => 
                           bht_13_22_port, B2 => n121, ZN => n483);
   U488 : AOI22_X1 port map( A1 => bht_10_22_port, A2 => n122, B1 => 
                           bht_11_22_port, B2 => n123, ZN => n482);
   U489 : AOI22_X1 port map( A1 => bht_8_22_port, A2 => n124, B1 => 
                           bht_9_22_port, B2 => n125_port, ZN => n481);
   U490 : NAND4_X1 port map( A1 => n485, A2 => n486, A3 => n487, A4 => n488, ZN
                           => n474);
   U491 : AOI22_X1 port map( A1 => bht_22_22_port, A2 => n154, B1 => 
                           bht_23_22_port, B2 => n155, ZN => n488);
   U492 : AOI22_X1 port map( A1 => bht_20_22_port, A2 => n156, B1 => 
                           bht_21_22_port, B2 => n157, ZN => n487);
   U493 : AOI22_X1 port map( A1 => bht_18_22_port, A2 => n158, B1 => 
                           bht_19_22_port, B2 => n159, ZN => n486);
   U494 : AOI22_X1 port map( A1 => bht_16_22_port, A2 => n160, B1 => 
                           bht_17_22_port, B2 => n161, ZN => n485);
   U495 : NAND4_X1 port map( A1 => n489, A2 => n490, A3 => n491, A4 => n492, ZN
                           => n473);
   U496 : AOI22_X1 port map( A1 => bht_30_22_port, A2 => n142_port, B1 => 
                           bht_31_22_port, B2 => n143_port, ZN => n492);
   U497 : AOI22_X1 port map( A1 => bht_28_22_port, A2 => n144_port, B1 => 
                           bht_29_22_port, B2 => n145_port, ZN => n491);
   U498 : AOI22_X1 port map( A1 => bht_26_22_port, A2 => n146_port, B1 => 
                           bht_27_22_port, B2 => n147_port, ZN => n490);
   U499 : AOI22_X1 port map( A1 => bht_24_22_port, A2 => n148_port, B1 => 
                           bht_25_22_port, B2 => n149_port, ZN => n489);
   U500 : INV_X1 port map( A => n493, ZN => n174);
   U501 : OR4_X1 port map( A1 => n494, A2 => n495, A3 => n496, A4 => n497, ZN 
                           => n88);
   U502 : NAND4_X1 port map( A1 => n498, A2 => n499, A3 => n500, A4 => n501, ZN
                           => n497);
   U503 : AOI22_X1 port map( A1 => bht_6_16_port, A2 => n130_port, B1 => 
                           bht_7_16_port, B2 => n131_port, ZN => n501);
   U504 : AOI22_X1 port map( A1 => bht_4_16_port, A2 => n132_port, B1 => 
                           bht_5_16_port, B2 => n133_port, ZN => n500);
   U505 : AOI22_X1 port map( A1 => bht_2_16_port, A2 => n134_port, B1 => 
                           bht_3_16_port, B2 => n135_port, ZN => n499);
   U506 : AOI22_X1 port map( A1 => bht_0_16_port, A2 => n136_port, B1 => 
                           bht_1_16_port, B2 => n137_port, ZN => n498);
   U507 : NAND4_X1 port map( A1 => n502, A2 => n503, A3 => n504, A4 => n505, ZN
                           => n496);
   U508 : AOI22_X1 port map( A1 => bht_14_16_port, A2 => n118, B1 => 
                           bht_15_16_port, B2 => n119, ZN => n505);
   U509 : AOI22_X1 port map( A1 => bht_12_16_port, A2 => n120, B1 => 
                           bht_13_16_port, B2 => n121, ZN => n504);
   U510 : AOI22_X1 port map( A1 => bht_10_16_port, A2 => n122, B1 => 
                           bht_11_16_port, B2 => n123, ZN => n503);
   U511 : AOI22_X1 port map( A1 => bht_8_16_port, A2 => n124, B1 => 
                           bht_9_16_port, B2 => n125_port, ZN => n502);
   U512 : NAND4_X1 port map( A1 => n506, A2 => n507, A3 => n508, A4 => n509, ZN
                           => n495);
   U513 : AOI22_X1 port map( A1 => bht_22_16_port, A2 => n154, B1 => 
                           bht_23_16_port, B2 => n155, ZN => n509);
   U514 : AOI22_X1 port map( A1 => bht_20_16_port, A2 => n156, B1 => 
                           bht_21_16_port, B2 => n157, ZN => n508);
   U515 : AOI22_X1 port map( A1 => bht_18_16_port, A2 => n158, B1 => 
                           bht_19_16_port, B2 => n159, ZN => n507);
   U516 : AOI22_X1 port map( A1 => bht_16_16_port, A2 => n160, B1 => 
                           bht_17_16_port, B2 => n161, ZN => n506);
   U517 : NAND4_X1 port map( A1 => n510, A2 => n511, A3 => n512, A4 => n513, ZN
                           => n494);
   U518 : AOI22_X1 port map( A1 => bht_30_16_port, A2 => n142_port, B1 => 
                           bht_31_16_port, B2 => n143_port, ZN => n513);
   U519 : AOI22_X1 port map( A1 => bht_28_16_port, A2 => n144_port, B1 => 
                           bht_29_16_port, B2 => n145_port, ZN => n512);
   U520 : AOI22_X1 port map( A1 => bht_26_16_port, A2 => n146_port, B1 => 
                           bht_27_16_port, B2 => n147_port, ZN => n511);
   U521 : AOI22_X1 port map( A1 => bht_24_16_port, A2 => n148_port, B1 => 
                           bht_25_16_port, B2 => n149_port, ZN => n510);
   U522 : INV_X1 port map( A => n514, ZN => n172);
   U523 : AOI222_X1 port map( A1 => n515, A2 => n96, B1 => n171, B2 => n87, C1 
                           => n173, C2 => n86, ZN => n302);
   U524 : OR4_X1 port map( A1 => n516, A2 => n517, A3 => n518, A4 => n519, ZN 
                           => n86);
   U525 : NAND4_X1 port map( A1 => n520, A2 => n521, A3 => n522, A4 => n523, ZN
                           => n519);
   U526 : AOI22_X1 port map( A1 => bht_6_18_port, A2 => n130_port, B1 => 
                           bht_7_18_port, B2 => n131_port, ZN => n523);
   U527 : AOI22_X1 port map( A1 => bht_4_18_port, A2 => n132_port, B1 => 
                           bht_5_18_port, B2 => n133_port, ZN => n522);
   U528 : AOI22_X1 port map( A1 => bht_2_18_port, A2 => n134_port, B1 => 
                           bht_3_18_port, B2 => n135_port, ZN => n521);
   U529 : AOI22_X1 port map( A1 => bht_0_18_port, A2 => n136_port, B1 => 
                           bht_1_18_port, B2 => n137_port, ZN => n520);
   U530 : NAND4_X1 port map( A1 => n524, A2 => n525, A3 => n526, A4 => n527, ZN
                           => n518);
   U531 : AOI22_X1 port map( A1 => bht_14_18_port, A2 => n118, B1 => 
                           bht_15_18_port, B2 => n119, ZN => n527);
   U532 : AOI22_X1 port map( A1 => bht_12_18_port, A2 => n120, B1 => 
                           bht_13_18_port, B2 => n121, ZN => n526);
   U533 : AOI22_X1 port map( A1 => bht_10_18_port, A2 => n122, B1 => 
                           bht_11_18_port, B2 => n123, ZN => n525);
   U534 : AOI22_X1 port map( A1 => bht_8_18_port, A2 => n124, B1 => 
                           bht_9_18_port, B2 => n125_port, ZN => n524);
   U535 : NAND4_X1 port map( A1 => n528, A2 => n529, A3 => n530, A4 => n531, ZN
                           => n517);
   U536 : AOI22_X1 port map( A1 => bht_22_18_port, A2 => n154, B1 => 
                           bht_23_18_port, B2 => n155, ZN => n531);
   U537 : AOI22_X1 port map( A1 => bht_20_18_port, A2 => n156, B1 => 
                           bht_21_18_port, B2 => n157, ZN => n530);
   U538 : AOI22_X1 port map( A1 => bht_18_18_port, A2 => n158, B1 => 
                           bht_19_18_port, B2 => n159, ZN => n529);
   U539 : AOI22_X1 port map( A1 => bht_16_18_port, A2 => n160, B1 => 
                           bht_17_18_port, B2 => n161, ZN => n528);
   U540 : NAND4_X1 port map( A1 => n532, A2 => n533, A3 => n534, A4 => n535, ZN
                           => n516);
   U541 : AOI22_X1 port map( A1 => bht_30_18_port, A2 => n142_port, B1 => 
                           bht_31_18_port, B2 => n143_port, ZN => n535);
   U542 : AOI22_X1 port map( A1 => bht_28_18_port, A2 => n144_port, B1 => 
                           bht_29_18_port, B2 => n145_port, ZN => n534);
   U543 : AOI22_X1 port map( A1 => bht_26_18_port, A2 => n146_port, B1 => 
                           bht_27_18_port, B2 => n147_port, ZN => n533);
   U544 : AOI22_X1 port map( A1 => bht_24_18_port, A2 => n148_port, B1 => 
                           bht_25_18_port, B2 => n149_port, ZN => n532);
   U545 : INV_X1 port map( A => n536, ZN => n173);
   U546 : OR4_X1 port map( A1 => n537, A2 => n538, A3 => n539, A4 => n540, ZN 
                           => n87);
   U547 : NAND4_X1 port map( A1 => n541, A2 => n542, A3 => n543, A4 => n544, ZN
                           => n540);
   U548 : AOI22_X1 port map( A1 => bht_6_17_port, A2 => n130_port, B1 => 
                           bht_7_17_port, B2 => n131_port, ZN => n544);
   U549 : AOI22_X1 port map( A1 => bht_4_17_port, A2 => n132_port, B1 => 
                           bht_5_17_port, B2 => n133_port, ZN => n543);
   U550 : AOI22_X1 port map( A1 => bht_2_17_port, A2 => n134_port, B1 => 
                           bht_3_17_port, B2 => n135_port, ZN => n542);
   U551 : AOI22_X1 port map( A1 => bht_0_17_port, A2 => n136_port, B1 => 
                           bht_1_17_port, B2 => n137_port, ZN => n541);
   U552 : NAND4_X1 port map( A1 => n545, A2 => n546, A3 => n547, A4 => n548, ZN
                           => n539);
   U553 : AOI22_X1 port map( A1 => bht_14_17_port, A2 => n118, B1 => 
                           bht_15_17_port, B2 => n119, ZN => n548);
   U554 : AOI22_X1 port map( A1 => bht_12_17_port, A2 => n120, B1 => 
                           bht_13_17_port, B2 => n121, ZN => n547);
   U555 : AOI22_X1 port map( A1 => bht_10_17_port, A2 => n122, B1 => 
                           bht_11_17_port, B2 => n123, ZN => n546);
   U556 : AOI22_X1 port map( A1 => bht_8_17_port, A2 => n124, B1 => 
                           bht_9_17_port, B2 => n125_port, ZN => n545);
   U557 : NAND4_X1 port map( A1 => n549, A2 => n550, A3 => n551, A4 => n552, ZN
                           => n538);
   U558 : AOI22_X1 port map( A1 => bht_22_17_port, A2 => n154, B1 => 
                           bht_23_17_port, B2 => n155, ZN => n552);
   U559 : AOI22_X1 port map( A1 => bht_20_17_port, A2 => n156, B1 => 
                           bht_21_17_port, B2 => n157, ZN => n551);
   U560 : AOI22_X1 port map( A1 => bht_18_17_port, A2 => n158, B1 => 
                           bht_19_17_port, B2 => n159, ZN => n550);
   U561 : AOI22_X1 port map( A1 => bht_16_17_port, A2 => n160, B1 => 
                           bht_17_17_port, B2 => n161, ZN => n549);
   U562 : NAND4_X1 port map( A1 => n553, A2 => n554, A3 => n555, A4 => n556, ZN
                           => n537);
   U563 : AOI22_X1 port map( A1 => bht_30_17_port, A2 => n142_port, B1 => 
                           bht_31_17_port, B2 => n143_port, ZN => n556);
   U564 : AOI22_X1 port map( A1 => bht_28_17_port, A2 => n144_port, B1 => 
                           bht_29_17_port, B2 => n145_port, ZN => n555);
   U565 : AOI22_X1 port map( A1 => bht_26_17_port, A2 => n146_port, B1 => 
                           bht_27_17_port, B2 => n147_port, ZN => n554);
   U566 : AOI22_X1 port map( A1 => bht_24_17_port, A2 => n148_port, B1 => 
                           bht_25_17_port, B2 => n149_port, ZN => n553);
   U567 : INV_X1 port map( A => n557, ZN => n171);
   U568 : INV_X1 port map( A => n558, ZN => n96);
   U569 : INV_X1 port map( A => n559, ZN => n515);
   U570 : NOR2_X1 port map( A1 => n560, A2 => n561, ZN => n196);
   U571 : NAND4_X1 port map( A1 => n562, A2 => n563, A3 => n564, A4 => n565, ZN
                           => n561);
   U572 : NOR4_X1 port map( A1 => n493, A2 => n536, A3 => n514, A4 => n557, ZN 
                           => n565);
   U573 : MUX2_X1 port map( A => reg_a(15), B => addr(22), S => sig_bal, Z => 
                           n557);
   U574 : MUX2_X1 port map( A => reg_a(14), B => addr(21), S => sig_bal, Z => 
                           n514);
   U575 : MUX2_X1 port map( A => reg_a(16), B => addr(23), S => sig_bal, Z => 
                           n536);
   U576 : MUX2_X1 port map( A => reg_a(20), B => addr(27), S => sig_bal, Z => 
                           n493);
   U577 : NOR4_X1 port map( A1 => n278, A2 => n559, A3 => n277, A4 => n280, ZN 
                           => n564);
   U578 : NOR4_X1 port map( A1 => n276, A2 => n279, A3 => n185, A4 => n281, ZN 
                           => n563);
   U579 : MUX2_X1 port map( A => reg_a(7), B => addr(14), S => sig_bal, Z => 
                           n281);
   U580 : NOR4_X1 port map( A1 => n192, A2 => n252, A3 => reg_a(1), A4 => n205,
                           ZN => n562);
   U581 : MUX2_X1 port map( A => reg_a(8), B => addr(15), S => sig_bal, Z => 
                           n192);
   U582 : NAND4_X1 port map( A1 => n566, A2 => n567, A3 => n568, A4 => n569, ZN
                           => n560);
   U583 : NOR4_X1 port map( A1 => reg_a(31), A2 => reg_a(30), A3 => reg_a(29), 
                           A4 => reg_a(28), ZN => n569);
   U584 : NOR4_X1 port map( A1 => reg_a(27), A2 => reg_a(26), A3 => reg_a(25), 
                           A4 => reg_a(0), ZN => n568);
   U585 : NOR4_X1 port map( A1 => n183, A2 => n182, A3 => n181, A4 => n409, ZN 
                           => n567);
   U586 : MUX2_X1 port map( A => reg_a(18), B => addr(25), S => sig_bal, Z => 
                           n409);
   U587 : MUX2_X1 port map( A => reg_a(22), B => addr(29), S => sig_bal, Z => 
                           n181);
   U588 : MUX2_X1 port map( A => reg_a(21), B => addr(28), S => sig_bal, Z => 
                           n182);
   U589 : MUX2_X1 port map( A => reg_a(23), B => addr(30), S => sig_bal, Z => 
                           n183);
   U590 : NOR4_X1 port map( A1 => n368, A2 => n430, A3 => n472, A4 => n451, ZN 
                           => n566);
   U591 : MUX2_X1 port map( A => reg_a(19), B => addr(26), S => sig_bal, Z => 
                           n451);
   U592 : MUX2_X1 port map( A => reg_a(13), B => addr(20), S => sig_bal, Z => 
                           n472);
   U593 : MUX2_X1 port map( A => reg_a(17), B => addr(24), S => sig_bal, Z => 
                           n430);
   U594 : MUX2_X1 port map( A => reg_a(24), B => addr(31), S => sig_bal, Z => 
                           n368);
   U595 : INV_X1 port map( A => n204, ZN => n103);
   U596 : NOR4_X1 port map( A1 => n570, A2 => n571, A3 => n572, A4 => n573, ZN 
                           => n204);
   U597 : NAND4_X1 port map( A1 => n574, A2 => n575, A3 => n576, A4 => n577, ZN
                           => n573);
   U598 : AOI22_X1 port map( A1 => bht_6_6_port, A2 => n130_port, B1 => 
                           bht_7_6_port, B2 => n131_port, ZN => n577);
   U599 : AOI22_X1 port map( A1 => bht_4_6_port, A2 => n132_port, B1 => 
                           bht_5_6_port, B2 => n133_port, ZN => n576);
   U600 : AOI22_X1 port map( A1 => bht_2_6_port, A2 => n134_port, B1 => 
                           bht_3_6_port, B2 => n135_port, ZN => n575);
   U601 : AOI22_X1 port map( A1 => bht_0_6_port, A2 => n136_port, B1 => 
                           bht_1_6_port, B2 => n137_port, ZN => n574);
   U602 : NAND4_X1 port map( A1 => n578, A2 => n579, A3 => n580, A4 => n581, ZN
                           => n572);
   U603 : AOI22_X1 port map( A1 => bht_14_6_port, A2 => n118, B1 => 
                           bht_15_6_port, B2 => n119, ZN => n581);
   U604 : AOI22_X1 port map( A1 => bht_12_6_port, A2 => n120, B1 => 
                           bht_13_6_port, B2 => n121, ZN => n580);
   U605 : AOI22_X1 port map( A1 => bht_10_6_port, A2 => n122, B1 => 
                           bht_11_6_port, B2 => n123, ZN => n579);
   U606 : AOI22_X1 port map( A1 => bht_8_6_port, A2 => n124, B1 => bht_9_6_port
                           , B2 => n125_port, ZN => n578);
   U607 : NAND4_X1 port map( A1 => n582, A2 => n583, A3 => n584, A4 => n585, ZN
                           => n571);
   U608 : AOI22_X1 port map( A1 => bht_22_6_port, A2 => n154, B1 => 
                           bht_23_6_port, B2 => n155, ZN => n585);
   U609 : AOI22_X1 port map( A1 => bht_20_6_port, A2 => n156, B1 => 
                           bht_21_6_port, B2 => n157, ZN => n584);
   U610 : AOI22_X1 port map( A1 => bht_18_6_port, A2 => n158, B1 => 
                           bht_19_6_port, B2 => n159, ZN => n583);
   U611 : AOI22_X1 port map( A1 => bht_16_6_port, A2 => n160, B1 => 
                           bht_17_6_port, B2 => n161, ZN => n582);
   U612 : NAND4_X1 port map( A1 => n586, A2 => n587, A3 => n588, A4 => n589, ZN
                           => n570);
   U613 : AOI22_X1 port map( A1 => bht_30_6_port, A2 => n142_port, B1 => 
                           bht_31_6_port, B2 => n143_port, ZN => n589);
   U614 : AOI22_X1 port map( A1 => bht_28_6_port, A2 => n144_port, B1 => 
                           bht_29_6_port, B2 => n145_port, ZN => n588);
   U615 : AOI22_X1 port map( A1 => bht_26_6_port, A2 => n146_port, B1 => 
                           bht_27_6_port, B2 => n147_port, ZN => n587);
   U616 : AOI22_X1 port map( A1 => bht_24_6_port, A2 => n148_port, B1 => 
                           bht_25_6_port, B2 => n149_port, ZN => n586);
   U617 : INV_X1 port map( A => n205, ZN => n194);
   U618 : MUX2_X1 port map( A => reg_a(4), B => addr(11), S => sig_bal, Z => 
                           n205);
   U619 : INV_X1 port map( A => n251, ZN => n104);
   U620 : NOR4_X1 port map( A1 => n590, A2 => n591, A3 => n592, A4 => n593, ZN 
                           => n251);
   U621 : NAND4_X1 port map( A1 => n594, A2 => n595, A3 => n596, A4 => n597, ZN
                           => n593);
   U622 : AOI22_X1 port map( A1 => bht_6_5_port, A2 => n130_port, B1 => 
                           bht_7_5_port, B2 => n131_port, ZN => n597);
   U623 : AOI22_X1 port map( A1 => bht_4_5_port, A2 => n132_port, B1 => 
                           bht_5_5_port, B2 => n133_port, ZN => n596);
   U624 : AOI22_X1 port map( A1 => bht_2_5_port, A2 => n134_port, B1 => 
                           bht_3_5_port, B2 => n135_port, ZN => n595);
   U625 : AOI22_X1 port map( A1 => bht_0_5_port, A2 => n136_port, B1 => 
                           bht_1_5_port, B2 => n137_port, ZN => n594);
   U626 : NAND4_X1 port map( A1 => n598, A2 => n599, A3 => n600, A4 => n601, ZN
                           => n592);
   U627 : AOI22_X1 port map( A1 => bht_14_5_port, A2 => n118, B1 => 
                           bht_15_5_port, B2 => n119, ZN => n601);
   U628 : AOI22_X1 port map( A1 => bht_12_5_port, A2 => n120, B1 => 
                           bht_13_5_port, B2 => n121, ZN => n600);
   U629 : AOI22_X1 port map( A1 => bht_10_5_port, A2 => n122, B1 => 
                           bht_11_5_port, B2 => n123, ZN => n599);
   U630 : AOI22_X1 port map( A1 => bht_8_5_port, A2 => n124, B1 => bht_9_5_port
                           , B2 => n125_port, ZN => n598);
   U631 : NAND4_X1 port map( A1 => n602, A2 => n603, A3 => n604, A4 => n605, ZN
                           => n591);
   U632 : AOI22_X1 port map( A1 => bht_22_5_port, A2 => n154, B1 => 
                           bht_23_5_port, B2 => n155, ZN => n605);
   U633 : AOI22_X1 port map( A1 => bht_20_5_port, A2 => n156, B1 => 
                           bht_21_5_port, B2 => n157, ZN => n604);
   U634 : AOI22_X1 port map( A1 => bht_18_5_port, A2 => n158, B1 => 
                           bht_19_5_port, B2 => n159, ZN => n603);
   U635 : AOI22_X1 port map( A1 => bht_16_5_port, A2 => n160, B1 => 
                           bht_17_5_port, B2 => n161, ZN => n602);
   U636 : NAND4_X1 port map( A1 => n606, A2 => n607, A3 => n608, A4 => n609, ZN
                           => n590);
   U637 : AOI22_X1 port map( A1 => bht_30_5_port, A2 => n142_port, B1 => 
                           bht_31_5_port, B2 => n143_port, ZN => n609);
   U638 : AOI22_X1 port map( A1 => bht_28_5_port, A2 => n144_port, B1 => 
                           bht_29_5_port, B2 => n145_port, ZN => n608);
   U639 : AOI22_X1 port map( A1 => bht_26_5_port, A2 => n146_port, B1 => 
                           bht_27_5_port, B2 => n147_port, ZN => n607);
   U640 : AOI22_X1 port map( A1 => bht_24_5_port, A2 => n148_port, B1 => 
                           bht_25_5_port, B2 => n149_port, ZN => n606);
   U641 : INV_X1 port map( A => n252, ZN => n193);
   U642 : MUX2_X1 port map( A => reg_a(3), B => addr(10), S => sig_bal, Z => 
                           n252);
   U643 : MUX2_X1 port map( A => reg_a(2), B => addr(9), S => sig_bal, Z => 
                           n185);
   U644 : NOR4_X1 port map( A1 => n610, A2 => n611, A3 => n612, A4 => n613, ZN 
                           => n106);
   U645 : NAND4_X1 port map( A1 => n614, A2 => n615, A3 => n616, A4 => n617, ZN
                           => n613);
   U646 : AOI22_X1 port map( A1 => bht_6_4_port, A2 => n130_port, B1 => 
                           bht_7_4_port, B2 => n131_port, ZN => n617);
   U647 : AOI22_X1 port map( A1 => bht_4_4_port, A2 => n132_port, B1 => 
                           bht_5_4_port, B2 => n133_port, ZN => n616);
   U648 : AOI22_X1 port map( A1 => bht_2_4_port, A2 => n134_port, B1 => 
                           bht_3_4_port, B2 => n135_port, ZN => n615);
   U649 : AOI22_X1 port map( A1 => bht_0_4_port, A2 => n136_port, B1 => 
                           bht_1_4_port, B2 => n137_port, ZN => n614);
   U650 : NAND4_X1 port map( A1 => n618, A2 => n619, A3 => n620, A4 => n621, ZN
                           => n612);
   U651 : AOI22_X1 port map( A1 => bht_14_4_port, A2 => n118, B1 => 
                           bht_15_4_port, B2 => n119, ZN => n621);
   U652 : AOI22_X1 port map( A1 => bht_12_4_port, A2 => n120, B1 => 
                           bht_13_4_port, B2 => n121, ZN => n620);
   U653 : AOI22_X1 port map( A1 => bht_10_4_port, A2 => n122, B1 => 
                           bht_11_4_port, B2 => n123, ZN => n619);
   U654 : AOI22_X1 port map( A1 => bht_8_4_port, A2 => n124, B1 => bht_9_4_port
                           , B2 => n125_port, ZN => n618);
   U655 : NAND4_X1 port map( A1 => n622, A2 => n623, A3 => n624, A4 => n625, ZN
                           => n611);
   U656 : AOI22_X1 port map( A1 => bht_22_4_port, A2 => n154, B1 => 
                           bht_23_4_port, B2 => n155, ZN => n625);
   U657 : AOI22_X1 port map( A1 => bht_20_4_port, A2 => n156, B1 => 
                           bht_21_4_port, B2 => n157, ZN => n624);
   U658 : AOI22_X1 port map( A1 => bht_18_4_port, A2 => n158, B1 => 
                           bht_19_4_port, B2 => n159, ZN => n623);
   U659 : AOI22_X1 port map( A1 => bht_16_4_port, A2 => n160, B1 => 
                           bht_17_4_port, B2 => n161, ZN => n622);
   U660 : NAND4_X1 port map( A1 => n626, A2 => n627, A3 => n628, A4 => n629, ZN
                           => n610);
   U661 : AOI22_X1 port map( A1 => bht_30_4_port, A2 => n142_port, B1 => 
                           bht_31_4_port, B2 => n143_port, ZN => n629);
   U662 : AOI22_X1 port map( A1 => bht_28_4_port, A2 => n144_port, B1 => 
                           bht_29_4_port, B2 => n145_port, ZN => n628);
   U663 : AOI22_X1 port map( A1 => bht_26_4_port, A2 => n146_port, B1 => 
                           bht_27_4_port, B2 => n147_port, ZN => n627);
   U664 : AOI22_X1 port map( A1 => bht_24_4_port, A2 => n148_port, B1 => 
                           bht_25_4_port, B2 => n149_port, ZN => n626);
   U665 : AOI222_X1 port map( A1 => n93, A2 => n278, B1 => n558, B2 => n559, C1
                           => n95, C2 => n277, ZN => n164);
   U666 : MUX2_X1 port map( A => reg_a(10), B => addr(17), S => sig_bal, Z => 
                           n277);
   U667 : NOR4_X1 port map( A1 => n630, A2 => n631, A3 => n632, A4 => n633, ZN 
                           => n95);
   U668 : NAND4_X1 port map( A1 => n634, A2 => n635, A3 => n636, A4 => n637, ZN
                           => n633);
   U669 : AOI22_X1 port map( A1 => bht_6_12_port, A2 => n130_port, B1 => 
                           bht_7_12_port, B2 => n131_port, ZN => n637);
   U670 : AOI22_X1 port map( A1 => bht_4_12_port, A2 => n132_port, B1 => 
                           bht_5_12_port, B2 => n133_port, ZN => n636);
   U671 : AOI22_X1 port map( A1 => bht_2_12_port, A2 => n134_port, B1 => 
                           bht_3_12_port, B2 => n135_port, ZN => n635);
   U672 : AOI22_X1 port map( A1 => bht_0_12_port, A2 => n136_port, B1 => 
                           bht_1_12_port, B2 => n137_port, ZN => n634);
   U673 : NAND4_X1 port map( A1 => n638, A2 => n639, A3 => n640, A4 => n641, ZN
                           => n632);
   U674 : AOI22_X1 port map( A1 => bht_14_12_port, A2 => n118, B1 => 
                           bht_15_12_port, B2 => n119, ZN => n641);
   U675 : AOI22_X1 port map( A1 => bht_12_12_port, A2 => n120, B1 => 
                           bht_13_12_port, B2 => n121, ZN => n640);
   U676 : AOI22_X1 port map( A1 => bht_10_12_port, A2 => n122, B1 => 
                           bht_11_12_port, B2 => n123, ZN => n639);
   U677 : AOI22_X1 port map( A1 => bht_8_12_port, A2 => n124, B1 => 
                           bht_9_12_port, B2 => n125_port, ZN => n638);
   U678 : NAND4_X1 port map( A1 => n642, A2 => n643, A3 => n644, A4 => n645, ZN
                           => n631);
   U679 : AOI22_X1 port map( A1 => bht_22_12_port, A2 => n154, B1 => 
                           bht_23_12_port, B2 => n155, ZN => n645);
   U680 : AOI22_X1 port map( A1 => bht_20_12_port, A2 => n156, B1 => 
                           bht_21_12_port, B2 => n157, ZN => n644);
   U681 : AOI22_X1 port map( A1 => bht_18_12_port, A2 => n158, B1 => 
                           bht_19_12_port, B2 => n159, ZN => n643);
   U682 : AOI22_X1 port map( A1 => bht_16_12_port, A2 => n160, B1 => 
                           bht_17_12_port, B2 => n161, ZN => n642);
   U683 : NAND4_X1 port map( A1 => n646, A2 => n647, A3 => n648, A4 => n649, ZN
                           => n630);
   U684 : AOI22_X1 port map( A1 => bht_30_12_port, A2 => n142_port, B1 => 
                           bht_31_12_port, B2 => n143_port, ZN => n649);
   U685 : AOI22_X1 port map( A1 => bht_28_12_port, A2 => n144_port, B1 => 
                           bht_29_12_port, B2 => n145_port, ZN => n648);
   U686 : AOI22_X1 port map( A1 => bht_26_12_port, A2 => n146_port, B1 => 
                           bht_27_12_port, B2 => n147_port, ZN => n647);
   U687 : AOI22_X1 port map( A1 => bht_24_12_port, A2 => n148_port, B1 => 
                           bht_25_12_port, B2 => n149_port, ZN => n646);
   U688 : MUX2_X1 port map( A => reg_a(9), B => addr(16), S => sig_bal, Z => 
                           n559);
   U689 : NOR4_X1 port map( A1 => n650, A2 => n651, A3 => n652, A4 => n653, ZN 
                           => n558);
   U690 : NAND4_X1 port map( A1 => n654, A2 => n655, A3 => n656, A4 => n657, ZN
                           => n653);
   U691 : AOI22_X1 port map( A1 => bht_6_11_port, A2 => n130_port, B1 => 
                           bht_7_11_port, B2 => n131_port, ZN => n657);
   U692 : AOI22_X1 port map( A1 => bht_4_11_port, A2 => n132_port, B1 => 
                           bht_5_11_port, B2 => n133_port, ZN => n656);
   U693 : AOI22_X1 port map( A1 => bht_2_11_port, A2 => n134_port, B1 => 
                           bht_3_11_port, B2 => n135_port, ZN => n655);
   U694 : AOI22_X1 port map( A1 => bht_0_11_port, A2 => n136_port, B1 => 
                           bht_1_11_port, B2 => n137_port, ZN => n654);
   U695 : NAND4_X1 port map( A1 => n658, A2 => n659, A3 => n660, A4 => n661, ZN
                           => n652);
   U696 : AOI22_X1 port map( A1 => bht_14_11_port, A2 => n118, B1 => 
                           bht_15_11_port, B2 => n119, ZN => n661);
   U697 : AOI22_X1 port map( A1 => bht_12_11_port, A2 => n120, B1 => 
                           bht_13_11_port, B2 => n121, ZN => n660);
   U698 : AOI22_X1 port map( A1 => bht_10_11_port, A2 => n122, B1 => 
                           bht_11_11_port, B2 => n123, ZN => n659);
   U699 : AOI22_X1 port map( A1 => bht_8_11_port, A2 => n124, B1 => 
                           bht_9_11_port, B2 => n125_port, ZN => n658);
   U700 : NAND4_X1 port map( A1 => n662, A2 => n663, A3 => n664, A4 => n665, ZN
                           => n651);
   U701 : AOI22_X1 port map( A1 => bht_22_11_port, A2 => n154, B1 => 
                           bht_23_11_port, B2 => n155, ZN => n665);
   U702 : AOI22_X1 port map( A1 => bht_20_11_port, A2 => n156, B1 => 
                           bht_21_11_port, B2 => n157, ZN => n664);
   U703 : AOI22_X1 port map( A1 => bht_18_11_port, A2 => n158, B1 => 
                           bht_19_11_port, B2 => n159, ZN => n663);
   U704 : AOI22_X1 port map( A1 => bht_16_11_port, A2 => n160, B1 => 
                           bht_17_11_port, B2 => n161, ZN => n662);
   U705 : NAND4_X1 port map( A1 => n666, A2 => n667, A3 => n668, A4 => n669, ZN
                           => n650);
   U706 : AOI22_X1 port map( A1 => bht_30_11_port, A2 => n142_port, B1 => 
                           bht_31_11_port, B2 => n143_port, ZN => n669);
   U707 : AOI22_X1 port map( A1 => bht_28_11_port, A2 => n144_port, B1 => 
                           bht_29_11_port, B2 => n145_port, ZN => n668);
   U708 : AOI22_X1 port map( A1 => bht_26_11_port, A2 => n146_port, B1 => 
                           bht_27_11_port, B2 => n147_port, ZN => n667);
   U709 : AOI22_X1 port map( A1 => bht_24_11_port, A2 => n148_port, B1 => 
                           bht_25_11_port, B2 => n149_port, ZN => n666);
   U710 : MUX2_X1 port map( A => reg_a(11), B => addr(18), S => sig_bal, Z => 
                           n278);
   U711 : NOR4_X1 port map( A1 => n670, A2 => n671, A3 => n672, A4 => n673, ZN 
                           => n93);
   U712 : NAND4_X1 port map( A1 => n674, A2 => n675, A3 => n676, A4 => n677, ZN
                           => n673);
   U713 : AOI22_X1 port map( A1 => bht_6_13_port, A2 => n130_port, B1 => 
                           bht_7_13_port, B2 => n131_port, ZN => n677);
   U714 : AOI22_X1 port map( A1 => bht_4_13_port, A2 => n132_port, B1 => 
                           bht_5_13_port, B2 => n133_port, ZN => n676);
   U715 : AOI22_X1 port map( A1 => bht_2_13_port, A2 => n134_port, B1 => 
                           bht_3_13_port, B2 => n135_port, ZN => n675);
   U716 : AOI22_X1 port map( A1 => bht_0_13_port, A2 => n136_port, B1 => 
                           bht_1_13_port, B2 => n137_port, ZN => n674);
   U717 : NAND4_X1 port map( A1 => n678, A2 => n679, A3 => n680, A4 => n681, ZN
                           => n672);
   U718 : AOI22_X1 port map( A1 => bht_14_13_port, A2 => n118, B1 => 
                           bht_15_13_port, B2 => n119, ZN => n681);
   U719 : AOI22_X1 port map( A1 => bht_12_13_port, A2 => n120, B1 => 
                           bht_13_13_port, B2 => n121, ZN => n680);
   U720 : AOI22_X1 port map( A1 => bht_10_13_port, A2 => n122, B1 => 
                           bht_11_13_port, B2 => n123, ZN => n679);
   U721 : AOI22_X1 port map( A1 => bht_8_13_port, A2 => n124, B1 => 
                           bht_9_13_port, B2 => n125_port, ZN => n678);
   U722 : NAND4_X1 port map( A1 => n682, A2 => n683, A3 => n684, A4 => n685, ZN
                           => n671);
   U723 : AOI22_X1 port map( A1 => bht_22_13_port, A2 => n154, B1 => 
                           bht_23_13_port, B2 => n155, ZN => n685);
   U724 : AOI22_X1 port map( A1 => bht_20_13_port, A2 => n156, B1 => 
                           bht_21_13_port, B2 => n157, ZN => n684);
   U725 : AOI22_X1 port map( A1 => bht_18_13_port, A2 => n158, B1 => 
                           bht_19_13_port, B2 => n159, ZN => n683);
   U726 : AOI22_X1 port map( A1 => bht_16_13_port, A2 => n160, B1 => 
                           bht_17_13_port, B2 => n161, ZN => n682);
   U727 : NAND4_X1 port map( A1 => n686, A2 => n687, A3 => n688, A4 => n689, ZN
                           => n670);
   U728 : AOI22_X1 port map( A1 => bht_30_13_port, A2 => n142_port, B1 => 
                           bht_31_13_port, B2 => n143_port, ZN => n689);
   U729 : AOI22_X1 port map( A1 => bht_28_13_port, A2 => n144_port, B1 => 
                           bht_29_13_port, B2 => n145_port, ZN => n688);
   U730 : AOI22_X1 port map( A1 => bht_26_13_port, A2 => n146_port, B1 => 
                           bht_27_13_port, B2 => n147_port, ZN => n687);
   U731 : AOI22_X1 port map( A1 => bht_24_13_port, A2 => n148_port, B1 => 
                           bht_25_13_port, B2 => n149_port, ZN => n686);
   U732 : AOI222_X1 port map( A1 => n100, A2 => n280, B1 => n91, B2 => n276, C1
                           => n102, C2 => n279, ZN => n163);
   U733 : MUX2_X1 port map( A => reg_a(5), B => addr(12), S => sig_bal, Z => 
                           n279);
   U734 : NOR4_X1 port map( A1 => n690, A2 => n691, A3 => n692, A4 => n693, ZN 
                           => n102);
   U735 : NAND4_X1 port map( A1 => n694, A2 => n695, A3 => n696, A4 => n697, ZN
                           => n693);
   U736 : AOI22_X1 port map( A1 => bht_6_7_port, A2 => n130_port, B1 => 
                           bht_7_7_port, B2 => n131_port, ZN => n697);
   U737 : AOI22_X1 port map( A1 => bht_4_7_port, A2 => n132_port, B1 => 
                           bht_5_7_port, B2 => n133_port, ZN => n696);
   U738 : AOI22_X1 port map( A1 => bht_2_7_port, A2 => n134_port, B1 => 
                           bht_3_7_port, B2 => n135_port, ZN => n695);
   U739 : AOI22_X1 port map( A1 => bht_0_7_port, A2 => n136_port, B1 => 
                           bht_1_7_port, B2 => n137_port, ZN => n694);
   U740 : NAND4_X1 port map( A1 => n698, A2 => n699, A3 => n700, A4 => n701, ZN
                           => n692);
   U741 : AOI22_X1 port map( A1 => bht_14_7_port, A2 => n118, B1 => 
                           bht_15_7_port, B2 => n119, ZN => n701);
   U742 : AOI22_X1 port map( A1 => bht_12_7_port, A2 => n120, B1 => 
                           bht_13_7_port, B2 => n121, ZN => n700);
   U743 : AOI22_X1 port map( A1 => bht_10_7_port, A2 => n122, B1 => 
                           bht_11_7_port, B2 => n123, ZN => n699);
   U744 : AOI22_X1 port map( A1 => bht_8_7_port, A2 => n124, B1 => bht_9_7_port
                           , B2 => n125_port, ZN => n698);
   U745 : NAND4_X1 port map( A1 => n702, A2 => n703, A3 => n704, A4 => n705, ZN
                           => n691);
   U746 : AOI22_X1 port map( A1 => bht_22_7_port, A2 => n154, B1 => 
                           bht_23_7_port, B2 => n155, ZN => n705);
   U747 : AOI22_X1 port map( A1 => bht_20_7_port, A2 => n156, B1 => 
                           bht_21_7_port, B2 => n157, ZN => n704);
   U748 : AOI22_X1 port map( A1 => bht_18_7_port, A2 => n158, B1 => 
                           bht_19_7_port, B2 => n159, ZN => n703);
   U749 : AOI22_X1 port map( A1 => bht_16_7_port, A2 => n160, B1 => 
                           bht_17_7_port, B2 => n161, ZN => n702);
   U750 : NAND4_X1 port map( A1 => n706, A2 => n707, A3 => n708, A4 => n709, ZN
                           => n690);
   U751 : AOI22_X1 port map( A1 => bht_30_7_port, A2 => n142_port, B1 => 
                           bht_31_7_port, B2 => n143_port, ZN => n709);
   U752 : AOI22_X1 port map( A1 => bht_28_7_port, A2 => n144_port, B1 => 
                           bht_29_7_port, B2 => n145_port, ZN => n708);
   U753 : AOI22_X1 port map( A1 => bht_26_7_port, A2 => n146_port, B1 => 
                           bht_27_7_port, B2 => n147_port, ZN => n707);
   U754 : AOI22_X1 port map( A1 => bht_24_7_port, A2 => n148_port, B1 => 
                           bht_25_7_port, B2 => n149_port, ZN => n706);
   U755 : MUX2_X1 port map( A => reg_a(12), B => addr(19), S => sig_bal, Z => 
                           n276);
   U756 : NOR4_X1 port map( A1 => n710, A2 => n711, A3 => n712, A4 => n713, ZN 
                           => n91);
   U757 : NAND4_X1 port map( A1 => n714, A2 => n715, A3 => n716, A4 => n717, ZN
                           => n713);
   U758 : AOI22_X1 port map( A1 => bht_6_14_port, A2 => n130_port, B1 => 
                           bht_7_14_port, B2 => n131_port, ZN => n717);
   U759 : AOI22_X1 port map( A1 => bht_4_14_port, A2 => n132_port, B1 => 
                           bht_5_14_port, B2 => n133_port, ZN => n716);
   U760 : AOI22_X1 port map( A1 => bht_2_14_port, A2 => n134_port, B1 => 
                           bht_3_14_port, B2 => n135_port, ZN => n715);
   U761 : AOI22_X1 port map( A1 => bht_0_14_port, A2 => n136_port, B1 => 
                           bht_1_14_port, B2 => n137_port, ZN => n714);
   U762 : NAND4_X1 port map( A1 => n718, A2 => n719, A3 => n720, A4 => n721, ZN
                           => n712);
   U763 : AOI22_X1 port map( A1 => bht_14_14_port, A2 => n118, B1 => 
                           bht_15_14_port, B2 => n119, ZN => n721);
   U764 : AOI22_X1 port map( A1 => bht_12_14_port, A2 => n120, B1 => 
                           bht_13_14_port, B2 => n121, ZN => n720);
   U765 : AOI22_X1 port map( A1 => bht_10_14_port, A2 => n122, B1 => 
                           bht_11_14_port, B2 => n123, ZN => n719);
   U766 : AOI22_X1 port map( A1 => bht_8_14_port, A2 => n124, B1 => 
                           bht_9_14_port, B2 => n125_port, ZN => n718);
   U767 : NAND4_X1 port map( A1 => n722, A2 => n723, A3 => n724, A4 => n725, ZN
                           => n711);
   U768 : AOI22_X1 port map( A1 => bht_22_14_port, A2 => n154, B1 => 
                           bht_23_14_port, B2 => n155, ZN => n725);
   U769 : AOI22_X1 port map( A1 => bht_20_14_port, A2 => n156, B1 => 
                           bht_21_14_port, B2 => n157, ZN => n724);
   U770 : AOI22_X1 port map( A1 => bht_18_14_port, A2 => n158, B1 => 
                           bht_19_14_port, B2 => n159, ZN => n723);
   U771 : AOI22_X1 port map( A1 => bht_16_14_port, A2 => n160, B1 => 
                           bht_17_14_port, B2 => n161, ZN => n722);
   U772 : NAND4_X1 port map( A1 => n726, A2 => n727, A3 => n728, A4 => n729, ZN
                           => n710);
   U773 : AOI22_X1 port map( A1 => bht_30_14_port, A2 => n142_port, B1 => 
                           bht_31_14_port, B2 => n143_port, ZN => n729);
   U774 : AOI22_X1 port map( A1 => bht_28_14_port, A2 => n144_port, B1 => 
                           bht_29_14_port, B2 => n145_port, ZN => n728);
   U775 : AOI22_X1 port map( A1 => bht_26_14_port, A2 => n146_port, B1 => 
                           bht_27_14_port, B2 => n147_port, ZN => n727);
   U776 : AOI22_X1 port map( A1 => bht_24_14_port, A2 => n148_port, B1 => 
                           bht_25_14_port, B2 => n149_port, ZN => n726);
   U777 : MUX2_X1 port map( A => reg_a(6), B => addr(13), S => sig_bal, Z => 
                           n280);
   U778 : NOR4_X1 port map( A1 => n730, A2 => n731, A3 => n732, A4 => n733, ZN 
                           => n100);
   U779 : NAND4_X1 port map( A1 => n734, A2 => n735, A3 => n736, A4 => n737, ZN
                           => n733);
   U780 : AOI22_X1 port map( A1 => bht_6_8_port, A2 => n130_port, B1 => 
                           bht_7_8_port, B2 => n131_port, ZN => n737);
   U781 : AOI22_X1 port map( A1 => bht_4_8_port, A2 => n132_port, B1 => 
                           bht_5_8_port, B2 => n133_port, ZN => n736);
   U782 : AOI22_X1 port map( A1 => bht_2_8_port, A2 => n134_port, B1 => 
                           bht_3_8_port, B2 => n135_port, ZN => n735);
   U783 : AOI22_X1 port map( A1 => bht_0_8_port, A2 => n136_port, B1 => 
                           bht_1_8_port, B2 => n137_port, ZN => n734);
   U784 : NAND4_X1 port map( A1 => n738, A2 => n739, A3 => n740, A4 => n741, ZN
                           => n732);
   U785 : AOI22_X1 port map( A1 => bht_14_8_port, A2 => n118, B1 => 
                           bht_15_8_port, B2 => n119, ZN => n741);
   U786 : AOI22_X1 port map( A1 => bht_12_8_port, A2 => n120, B1 => 
                           bht_13_8_port, B2 => n121, ZN => n740);
   U787 : AOI22_X1 port map( A1 => bht_10_8_port, A2 => n122, B1 => 
                           bht_11_8_port, B2 => n123, ZN => n739);
   U788 : AOI22_X1 port map( A1 => bht_8_8_port, A2 => n124, B1 => bht_9_8_port
                           , B2 => n125_port, ZN => n738);
   U789 : NAND4_X1 port map( A1 => n742, A2 => n743, A3 => n744, A4 => n745, ZN
                           => n731);
   U790 : AOI22_X1 port map( A1 => bht_22_8_port, A2 => n154, B1 => 
                           bht_23_8_port, B2 => n155, ZN => n745);
   U791 : AOI22_X1 port map( A1 => bht_20_8_port, A2 => n156, B1 => 
                           bht_21_8_port, B2 => n157, ZN => n744);
   U792 : AOI22_X1 port map( A1 => bht_18_8_port, A2 => n158, B1 => 
                           bht_19_8_port, B2 => n159, ZN => n743);
   U793 : AOI22_X1 port map( A1 => bht_16_8_port, A2 => n160, B1 => 
                           bht_17_8_port, B2 => n161, ZN => n742);
   U794 : NAND4_X1 port map( A1 => n746, A2 => n747, A3 => n748, A4 => n749, ZN
                           => n730);
   U795 : AOI22_X1 port map( A1 => bht_30_8_port, A2 => n142_port, B1 => 
                           bht_31_8_port, B2 => n143_port, ZN => n749);
   U796 : AOI22_X1 port map( A1 => bht_28_8_port, A2 => n144_port, B1 => 
                           bht_29_8_port, B2 => n145_port, ZN => n748);
   U797 : AOI22_X1 port map( A1 => bht_26_8_port, A2 => n146_port, B1 => 
                           bht_27_8_port, B2 => n147_port, ZN => n747);
   U798 : AOI22_X1 port map( A1 => bht_24_8_port, A2 => n148_port, B1 => 
                           bht_25_8_port, B2 => n149_port, ZN => n746);
   U799 : NOR4_X1 port map( A1 => n750, A2 => n751, A3 => n752, A4 => n753, ZN 
                           => n162);
   U800 : NAND4_X1 port map( A1 => n754, A2 => n755, A3 => n756, A4 => n757, ZN
                           => n753);
   U801 : AOI22_X1 port map( A1 => bht_14_0_port, A2 => n118, B1 => 
                           bht_15_0_port, B2 => n119, ZN => n757);
   U802 : AOI22_X1 port map( A1 => bht_12_0_port, A2 => n120, B1 => 
                           bht_13_0_port, B2 => n121, ZN => n756);
   U803 : AOI22_X1 port map( A1 => bht_10_0_port, A2 => n122, B1 => 
                           bht_11_0_port, B2 => n123, ZN => n755);
   U804 : AOI22_X1 port map( A1 => bht_8_0_port, A2 => n124, B1 => bht_9_0_port
                           , B2 => n125_port, ZN => n754);
   U805 : NOR3_X1 port map( A1 => n764, A2 => addr(6), A3 => n765, ZN => n758);
   U806 : NOR3_X1 port map( A1 => addr(2), A2 => addr(6), A3 => n764, ZN => 
                           n760);
   U807 : NAND4_X1 port map( A1 => n766, A2 => n767, A3 => n768, A4 => n769, ZN
                           => n752);
   U808 : AOI22_X1 port map( A1 => bht_6_0_port, A2 => n130_port, B1 => 
                           bht_7_0_port, B2 => n131_port, ZN => n769);
   U809 : AOI22_X1 port map( A1 => bht_4_0_port, A2 => n132_port, B1 => 
                           bht_5_0_port, B2 => n133_port, ZN => n768);
   U810 : AOI22_X1 port map( A1 => bht_2_0_port, A2 => n134_port, B1 => 
                           bht_3_0_port, B2 => n135_port, ZN => n767);
   U811 : AOI22_X1 port map( A1 => bht_0_0_port, A2 => n136_port, B1 => 
                           bht_1_0_port, B2 => n137_port, ZN => n766);
   U812 : NOR3_X1 port map( A1 => addr(5), A2 => addr(6), A3 => n765, ZN => 
                           n770);
   U813 : NOR3_X1 port map( A1 => addr(5), A2 => addr(6), A3 => addr(2), ZN => 
                           n771);
   U814 : NAND4_X1 port map( A1 => n772, A2 => n773, A3 => n774, A4 => n775, ZN
                           => n751);
   U815 : AOI22_X1 port map( A1 => bht_30_0_port, A2 => n142_port, B1 => 
                           bht_31_0_port, B2 => n143_port, ZN => n775);
   U816 : AOI22_X1 port map( A1 => bht_28_0_port, A2 => n144_port, B1 => 
                           bht_29_0_port, B2 => n145_port, ZN => n774);
   U817 : AOI22_X1 port map( A1 => bht_26_0_port, A2 => n146_port, B1 => 
                           bht_27_0_port, B2 => n147_port, ZN => n773);
   U818 : AOI22_X1 port map( A1 => bht_24_0_port, A2 => n148_port, B1 => 
                           bht_25_0_port, B2 => n149_port, ZN => n772);
   U819 : NOR3_X1 port map( A1 => n765, A2 => n764, A3 => n778, ZN => n776);
   U820 : NOR3_X1 port map( A1 => n764, A2 => addr(2), A3 => n778, ZN => n777);
   U821 : INV_X1 port map( A => addr(5), ZN => n764);
   U822 : NAND4_X1 port map( A1 => n779, A2 => n780, A3 => n781, A4 => n782, ZN
                           => n750);
   U823 : AOI22_X1 port map( A1 => bht_22_0_port, A2 => n154, B1 => 
                           bht_23_0_port, B2 => n155, ZN => n782);
   U824 : AND2_X1 port map( A1 => addr(4), A2 => addr(3), ZN => n759);
   U825 : AOI22_X1 port map( A1 => bht_20_0_port, A2 => n156, B1 => 
                           bht_21_0_port, B2 => n157, ZN => n781);
   U826 : AND2_X1 port map( A1 => addr(4), A2 => n785, ZN => n761);
   U827 : AOI22_X1 port map( A1 => bht_18_0_port, A2 => n158, B1 => 
                           bht_19_0_port, B2 => n159, ZN => n780);
   U828 : NOR2_X1 port map( A1 => n785, A2 => addr(4), ZN => n762);
   U829 : INV_X1 port map( A => addr(3), ZN => n785);
   U830 : AOI22_X1 port map( A1 => bht_16_0_port, A2 => n160, B1 => 
                           bht_17_0_port, B2 => n161, ZN => n779);
   U831 : NOR3_X1 port map( A1 => n765, A2 => addr(5), A3 => n778, ZN => n783);
   U832 : INV_X1 port map( A => addr(2), ZN => n765);
   U833 : NOR2_X1 port map( A1 => addr(3), A2 => addr(4), ZN => n763);
   U834 : NOR3_X1 port map( A1 => addr(2), A2 => addr(5), A3 => n778, ZN => 
                           n784);
   U835 : INV_X1 port map( A => addr(6), ZN => n778);

end SYN_branch_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity StallGenerator_CWRD_SIZE20 is

   port( rst, clk, sig_ral, sig_bpw, sig_jral, sig_mul, sig_div, sig_sqrt : in 
         std_logic;  stall_flag : out std_logic_vector (4 downto 0));

end StallGenerator_CWRD_SIZE20;

architecture SYN_stall_generator_arch of StallGenerator_CWRD_SIZE20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X4
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component StallGenerator_CWRD_SIZE20_DW01_inc_5
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component StallGenerator_CWRD_SIZE20_DW01_inc_4
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component StallGenerator_CWRD_SIZE20_DW01_inc_3
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component StallGenerator_CWRD_SIZE20_DW01_inc_2
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component StallGenerator_CWRD_SIZE20_DW01_inc_1
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component StallGenerator_CWRD_SIZE20_DW01_inc_0
      port( A : in std_logic_vector (31 downto 0);  SUM : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal stall_flag_3_port, stall_flag_2_port, stall_flag_1_port, 
      stall_flag_0_port, n_state_ral_31_port, n_state_ral_30_port, 
      n_state_ral_29_port, n_state_ral_28_port, n_state_ral_27_port, 
      n_state_ral_26_port, n_state_ral_25_port, n_state_ral_24_port, 
      n_state_ral_23_port, n_state_ral_22_port, n_state_ral_21_port, 
      n_state_ral_20_port, n_state_ral_19_port, n_state_ral_18_port, 
      n_state_ral_17_port, n_state_ral_16_port, n_state_ral_15_port, 
      n_state_ral_14_port, n_state_ral_13_port, n_state_ral_12_port, 
      n_state_ral_11_port, n_state_ral_10_port, n_state_ral_9_port, 
      n_state_ral_8_port, n_state_ral_7_port, n_state_ral_6_port, 
      n_state_ral_5_port, n_state_ral_4_port, n_state_ral_3_port, 
      n_state_ral_2_port, n_state_ral_1_port, n_state_ral_0_port, 
      c_state_ral_31_port, c_state_ral_30_port, c_state_ral_29_port, 
      c_state_ral_28_port, c_state_ral_27_port, c_state_ral_26_port, 
      c_state_ral_25_port, c_state_ral_24_port, c_state_ral_23_port, 
      c_state_ral_22_port, c_state_ral_21_port, c_state_ral_20_port, 
      c_state_ral_19_port, c_state_ral_18_port, c_state_ral_17_port, 
      c_state_ral_16_port, c_state_ral_15_port, c_state_ral_14_port, 
      c_state_ral_13_port, c_state_ral_12_port, c_state_ral_11_port, 
      c_state_ral_10_port, c_state_ral_9_port, c_state_ral_8_port, 
      c_state_ral_7_port, c_state_ral_6_port, c_state_ral_5_port, 
      c_state_ral_4_port, c_state_ral_3_port, c_state_ral_2_port, 
      c_state_ral_1_port, c_state_ral_0_port, N46, N47, N48, N49, N50, N51, N52
      , N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64, N65, N66, 
      N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77, 
      n_state_bpw_31_port, n_state_bpw_30_port, n_state_bpw_29_port, 
      n_state_bpw_28_port, n_state_bpw_27_port, n_state_bpw_26_port, 
      n_state_bpw_25_port, n_state_bpw_24_port, n_state_bpw_23_port, 
      n_state_bpw_22_port, n_state_bpw_21_port, n_state_bpw_20_port, 
      n_state_bpw_19_port, n_state_bpw_18_port, n_state_bpw_17_port, 
      n_state_bpw_16_port, n_state_bpw_15_port, n_state_bpw_14_port, 
      n_state_bpw_13_port, n_state_bpw_12_port, n_state_bpw_11_port, 
      n_state_bpw_10_port, n_state_bpw_9_port, n_state_bpw_8_port, 
      n_state_bpw_7_port, n_state_bpw_6_port, n_state_bpw_5_port, 
      n_state_bpw_4_port, n_state_bpw_3_port, n_state_bpw_2_port, 
      n_state_bpw_1_port, n_state_bpw_0_port, c_state_bpw_31_port, 
      c_state_bpw_30_port, c_state_bpw_29_port, c_state_bpw_28_port, 
      c_state_bpw_27_port, c_state_bpw_26_port, c_state_bpw_25_port, 
      c_state_bpw_24_port, c_state_bpw_23_port, c_state_bpw_22_port, 
      c_state_bpw_21_port, c_state_bpw_20_port, c_state_bpw_19_port, 
      c_state_bpw_18_port, c_state_bpw_17_port, c_state_bpw_16_port, 
      c_state_bpw_15_port, c_state_bpw_14_port, c_state_bpw_13_port, 
      c_state_bpw_12_port, c_state_bpw_11_port, c_state_bpw_10_port, 
      c_state_bpw_9_port, c_state_bpw_8_port, c_state_bpw_7_port, 
      c_state_bpw_6_port, c_state_bpw_5_port, c_state_bpw_4_port, 
      c_state_bpw_3_port, c_state_bpw_2_port, c_state_bpw_1_port, 
      c_state_bpw_0_port, N119, N120, N121, N122, N123, N124, N125, N126, N127,
      N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139, 
      N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150, 
      c_state_mul_31_port, c_state_mul_30_port, c_state_mul_29_port, 
      c_state_mul_28_port, c_state_mul_27_port, c_state_mul_26_port, 
      c_state_mul_25_port, c_state_mul_24_port, c_state_mul_23_port, 
      c_state_mul_22_port, c_state_mul_21_port, c_state_mul_20_port, 
      c_state_mul_19_port, c_state_mul_18_port, c_state_mul_17_port, 
      c_state_mul_16_port, c_state_mul_15_port, c_state_mul_14_port, 
      c_state_mul_13_port, c_state_mul_12_port, c_state_mul_11_port, 
      c_state_mul_10_port, c_state_mul_9_port, c_state_mul_8_port, 
      c_state_mul_7_port, c_state_mul_6_port, c_state_mul_5_port, 
      c_state_mul_4_port, c_state_mul_3_port, c_state_mul_2_port, 
      c_state_mul_1_port, c_state_mul_0_port, n_state_mul_31_port, 
      n_state_mul_30_port, n_state_mul_29_port, n_state_mul_28_port, 
      n_state_mul_27_port, n_state_mul_26_port, n_state_mul_25_port, 
      n_state_mul_24_port, n_state_mul_23_port, n_state_mul_22_port, 
      n_state_mul_21_port, n_state_mul_20_port, n_state_mul_19_port, 
      n_state_mul_18_port, n_state_mul_17_port, n_state_mul_16_port, 
      n_state_mul_15_port, n_state_mul_14_port, n_state_mul_13_port, 
      n_state_mul_12_port, n_state_mul_11_port, n_state_mul_10_port, 
      n_state_mul_9_port, n_state_mul_8_port, n_state_mul_7_port, 
      n_state_mul_6_port, n_state_mul_5_port, n_state_mul_4_port, 
      n_state_mul_3_port, n_state_mul_2_port, n_state_mul_1_port, 
      n_state_mul_0_port, N193, N194, N195, N196, N197, N198, N199, N200, N201,
      N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212, N213, 
      N214, N215, N216, N217, N218, N219, N220, N221, N222, N223, N224, 
      c_state_div_31_port, c_state_div_30_port, c_state_div_29_port, 
      c_state_div_28_port, c_state_div_27_port, c_state_div_26_port, 
      c_state_div_25_port, c_state_div_24_port, c_state_div_23_port, 
      c_state_div_22_port, c_state_div_21_port, c_state_div_20_port, 
      c_state_div_19_port, c_state_div_18_port, c_state_div_17_port, 
      c_state_div_16_port, c_state_div_15_port, c_state_div_14_port, 
      c_state_div_13_port, c_state_div_12_port, c_state_div_11_port, 
      c_state_div_10_port, c_state_div_9_port, c_state_div_8_port, 
      c_state_div_7_port, c_state_div_6_port, c_state_div_5_port, 
      c_state_div_4_port, c_state_div_3_port, c_state_div_2_port, 
      c_state_div_1_port, c_state_div_0_port, n_state_div_31_port, 
      n_state_div_30_port, n_state_div_29_port, n_state_div_28_port, 
      n_state_div_27_port, n_state_div_26_port, n_state_div_25_port, 
      n_state_div_24_port, n_state_div_23_port, n_state_div_22_port, 
      n_state_div_21_port, n_state_div_20_port, n_state_div_19_port, 
      n_state_div_18_port, n_state_div_17_port, n_state_div_16_port, 
      n_state_div_15_port, n_state_div_14_port, n_state_div_13_port, 
      n_state_div_12_port, n_state_div_11_port, n_state_div_10_port, 
      n_state_div_9_port, n_state_div_8_port, n_state_div_7_port, 
      n_state_div_6_port, n_state_div_5_port, n_state_div_4_port, 
      n_state_div_3_port, n_state_div_2_port, n_state_div_1_port, 
      n_state_div_0_port, N278, N279, N280, N281, N282, N283, N284, N285, N286,
      N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, 
      N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N309, 
      c_state_sqrt_31_port, c_state_sqrt_30_port, c_state_sqrt_29_port, 
      c_state_sqrt_28_port, c_state_sqrt_27_port, c_state_sqrt_26_port, 
      c_state_sqrt_25_port, c_state_sqrt_24_port, c_state_sqrt_23_port, 
      c_state_sqrt_22_port, c_state_sqrt_21_port, c_state_sqrt_20_port, 
      c_state_sqrt_19_port, c_state_sqrt_18_port, c_state_sqrt_17_port, 
      c_state_sqrt_16_port, c_state_sqrt_15_port, c_state_sqrt_14_port, 
      c_state_sqrt_13_port, c_state_sqrt_12_port, c_state_sqrt_11_port, 
      c_state_sqrt_10_port, c_state_sqrt_9_port, c_state_sqrt_8_port, 
      c_state_sqrt_7_port, c_state_sqrt_6_port, c_state_sqrt_5_port, 
      c_state_sqrt_4_port, c_state_sqrt_3_port, c_state_sqrt_2_port, 
      c_state_sqrt_1_port, c_state_sqrt_0_port, n_state_sqrt_31_port, 
      n_state_sqrt_30_port, n_state_sqrt_29_port, n_state_sqrt_28_port, 
      n_state_sqrt_27_port, n_state_sqrt_26_port, n_state_sqrt_25_port, 
      n_state_sqrt_24_port, n_state_sqrt_23_port, n_state_sqrt_22_port, 
      n_state_sqrt_21_port, n_state_sqrt_20_port, n_state_sqrt_19_port, 
      n_state_sqrt_18_port, n_state_sqrt_17_port, n_state_sqrt_16_port, 
      n_state_sqrt_15_port, n_state_sqrt_14_port, n_state_sqrt_13_port, 
      n_state_sqrt_12_port, n_state_sqrt_11_port, n_state_sqrt_10_port, 
      n_state_sqrt_9_port, n_state_sqrt_8_port, n_state_sqrt_7_port, 
      n_state_sqrt_6_port, n_state_sqrt_5_port, n_state_sqrt_4_port, 
      n_state_sqrt_3_port, n_state_sqrt_2_port, n_state_sqrt_1_port, 
      n_state_sqrt_0_port, N363, N364, N365, N366, N367, N368, N369, N370, N371
      , N372, N373, N374, N375, N376, N377, N378, N379, N380, N381, N382, N383,
      N384, N385, N386, N387, N388, N389, N390, N391, N392, N393, N394, 
      c_state_stu_31_port, c_state_stu_30_port, c_state_stu_29_port, 
      c_state_stu_28_port, c_state_stu_27_port, c_state_stu_26_port, 
      c_state_stu_25_port, c_state_stu_24_port, c_state_stu_23_port, 
      c_state_stu_22_port, c_state_stu_21_port, c_state_stu_20_port, 
      c_state_stu_19_port, c_state_stu_18_port, c_state_stu_17_port, 
      c_state_stu_16_port, c_state_stu_15_port, c_state_stu_14_port, 
      c_state_stu_13_port, c_state_stu_12_port, c_state_stu_11_port, 
      c_state_stu_10_port, c_state_stu_9_port, c_state_stu_8_port, 
      c_state_stu_7_port, c_state_stu_6_port, c_state_stu_5_port, 
      c_state_stu_4_port, c_state_stu_3_port, c_state_stu_2_port, 
      c_state_stu_1_port, c_state_stu_0_port, n_state_stu_31_port, 
      n_state_stu_30_port, n_state_stu_29_port, n_state_stu_28_port, 
      n_state_stu_27_port, n_state_stu_26_port, n_state_stu_25_port, 
      n_state_stu_24_port, n_state_stu_23_port, n_state_stu_22_port, 
      n_state_stu_21_port, n_state_stu_20_port, n_state_stu_19_port, 
      n_state_stu_18_port, n_state_stu_17_port, n_state_stu_16_port, 
      n_state_stu_15_port, n_state_stu_14_port, n_state_stu_13_port, 
      n_state_stu_12_port, n_state_stu_11_port, n_state_stu_10_port, 
      n_state_stu_9_port, n_state_stu_8_port, n_state_stu_7_port, 
      n_state_stu_6_port, n_state_stu_5_port, n_state_stu_4_port, 
      n_state_stu_3_port, n_state_stu_2_port, n_state_stu_1_port, 
      n_state_stu_0_port, N444, N445, N446, N447, N448, N449, N450, N451, N452,
      N453, N454, N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, 
      N465, N466, N467, N468, N469, N470, N471, N472, N473, N474, N475, n192, 
      n194_port, n195_port, n197_port, n214_port, n222_port, n230, n231, n232, 
      n247, n261, n262, n263, n264, n266, n267, n271, n276, n294_port, 
      n307_port, n308_port, n309_port, n310, n311, n312, n316, n317, n318, n323
      , n328, n342, n343, n344, n345, n347, n348, n352, n357, n1, n2, n3, n4, 
      n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20
      , n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, 
      n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46_port, n47_port
      , n48_port, n49_port, n50_port, n51_port, n52_port, n53_port, n54_port, 
      n55_port, n56_port, n57_port, n58_port, n59_port, n60_port, n61_port, 
      n62_port, n63_port, n64_port, n65_port, n66_port, n67_port, n68_port, 
      n69_port, n70_port, n71_port, n72_port, n73_port, n74_port, n75_port, 
      n76_port, n77_port, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88
      , n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102
      , n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
      n115, n116, n117, n118, n119_port, n120_port, n121_port, n122_port, 
      n123_port, n124_port, n125_port, n126_port, n127_port, n128_port, 
      n129_port, n130_port, n131_port, n132_port, n133_port, n134_port, 
      n135_port, n136_port, n137_port, n138_port, n139_port, n140_port, 
      n141_port, n142_port, n143_port, n144_port, n145_port, n146_port, 
      n147_port, n148_port, n149_port, n150_port, n151, n152, n153, n154, n155,
      n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, 
      n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n193_port, n196_port, n198_port, n199_port, n200_port, n201_port, 
      n202_port, n203_port, n204_port, n205_port, n206_port, n207_port, 
      n208_port, n209_port, n210_port, n211_port, n212_port, n213_port, 
      n215_port, n216_port, n217_port, n218_port, n219_port, n220_port, 
      n221_port, n223_port, n224_port, n225, n226, n227, n228, n229, n233, n234
      , n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
      n248, n249, net107995, net107996, net107997, net107998, net107999, 
      net108000, net108001, net108002, net108003, net108004, net108005, 
      net108006, net108007, net108008, net108009, net108010, net108011, 
      net108012, net108013, net108014, net108015, net108016, net108017, 
      net108018, net108019, net108020, net108021, net108022, net108023, 
      net108024, net108025, net108026, net108027, net108028, net108029, 
      net108030, net108031, net108032, net108033, net108034, net108035, 
      net108036, net108037, net108038, net108039, net108040, net108041, 
      net108042, net108043, net108044, net108045, net108046, net108047, 
      net108048, net108049, net108050, net108051, net108052, net108053, 
      net108054, net108055, net108056, net108057, net108058, net108059, 
      net108060, net108061, net108062, net108063 : std_logic;

begin
   stall_flag <= ( stall_flag_3_port, stall_flag_3_port, stall_flag_2_port, 
      stall_flag_1_port, stall_flag_0_port );
   
   c_state_ral_reg_0_inst : DFFR_X1 port map( D => n_state_ral_0_port, CK => 
                           clk, RN => rst, Q => c_state_ral_0_port, QN => 
                           n195_port);
   c_state_ral_reg_10_inst : DFFR_X1 port map( D => n_state_ral_10_port, CK => 
                           clk, RN => rst, Q => c_state_ral_10_port, QN => 
                           net108063);
   c_state_ral_reg_1_inst : DFFR_X1 port map( D => n_state_ral_1_port, CK => 
                           clk, RN => rst, Q => c_state_ral_1_port, QN => n231)
                           ;
   c_state_ral_reg_2_inst : DFFR_X1 port map( D => n_state_ral_2_port, CK => 
                           clk, RN => rst, Q => c_state_ral_2_port, QN => 
                           net108062);
   c_state_ral_reg_3_inst : DFFR_X1 port map( D => n_state_ral_3_port, CK => 
                           clk, RN => rst, Q => c_state_ral_3_port, QN => 
                           net108061);
   c_state_ral_reg_4_inst : DFFR_X1 port map( D => n_state_ral_4_port, CK => 
                           clk, RN => rst, Q => c_state_ral_4_port, QN => 
                           n209_port);
   c_state_ral_reg_5_inst : DFFR_X1 port map( D => n_state_ral_5_port, CK => 
                           clk, RN => rst, Q => c_state_ral_5_port, QN => 
                           n208_port);
   c_state_ral_reg_6_inst : DFFR_X1 port map( D => n_state_ral_6_port, CK => 
                           clk, RN => rst, Q => c_state_ral_6_port, QN => 
                           n207_port);
   c_state_ral_reg_7_inst : DFFR_X1 port map( D => n_state_ral_7_port, CK => 
                           clk, RN => rst, Q => c_state_ral_7_port, QN => 
                           n206_port);
   c_state_ral_reg_8_inst : DFFR_X1 port map( D => n_state_ral_8_port, CK => 
                           clk, RN => rst, Q => c_state_ral_8_port, QN => 
                           net108060);
   c_state_ral_reg_9_inst : DFFR_X1 port map( D => n_state_ral_9_port, CK => 
                           clk, RN => rst, Q => c_state_ral_9_port, QN => 
                           net108059);
   c_state_ral_reg_11_inst : DFFR_X1 port map( D => n_state_ral_11_port, CK => 
                           clk, RN => rst, Q => c_state_ral_11_port, QN => 
                           net108058);
   c_state_ral_reg_12_inst : DFFR_X1 port map( D => n_state_ral_12_port, CK => 
                           clk, RN => rst, Q => c_state_ral_12_port, QN => 
                           n205_port);
   c_state_ral_reg_13_inst : DFFR_X1 port map( D => n_state_ral_13_port, CK => 
                           clk, RN => rst, Q => c_state_ral_13_port, QN => 
                           n204_port);
   c_state_ral_reg_14_inst : DFFR_X1 port map( D => n_state_ral_14_port, CK => 
                           clk, RN => rst, Q => c_state_ral_14_port, QN => 
                           n203_port);
   c_state_ral_reg_15_inst : DFFR_X1 port map( D => n_state_ral_15_port, CK => 
                           clk, RN => rst, Q => c_state_ral_15_port, QN => 
                           n202_port);
   c_state_ral_reg_16_inst : DFFR_X1 port map( D => n_state_ral_16_port, CK => 
                           clk, RN => rst, Q => c_state_ral_16_port, QN => 
                           net108057);
   c_state_ral_reg_17_inst : DFFR_X1 port map( D => n_state_ral_17_port, CK => 
                           clk, RN => rst, Q => c_state_ral_17_port, QN => 
                           net108056);
   c_state_ral_reg_18_inst : DFFR_X1 port map( D => n_state_ral_18_port, CK => 
                           clk, RN => rst, Q => c_state_ral_18_port, QN => 
                           net108055);
   c_state_ral_reg_19_inst : DFFR_X1 port map( D => n_state_ral_19_port, CK => 
                           clk, RN => rst, Q => c_state_ral_19_port, QN => 
                           n201_port);
   c_state_ral_reg_20_inst : DFFR_X1 port map( D => n_state_ral_20_port, CK => 
                           clk, RN => rst, Q => c_state_ral_20_port, QN => 
                           n200_port);
   c_state_ral_reg_21_inst : DFFR_X1 port map( D => n_state_ral_21_port, CK => 
                           clk, RN => rst, Q => c_state_ral_21_port, QN => 
                           n199_port);
   c_state_ral_reg_22_inst : DFFR_X1 port map( D => n_state_ral_22_port, CK => 
                           clk, RN => rst, Q => c_state_ral_22_port, QN => 
                           n198_port);
   c_state_ral_reg_23_inst : DFFR_X1 port map( D => n_state_ral_23_port, CK => 
                           clk, RN => rst, Q => c_state_ral_23_port, QN => 
                           n196_port);
   c_state_ral_reg_24_inst : DFFR_X1 port map( D => n_state_ral_24_port, CK => 
                           clk, RN => rst, Q => c_state_ral_24_port, QN => 
                           n193_port);
   c_state_ral_reg_25_inst : DFFR_X1 port map( D => n_state_ral_25_port, CK => 
                           clk, RN => rst, Q => c_state_ral_25_port, QN => n191
                           );
   c_state_ral_reg_26_inst : DFFR_X1 port map( D => n_state_ral_26_port, CK => 
                           clk, RN => rst, Q => c_state_ral_26_port, QN => n190
                           );
   c_state_ral_reg_27_inst : DFFR_X1 port map( D => n_state_ral_27_port, CK => 
                           clk, RN => rst, Q => c_state_ral_27_port, QN => n189
                           );
   c_state_ral_reg_28_inst : DFFR_X1 port map( D => n_state_ral_28_port, CK => 
                           clk, RN => rst, Q => c_state_ral_28_port, QN => n188
                           );
   c_state_ral_reg_29_inst : DFFR_X1 port map( D => n_state_ral_29_port, CK => 
                           clk, RN => rst, Q => c_state_ral_29_port, QN => n187
                           );
   c_state_ral_reg_30_inst : DFFR_X1 port map( D => n_state_ral_30_port, CK => 
                           clk, RN => rst, Q => c_state_ral_30_port, QN => n186
                           );
   c_state_ral_reg_31_inst : DFFR_X1 port map( D => n_state_ral_31_port, CK => 
                           clk, RN => rst, Q => c_state_ral_31_port, QN => n185
                           );
   c_state_bpw_reg_0_inst : DFFR_X1 port map( D => n_state_bpw_0_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_0_port, QN => 
                           n197_port);
   c_state_bpw_reg_10_inst : DFFR_X1 port map( D => n_state_bpw_10_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_10_port, QN => 
                           net108054);
   c_state_bpw_reg_1_inst : DFFR_X1 port map( D => n_state_bpw_1_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_1_port, QN => n232)
                           ;
   c_state_bpw_reg_2_inst : DFFR_X1 port map( D => n_state_bpw_2_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_2_port, QN => 
                           net108053);
   c_state_bpw_reg_3_inst : DFFR_X1 port map( D => n_state_bpw_3_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_3_port, QN => 
                           net108052);
   c_state_bpw_reg_4_inst : DFFR_X1 port map( D => n_state_bpw_4_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_4_port, QN => n184)
                           ;
   c_state_bpw_reg_5_inst : DFFR_X1 port map( D => n_state_bpw_5_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_5_port, QN => n183)
                           ;
   c_state_bpw_reg_6_inst : DFFR_X1 port map( D => n_state_bpw_6_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_6_port, QN => n182)
                           ;
   c_state_bpw_reg_7_inst : DFFR_X1 port map( D => n_state_bpw_7_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_7_port, QN => n181)
                           ;
   c_state_bpw_reg_8_inst : DFFR_X1 port map( D => n_state_bpw_8_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_8_port, QN => 
                           net108051);
   c_state_bpw_reg_9_inst : DFFR_X1 port map( D => n_state_bpw_9_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_9_port, QN => 
                           net108050);
   c_state_bpw_reg_11_inst : DFFR_X1 port map( D => n_state_bpw_11_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_11_port, QN => 
                           net108049);
   c_state_bpw_reg_12_inst : DFFR_X1 port map( D => n_state_bpw_12_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_12_port, QN => n180
                           );
   c_state_bpw_reg_13_inst : DFFR_X1 port map( D => n_state_bpw_13_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_13_port, QN => n179
                           );
   c_state_bpw_reg_14_inst : DFFR_X1 port map( D => n_state_bpw_14_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_14_port, QN => n178
                           );
   c_state_bpw_reg_15_inst : DFFR_X1 port map( D => n_state_bpw_15_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_15_port, QN => n177
                           );
   c_state_bpw_reg_16_inst : DFFR_X1 port map( D => n_state_bpw_16_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_16_port, QN => 
                           net108048);
   c_state_bpw_reg_17_inst : DFFR_X1 port map( D => n_state_bpw_17_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_17_port, QN => 
                           net108047);
   c_state_bpw_reg_18_inst : DFFR_X1 port map( D => n_state_bpw_18_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_18_port, QN => 
                           net108046);
   c_state_bpw_reg_19_inst : DFFR_X1 port map( D => n_state_bpw_19_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_19_port, QN => n176
                           );
   c_state_bpw_reg_20_inst : DFFR_X1 port map( D => n_state_bpw_20_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_20_port, QN => n175
                           );
   c_state_bpw_reg_21_inst : DFFR_X1 port map( D => n_state_bpw_21_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_21_port, QN => n174
                           );
   c_state_bpw_reg_22_inst : DFFR_X1 port map( D => n_state_bpw_22_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_22_port, QN => n173
                           );
   c_state_bpw_reg_23_inst : DFFR_X1 port map( D => n_state_bpw_23_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_23_port, QN => n172
                           );
   c_state_bpw_reg_24_inst : DFFR_X1 port map( D => n_state_bpw_24_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_24_port, QN => n171
                           );
   c_state_bpw_reg_25_inst : DFFR_X1 port map( D => n_state_bpw_25_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_25_port, QN => n170
                           );
   c_state_bpw_reg_26_inst : DFFR_X1 port map( D => n_state_bpw_26_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_26_port, QN => n169
                           );
   c_state_bpw_reg_27_inst : DFFR_X1 port map( D => n_state_bpw_27_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_27_port, QN => n168
                           );
   c_state_bpw_reg_28_inst : DFFR_X1 port map( D => n_state_bpw_28_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_28_port, QN => n167
                           );
   c_state_bpw_reg_29_inst : DFFR_X1 port map( D => n_state_bpw_29_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_29_port, QN => n166
                           );
   c_state_bpw_reg_30_inst : DFFR_X1 port map( D => n_state_bpw_30_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_30_port, QN => n165
                           );
   c_state_bpw_reg_31_inst : DFFR_X1 port map( D => n_state_bpw_31_port, CK => 
                           clk, RN => rst, Q => c_state_bpw_31_port, QN => n164
                           );
   c_state_mul_reg_0_inst : DFFR_X1 port map( D => n_state_mul_0_port, CK => 
                           clk, RN => rst, Q => c_state_mul_0_port, QN => 
                           n294_port);
   c_state_mul_reg_10_inst : DFFR_X1 port map( D => n_state_mul_10_port, CK => 
                           clk, RN => rst, Q => c_state_mul_10_port, QN => n323
                           );
   c_state_mul_reg_1_inst : DFFR_X1 port map( D => n_state_mul_1_port, CK => 
                           clk, RN => rst, Q => c_state_mul_1_port, QN => n163)
                           ;
   c_state_mul_reg_2_inst : DFFR_X1 port map( D => n_state_mul_2_port, CK => 
                           clk, RN => rst, Q => c_state_mul_2_port, QN => n310)
                           ;
   c_state_mul_reg_3_inst : DFFR_X1 port map( D => n_state_mul_3_port, CK => 
                           clk, RN => rst, Q => c_state_mul_3_port, QN => 
                           n222_port);
   c_state_mul_reg_4_inst : DFFR_X1 port map( D => n_state_mul_4_port, CK => 
                           clk, RN => rst, Q => c_state_mul_4_port, QN => 
                           net108045);
   c_state_mul_reg_5_inst : DFFR_X1 port map( D => n_state_mul_5_port, CK => 
                           clk, RN => rst, Q => c_state_mul_5_port, QN => 
                           net108044);
   c_state_mul_reg_6_inst : DFFR_X1 port map( D => n_state_mul_6_port, CK => 
                           clk, RN => rst, Q => c_state_mul_6_port, QN => 
                           net108043);
   c_state_mul_reg_7_inst : DFFR_X1 port map( D => n_state_mul_7_port, CK => 
                           clk, RN => rst, Q => c_state_mul_7_port, QN => n316)
                           ;
   c_state_mul_reg_8_inst : DFFR_X1 port map( D => n_state_mul_8_port, CK => 
                           clk, RN => rst, Q => c_state_mul_8_port, QN => n317)
                           ;
   c_state_mul_reg_9_inst : DFFR_X1 port map( D => n_state_mul_9_port, CK => 
                           clk, RN => rst, Q => c_state_mul_9_port, QN => n318)
                           ;
   c_state_mul_reg_11_inst : DFFR_X1 port map( D => n_state_mul_11_port, CK => 
                           clk, RN => rst, Q => c_state_mul_11_port, QN => 
                           net108042);
   c_state_mul_reg_12_inst : DFFR_X1 port map( D => n_state_mul_12_port, CK => 
                           clk, RN => rst, Q => c_state_mul_12_port, QN => 
                           net108041);
   c_state_mul_reg_13_inst : DFFR_X1 port map( D => n_state_mul_13_port, CK => 
                           clk, RN => rst, Q => c_state_mul_13_port, QN => 
                           net108040);
   c_state_mul_reg_14_inst : DFFR_X1 port map( D => n_state_mul_14_port, CK => 
                           clk, RN => rst, Q => c_state_mul_14_port, QN => n162
                           );
   c_state_mul_reg_15_inst : DFFR_X1 port map( D => n_state_mul_15_port, CK => 
                           clk, RN => rst, Q => c_state_mul_15_port, QN => n161
                           );
   c_state_mul_reg_16_inst : DFFR_X1 port map( D => n_state_mul_16_port, CK => 
                           clk, RN => rst, Q => c_state_mul_16_port, QN => n160
                           );
   c_state_mul_reg_17_inst : DFFR_X1 port map( D => n_state_mul_17_port, CK => 
                           clk, RN => rst, Q => c_state_mul_17_port, QN => 
                           net108039);
   c_state_mul_reg_18_inst : DFFR_X1 port map( D => n_state_mul_18_port, CK => 
                           clk, RN => rst, Q => c_state_mul_18_port, QN => 
                           net108038);
   c_state_mul_reg_19_inst : DFFR_X1 port map( D => n_state_mul_19_port, CK => 
                           clk, RN => rst, Q => c_state_mul_19_port, QN => 
                           net108037);
   c_state_mul_reg_20_inst : DFFR_X1 port map( D => n_state_mul_20_port, CK => 
                           clk, RN => rst, Q => c_state_mul_20_port, QN => n159
                           );
   c_state_mul_reg_21_inst : DFFR_X1 port map( D => n_state_mul_21_port, CK => 
                           clk, RN => rst, Q => c_state_mul_21_port, QN => n158
                           );
   c_state_mul_reg_22_inst : DFFR_X1 port map( D => n_state_mul_22_port, CK => 
                           clk, RN => rst, Q => c_state_mul_22_port, QN => n157
                           );
   c_state_mul_reg_23_inst : DFFR_X1 port map( D => n_state_mul_23_port, CK => 
                           clk, RN => rst, Q => c_state_mul_23_port, QN => n156
                           );
   c_state_mul_reg_24_inst : DFFR_X1 port map( D => n_state_mul_24_port, CK => 
                           clk, RN => rst, Q => c_state_mul_24_port, QN => 
                           net108036);
   c_state_mul_reg_25_inst : DFFR_X1 port map( D => n_state_mul_25_port, CK => 
                           clk, RN => rst, Q => c_state_mul_25_port, QN => 
                           net108035);
   c_state_mul_reg_26_inst : DFFR_X1 port map( D => n_state_mul_26_port, CK => 
                           clk, RN => rst, Q => c_state_mul_26_port, QN => 
                           net108034);
   c_state_mul_reg_27_inst : DFFR_X1 port map( D => n_state_mul_27_port, CK => 
                           clk, RN => rst, Q => c_state_mul_27_port, QN => 
                           n307_port);
   c_state_mul_reg_28_inst : DFFR_X1 port map( D => n_state_mul_28_port, CK => 
                           clk, RN => rst, Q => c_state_mul_28_port, QN => 
                           n308_port);
   c_state_mul_reg_29_inst : DFFR_X1 port map( D => n_state_mul_29_port, CK => 
                           clk, RN => rst, Q => c_state_mul_29_port, QN => 
                           n309_port);
   c_state_mul_reg_30_inst : DFFR_X1 port map( D => n_state_mul_30_port, CK => 
                           clk, RN => rst, Q => c_state_mul_30_port, QN => n311
                           );
   c_state_mul_reg_31_inst : DFFR_X1 port map( D => n_state_mul_31_port, CK => 
                           clk, RN => rst, Q => c_state_mul_31_port, QN => n312
                           );
   c_state_div_reg_0_inst : DFFR_X1 port map( D => n_state_div_0_port, CK => 
                           clk, RN => rst, Q => c_state_div_0_port, QN => n328)
                           ;
   c_state_div_reg_10_inst : DFFR_X1 port map( D => n_state_div_10_port, CK => 
                           clk, RN => rst, Q => c_state_div_10_port, QN => n357
                           );
   c_state_div_reg_1_inst : DFFR_X1 port map( D => n_state_div_1_port, CK => 
                           clk, RN => rst, Q => c_state_div_1_port, QN => n155)
                           ;
   c_state_div_reg_2_inst : DFFR_X1 port map( D => n_state_div_2_port, CK => 
                           clk, RN => rst, Q => c_state_div_2_port, QN => n344)
                           ;
   c_state_div_reg_3_inst : DFFR_X1 port map( D => n_state_div_3_port, CK => 
                           clk, RN => rst, Q => c_state_div_3_port, QN => n347)
                           ;
   c_state_div_reg_4_inst : DFFR_X1 port map( D => n_state_div_4_port, CK => 
                           clk, RN => rst, Q => c_state_div_4_port, QN => n348)
                           ;
   c_state_div_reg_5_inst : DFFR_X1 port map( D => n_state_div_5_port, CK => 
                           clk, RN => rst, Q => c_state_div_5_port, QN => n230)
                           ;
   c_state_div_reg_6_inst : DFFR_X1 port map( D => n_state_div_6_port, CK => 
                           clk, RN => rst, Q => c_state_div_6_port, QN => 
                           net108033);
   c_state_div_reg_7_inst : DFFR_X1 port map( D => n_state_div_7_port, CK => 
                           clk, RN => rst, Q => c_state_div_7_port, QN => 
                           net108032);
   c_state_div_reg_8_inst : DFFR_X1 port map( D => n_state_div_8_port, CK => 
                           clk, RN => rst, Q => c_state_div_8_port, QN => 
                           net108031);
   c_state_div_reg_9_inst : DFFR_X1 port map( D => n_state_div_9_port, CK => 
                           clk, RN => rst, Q => c_state_div_9_port, QN => n352)
                           ;
   c_state_div_reg_11_inst : DFFR_X1 port map( D => n_state_div_11_port, CK => 
                           clk, RN => rst, Q => c_state_div_11_port, QN => 
                           net108030);
   c_state_div_reg_12_inst : DFFR_X1 port map( D => n_state_div_12_port, CK => 
                           clk, RN => rst, Q => c_state_div_12_port, QN => 
                           net108029);
   c_state_div_reg_13_inst : DFFR_X1 port map( D => n_state_div_13_port, CK => 
                           clk, RN => rst, Q => c_state_div_13_port, QN => n249
                           );
   c_state_div_reg_14_inst : DFFR_X1 port map( D => n_state_div_14_port, CK => 
                           clk, RN => rst, Q => c_state_div_14_port, QN => n248
                           );
   c_state_div_reg_15_inst : DFFR_X1 port map( D => n_state_div_15_port, CK => 
                           clk, RN => rst, Q => c_state_div_15_port, QN => n246
                           );
   c_state_div_reg_16_inst : DFFR_X1 port map( D => n_state_div_16_port, CK => 
                           clk, RN => rst, Q => c_state_div_16_port, QN => 
                           net108028);
   c_state_div_reg_17_inst : DFFR_X1 port map( D => n_state_div_17_port, CK => 
                           clk, RN => rst, Q => c_state_div_17_port, QN => 
                           net108027);
   c_state_div_reg_18_inst : DFFR_X1 port map( D => n_state_div_18_port, CK => 
                           clk, RN => rst, Q => c_state_div_18_port, QN => 
                           net108026);
   c_state_div_reg_19_inst : DFFR_X1 port map( D => n_state_div_19_port, CK => 
                           clk, RN => rst, Q => c_state_div_19_port, QN => n245
                           );
   c_state_div_reg_20_inst : DFFR_X1 port map( D => n_state_div_20_port, CK => 
                           clk, RN => rst, Q => c_state_div_20_port, QN => n244
                           );
   c_state_div_reg_21_inst : DFFR_X1 port map( D => n_state_div_21_port, CK => 
                           clk, RN => rst, Q => c_state_div_21_port, QN => n243
                           );
   c_state_div_reg_22_inst : DFFR_X1 port map( D => n_state_div_22_port, CK => 
                           clk, RN => rst, Q => c_state_div_22_port, QN => 
                           net108025);
   c_state_div_reg_23_inst : DFFR_X1 port map( D => n_state_div_23_port, CK => 
                           clk, RN => rst, Q => c_state_div_23_port, QN => 
                           net108024);
   c_state_div_reg_24_inst : DFFR_X1 port map( D => n_state_div_24_port, CK => 
                           clk, RN => rst, Q => c_state_div_24_port, QN => 
                           net108023);
   c_state_div_reg_25_inst : DFFR_X1 port map( D => n_state_div_25_port, CK => 
                           clk, RN => rst, Q => c_state_div_25_port, QN => n242
                           );
   c_state_div_reg_26_inst : DFFR_X1 port map( D => n_state_div_26_port, CK => 
                           clk, RN => rst, Q => c_state_div_26_port, QN => n241
                           );
   c_state_div_reg_27_inst : DFFR_X1 port map( D => n_state_div_27_port, CK => 
                           clk, RN => rst, Q => c_state_div_27_port, QN => 
                           net108022);
   c_state_div_reg_28_inst : DFFR_X1 port map( D => n_state_div_28_port, CK => 
                           clk, RN => rst, Q => c_state_div_28_port, QN => n342
                           );
   c_state_div_reg_29_inst : DFFR_X1 port map( D => n_state_div_29_port, CK => 
                           clk, RN => rst, Q => c_state_div_29_port, QN => n343
                           );
   c_state_div_reg_30_inst : DFFR_X1 port map( D => n_state_div_30_port, CK => 
                           clk, RN => rst, Q => c_state_div_30_port, QN => n345
                           );
   c_state_div_reg_31_inst : DFFR_X1 port map( D => n_state_div_31_port, CK => 
                           clk, RN => rst, Q => c_state_div_31_port, QN => 
                           net108021);
   c_state_sqrt_reg_0_inst : DFFR_X1 port map( D => n_state_sqrt_0_port, CK => 
                           clk, RN => rst, Q => c_state_sqrt_0_port, QN => n247
                           );
   c_state_sqrt_reg_10_inst : DFFR_X1 port map( D => n_state_sqrt_10_port, CK 
                           => clk, RN => rst, Q => c_state_sqrt_10_port, QN => 
                           n276);
   c_state_sqrt_reg_1_inst : DFFR_X1 port map( D => n_state_sqrt_1_port, CK => 
                           clk, RN => rst, Q => c_state_sqrt_1_port, QN => n240
                           );
   c_state_sqrt_reg_2_inst : DFFR_X1 port map( D => n_state_sqrt_2_port, CK => 
                           clk, RN => rst, Q => c_state_sqrt_2_port, QN => n263
                           );
   c_state_sqrt_reg_3_inst : DFFR_X1 port map( D => n_state_sqrt_3_port, CK => 
                           clk, RN => rst, Q => c_state_sqrt_3_port, QN => n266
                           );
   c_state_sqrt_reg_4_inst : DFFR_X1 port map( D => n_state_sqrt_4_port, CK => 
                           clk, RN => rst, Q => c_state_sqrt_4_port, QN => 
                           net108020);
   c_state_sqrt_reg_5_inst : DFFR_X1 port map( D => n_state_sqrt_5_port, CK => 
                           clk, RN => rst, Q => c_state_sqrt_5_port, QN => n267
                           );
   c_state_sqrt_reg_6_inst : DFFR_X1 port map( D => n_state_sqrt_6_port, CK => 
                           clk, RN => rst, Q => c_state_sqrt_6_port, QN => 
                           net108019);
   c_state_sqrt_reg_7_inst : DFFR_X1 port map( D => n_state_sqrt_7_port, CK => 
                           clk, RN => rst, Q => c_state_sqrt_7_port, QN => 
                           net108018);
   c_state_sqrt_reg_8_inst : DFFR_X1 port map( D => n_state_sqrt_8_port, CK => 
                           clk, RN => rst, Q => c_state_sqrt_8_port, QN => 
                           net108017);
   c_state_sqrt_reg_9_inst : DFFR_X1 port map( D => n_state_sqrt_9_port, CK => 
                           clk, RN => rst, Q => c_state_sqrt_9_port, QN => n271
                           );
   c_state_sqrt_reg_11_inst : DFFR_X1 port map( D => n_state_sqrt_11_port, CK 
                           => clk, RN => rst, Q => c_state_sqrt_11_port, QN => 
                           net108016);
   c_state_sqrt_reg_12_inst : DFFR_X1 port map( D => n_state_sqrt_12_port, CK 
                           => clk, RN => rst, Q => c_state_sqrt_12_port, QN => 
                           net108015);
   c_state_sqrt_reg_13_inst : DFFR_X1 port map( D => n_state_sqrt_13_port, CK 
                           => clk, RN => rst, Q => c_state_sqrt_13_port, QN => 
                           n239);
   c_state_sqrt_reg_14_inst : DFFR_X1 port map( D => n_state_sqrt_14_port, CK 
                           => clk, RN => rst, Q => c_state_sqrt_14_port, QN => 
                           n238);
   c_state_sqrt_reg_15_inst : DFFR_X1 port map( D => n_state_sqrt_15_port, CK 
                           => clk, RN => rst, Q => c_state_sqrt_15_port, QN => 
                           n237);
   c_state_sqrt_reg_16_inst : DFFR_X1 port map( D => n_state_sqrt_16_port, CK 
                           => clk, RN => rst, Q => c_state_sqrt_16_port, QN => 
                           net108014);
   c_state_sqrt_reg_17_inst : DFFR_X1 port map( D => n_state_sqrt_17_port, CK 
                           => clk, RN => rst, Q => c_state_sqrt_17_port, QN => 
                           net108013);
   c_state_sqrt_reg_18_inst : DFFR_X1 port map( D => n_state_sqrt_18_port, CK 
                           => clk, RN => rst, Q => c_state_sqrt_18_port, QN => 
                           net108012);
   c_state_sqrt_reg_19_inst : DFFR_X1 port map( D => n_state_sqrt_19_port, CK 
                           => clk, RN => rst, Q => c_state_sqrt_19_port, QN => 
                           n236);
   c_state_sqrt_reg_20_inst : DFFR_X1 port map( D => n_state_sqrt_20_port, CK 
                           => clk, RN => rst, Q => c_state_sqrt_20_port, QN => 
                           n235);
   c_state_sqrt_reg_21_inst : DFFR_X1 port map( D => n_state_sqrt_21_port, CK 
                           => clk, RN => rst, Q => c_state_sqrt_21_port, QN => 
                           n234);
   c_state_sqrt_reg_22_inst : DFFR_X1 port map( D => n_state_sqrt_22_port, CK 
                           => clk, RN => rst, Q => c_state_sqrt_22_port, QN => 
                           net108011);
   c_state_sqrt_reg_23_inst : DFFR_X1 port map( D => n_state_sqrt_23_port, CK 
                           => clk, RN => rst, Q => c_state_sqrt_23_port, QN => 
                           net108010);
   c_state_sqrt_reg_24_inst : DFFR_X1 port map( D => n_state_sqrt_24_port, CK 
                           => clk, RN => rst, Q => c_state_sqrt_24_port, QN => 
                           net108009);
   c_state_sqrt_reg_25_inst : DFFR_X1 port map( D => n_state_sqrt_25_port, CK 
                           => clk, RN => rst, Q => c_state_sqrt_25_port, QN => 
                           n233);
   c_state_sqrt_reg_26_inst : DFFR_X1 port map( D => n_state_sqrt_26_port, CK 
                           => clk, RN => rst, Q => c_state_sqrt_26_port, QN => 
                           n229);
   c_state_sqrt_reg_27_inst : DFFR_X1 port map( D => n_state_sqrt_27_port, CK 
                           => clk, RN => rst, Q => c_state_sqrt_27_port, QN => 
                           net108008);
   c_state_sqrt_reg_28_inst : DFFR_X1 port map( D => n_state_sqrt_28_port, CK 
                           => clk, RN => rst, Q => c_state_sqrt_28_port, QN => 
                           n261);
   c_state_sqrt_reg_29_inst : DFFR_X1 port map( D => n_state_sqrt_29_port, CK 
                           => clk, RN => rst, Q => c_state_sqrt_29_port, QN => 
                           n262);
   c_state_sqrt_reg_30_inst : DFFR_X1 port map( D => n_state_sqrt_30_port, CK 
                           => clk, RN => rst, Q => c_state_sqrt_30_port, QN => 
                           n264);
   c_state_sqrt_reg_31_inst : DFFR_X1 port map( D => n_state_sqrt_31_port, CK 
                           => clk, RN => rst, Q => c_state_sqrt_31_port, QN => 
                           net108007);
   c_state_stu_reg_0_inst : DFFR_X1 port map( D => n_state_stu_0_port, CK => 
                           clk, RN => rst, Q => c_state_stu_0_port, QN => n192)
                           ;
   c_state_stu_reg_31_inst : DFFR_X1 port map( D => n_state_stu_31_port, CK => 
                           clk, RN => rst, Q => c_state_stu_31_port, QN => n228
                           );
   c_state_stu_reg_2_inst : DFFR_X1 port map( D => n_state_stu_2_port, CK => 
                           clk, RN => rst, Q => c_state_stu_2_port, QN => 
                           n214_port);
   c_state_stu_reg_9_inst : DFFR_X1 port map( D => n_state_stu_9_port, CK => 
                           clk, RN => rst, Q => c_state_stu_9_port, QN => 
                           net108006);
   c_state_stu_reg_8_inst : DFFR_X1 port map( D => n_state_stu_8_port, CK => 
                           clk, RN => rst, Q => c_state_stu_8_port, QN => 
                           net108005);
   c_state_stu_reg_7_inst : DFFR_X1 port map( D => n_state_stu_7_port, CK => 
                           clk, RN => rst, Q => c_state_stu_7_port, QN => 
                           net108004);
   c_state_stu_reg_6_inst : DFFR_X1 port map( D => n_state_stu_6_port, CK => 
                           clk, RN => rst, Q => c_state_stu_6_port, QN => n227)
                           ;
   c_state_stu_reg_5_inst : DFFR_X1 port map( D => n_state_stu_5_port, CK => 
                           clk, RN => rst, Q => c_state_stu_5_port, QN => n226)
                           ;
   c_state_stu_reg_4_inst : DFFR_X1 port map( D => n_state_stu_4_port, CK => 
                           clk, RN => rst, Q => c_state_stu_4_port, QN => n225)
                           ;
   c_state_stu_reg_3_inst : DFFR_X1 port map( D => n_state_stu_3_port, CK => 
                           clk, RN => rst, Q => c_state_stu_3_port, QN => 
                           n224_port);
   c_state_stu_reg_30_inst : DFFR_X1 port map( D => n_state_stu_30_port, CK => 
                           clk, RN => rst, Q => c_state_stu_30_port, QN => 
                           net108003);
   c_state_stu_reg_29_inst : DFFR_X1 port map( D => n_state_stu_29_port, CK => 
                           clk, RN => rst, Q => c_state_stu_29_port, QN => 
                           net108002);
   c_state_stu_reg_28_inst : DFFR_X1 port map( D => n_state_stu_28_port, CK => 
                           clk, RN => rst, Q => c_state_stu_28_port, QN => 
                           net108001);
   c_state_stu_reg_27_inst : DFFR_X1 port map( D => n_state_stu_27_port, CK => 
                           clk, RN => rst, Q => c_state_stu_27_port, QN => 
                           n223_port);
   c_state_stu_reg_26_inst : DFFR_X1 port map( D => n_state_stu_26_port, CK => 
                           clk, RN => rst, Q => c_state_stu_26_port, QN => 
                           n221_port);
   c_state_stu_reg_25_inst : DFFR_X1 port map( D => n_state_stu_25_port, CK => 
                           clk, RN => rst, Q => c_state_stu_25_port, QN => 
                           n220_port);
   c_state_stu_reg_24_inst : DFFR_X1 port map( D => n_state_stu_24_port, CK => 
                           clk, RN => rst, Q => c_state_stu_24_port, QN => 
                           n219_port);
   c_state_stu_reg_23_inst : DFFR_X1 port map( D => n_state_stu_23_port, CK => 
                           clk, RN => rst, Q => c_state_stu_23_port, QN => 
                           net108000);
   c_state_stu_reg_22_inst : DFFR_X1 port map( D => n_state_stu_22_port, CK => 
                           clk, RN => rst, Q => c_state_stu_22_port, QN => 
                           net107999);
   c_state_stu_reg_21_inst : DFFR_X1 port map( D => n_state_stu_21_port, CK => 
                           clk, RN => rst, Q => c_state_stu_21_port, QN => 
                           net107998);
   c_state_stu_reg_20_inst : DFFR_X1 port map( D => n_state_stu_20_port, CK => 
                           clk, RN => rst, Q => c_state_stu_20_port, QN => 
                           n218_port);
   c_state_stu_reg_1_inst : DFFR_X1 port map( D => n_state_stu_1_port, CK => 
                           clk, RN => rst, Q => c_state_stu_1_port, QN => 
                           n194_port);
   c_state_stu_reg_19_inst : DFFR_X1 port map( D => n_state_stu_19_port, CK => 
                           clk, RN => rst, Q => c_state_stu_19_port, QN => 
                           n217_port);
   c_state_stu_reg_18_inst : DFFR_X1 port map( D => n_state_stu_18_port, CK => 
                           clk, RN => rst, Q => c_state_stu_18_port, QN => 
                           n216_port);
   c_state_stu_reg_17_inst : DFFR_X1 port map( D => n_state_stu_17_port, CK => 
                           clk, RN => rst, Q => c_state_stu_17_port, QN => 
                           n215_port);
   c_state_stu_reg_16_inst : DFFR_X1 port map( D => n_state_stu_16_port, CK => 
                           clk, RN => rst, Q => c_state_stu_16_port, QN => 
                           net107997);
   c_state_stu_reg_15_inst : DFFR_X1 port map( D => n_state_stu_15_port, CK => 
                           clk, RN => rst, Q => c_state_stu_15_port, QN => 
                           net107996);
   c_state_stu_reg_14_inst : DFFR_X1 port map( D => n_state_stu_14_port, CK => 
                           clk, RN => rst, Q => c_state_stu_14_port, QN => 
                           net107995);
   c_state_stu_reg_13_inst : DFFR_X1 port map( D => n_state_stu_13_port, CK => 
                           clk, RN => rst, Q => c_state_stu_13_port, QN => 
                           n213_port);
   c_state_stu_reg_12_inst : DFFR_X1 port map( D => n_state_stu_12_port, CK => 
                           clk, RN => rst, Q => c_state_stu_12_port, QN => 
                           n212_port);
   c_state_stu_reg_11_inst : DFFR_X1 port map( D => n_state_stu_11_port, CK => 
                           clk, RN => rst, Q => c_state_stu_11_port, QN => 
                           n211_port);
   c_state_stu_reg_10_inst : DFFR_X1 port map( D => n_state_stu_10_port, CK => 
                           clk, RN => rst, Q => c_state_stu_10_port, QN => 
                           n210_port);
   add_319 : StallGenerator_CWRD_SIZE20_DW01_inc_0 port map( A(31) => 
                           c_state_stu_31_port, A(30) => c_state_stu_30_port, 
                           A(29) => c_state_stu_29_port, A(28) => 
                           c_state_stu_28_port, A(27) => c_state_stu_27_port, 
                           A(26) => c_state_stu_26_port, A(25) => 
                           c_state_stu_25_port, A(24) => c_state_stu_24_port, 
                           A(23) => c_state_stu_23_port, A(22) => 
                           c_state_stu_22_port, A(21) => c_state_stu_21_port, 
                           A(20) => c_state_stu_20_port, A(19) => 
                           c_state_stu_19_port, A(18) => c_state_stu_18_port, 
                           A(17) => c_state_stu_17_port, A(16) => 
                           c_state_stu_16_port, A(15) => c_state_stu_15_port, 
                           A(14) => c_state_stu_14_port, A(13) => 
                           c_state_stu_13_port, A(12) => c_state_stu_12_port, 
                           A(11) => c_state_stu_11_port, A(10) => 
                           c_state_stu_10_port, A(9) => c_state_stu_9_port, 
                           A(8) => c_state_stu_8_port, A(7) => 
                           c_state_stu_7_port, A(6) => c_state_stu_6_port, A(5)
                           => c_state_stu_5_port, A(4) => c_state_stu_4_port, 
                           A(3) => c_state_stu_3_port, A(2) => 
                           c_state_stu_2_port, A(1) => c_state_stu_1_port, A(0)
                           => c_state_stu_0_port, SUM(31) => N475, SUM(30) => 
                           N474, SUM(29) => N473, SUM(28) => N472, SUM(27) => 
                           N471, SUM(26) => N470, SUM(25) => N469, SUM(24) => 
                           N468, SUM(23) => N467, SUM(22) => N466, SUM(21) => 
                           N465, SUM(20) => N464, SUM(19) => N463, SUM(18) => 
                           N462, SUM(17) => N461, SUM(16) => N460, SUM(15) => 
                           N459, SUM(14) => N458, SUM(13) => N457, SUM(12) => 
                           N456, SUM(11) => N455, SUM(10) => N454, SUM(9) => 
                           N453, SUM(8) => N452, SUM(7) => N451, SUM(6) => N450
                           , SUM(5) => N449, SUM(4) => N448, SUM(3) => N447, 
                           SUM(2) => N446, SUM(1) => N445, SUM(0) => N444);
   add_277 : StallGenerator_CWRD_SIZE20_DW01_inc_1 port map( A(31) => 
                           c_state_sqrt_31_port, A(30) => c_state_sqrt_30_port,
                           A(29) => c_state_sqrt_29_port, A(28) => 
                           c_state_sqrt_28_port, A(27) => c_state_sqrt_27_port,
                           A(26) => c_state_sqrt_26_port, A(25) => 
                           c_state_sqrt_25_port, A(24) => c_state_sqrt_24_port,
                           A(23) => c_state_sqrt_23_port, A(22) => 
                           c_state_sqrt_22_port, A(21) => c_state_sqrt_21_port,
                           A(20) => c_state_sqrt_20_port, A(19) => 
                           c_state_sqrt_19_port, A(18) => c_state_sqrt_18_port,
                           A(17) => c_state_sqrt_17_port, A(16) => 
                           c_state_sqrt_16_port, A(15) => c_state_sqrt_15_port,
                           A(14) => c_state_sqrt_14_port, A(13) => 
                           c_state_sqrt_13_port, A(12) => c_state_sqrt_12_port,
                           A(11) => c_state_sqrt_11_port, A(10) => 
                           c_state_sqrt_10_port, A(9) => c_state_sqrt_9_port, 
                           A(8) => c_state_sqrt_8_port, A(7) => 
                           c_state_sqrt_7_port, A(6) => c_state_sqrt_6_port, 
                           A(5) => c_state_sqrt_5_port, A(4) => 
                           c_state_sqrt_4_port, A(3) => c_state_sqrt_3_port, 
                           A(2) => c_state_sqrt_2_port, A(1) => 
                           c_state_sqrt_1_port, A(0) => c_state_sqrt_0_port, 
                           SUM(31) => N394, SUM(30) => N393, SUM(29) => N392, 
                           SUM(28) => N391, SUM(27) => N390, SUM(26) => N389, 
                           SUM(25) => N388, SUM(24) => N387, SUM(23) => N386, 
                           SUM(22) => N385, SUM(21) => N384, SUM(20) => N383, 
                           SUM(19) => N382, SUM(18) => N381, SUM(17) => N380, 
                           SUM(16) => N379, SUM(15) => N378, SUM(14) => N377, 
                           SUM(13) => N376, SUM(12) => N375, SUM(11) => N374, 
                           SUM(10) => N373, SUM(9) => N372, SUM(8) => N371, 
                           SUM(7) => N370, SUM(6) => N369, SUM(5) => N368, 
                           SUM(4) => N367, SUM(3) => N366, SUM(2) => N365, 
                           SUM(1) => N364, SUM(0) => N363);
   add_232 : StallGenerator_CWRD_SIZE20_DW01_inc_2 port map( A(31) => 
                           c_state_div_31_port, A(30) => c_state_div_30_port, 
                           A(29) => c_state_div_29_port, A(28) => 
                           c_state_div_28_port, A(27) => c_state_div_27_port, 
                           A(26) => c_state_div_26_port, A(25) => 
                           c_state_div_25_port, A(24) => c_state_div_24_port, 
                           A(23) => c_state_div_23_port, A(22) => 
                           c_state_div_22_port, A(21) => c_state_div_21_port, 
                           A(20) => c_state_div_20_port, A(19) => 
                           c_state_div_19_port, A(18) => c_state_div_18_port, 
                           A(17) => c_state_div_17_port, A(16) => 
                           c_state_div_16_port, A(15) => c_state_div_15_port, 
                           A(14) => c_state_div_14_port, A(13) => 
                           c_state_div_13_port, A(12) => c_state_div_12_port, 
                           A(11) => c_state_div_11_port, A(10) => 
                           c_state_div_10_port, A(9) => c_state_div_9_port, 
                           A(8) => c_state_div_8_port, A(7) => 
                           c_state_div_7_port, A(6) => c_state_div_6_port, A(5)
                           => c_state_div_5_port, A(4) => c_state_div_4_port, 
                           A(3) => c_state_div_3_port, A(2) => 
                           c_state_div_2_port, A(1) => c_state_div_1_port, A(0)
                           => c_state_div_0_port, SUM(31) => N309, SUM(30) => 
                           N308, SUM(29) => N307, SUM(28) => N306, SUM(27) => 
                           N305, SUM(26) => N304, SUM(25) => N303, SUM(24) => 
                           N302, SUM(23) => N301, SUM(22) => N300, SUM(21) => 
                           N299, SUM(20) => N298, SUM(19) => N297, SUM(18) => 
                           N296, SUM(17) => N295, SUM(16) => N294, SUM(15) => 
                           N293, SUM(14) => N292, SUM(13) => N291, SUM(12) => 
                           N290, SUM(11) => N289, SUM(10) => N288, SUM(9) => 
                           N287, SUM(8) => N286, SUM(7) => N285, SUM(6) => N284
                           , SUM(5) => N283, SUM(4) => N282, SUM(3) => N281, 
                           SUM(2) => N280, SUM(1) => N279, SUM(0) => N278);
   add_187 : StallGenerator_CWRD_SIZE20_DW01_inc_3 port map( A(31) => 
                           c_state_mul_31_port, A(30) => c_state_mul_30_port, 
                           A(29) => c_state_mul_29_port, A(28) => 
                           c_state_mul_28_port, A(27) => c_state_mul_27_port, 
                           A(26) => c_state_mul_26_port, A(25) => 
                           c_state_mul_25_port, A(24) => c_state_mul_24_port, 
                           A(23) => c_state_mul_23_port, A(22) => 
                           c_state_mul_22_port, A(21) => c_state_mul_21_port, 
                           A(20) => c_state_mul_20_port, A(19) => 
                           c_state_mul_19_port, A(18) => c_state_mul_18_port, 
                           A(17) => c_state_mul_17_port, A(16) => 
                           c_state_mul_16_port, A(15) => c_state_mul_15_port, 
                           A(14) => c_state_mul_14_port, A(13) => 
                           c_state_mul_13_port, A(12) => c_state_mul_12_port, 
                           A(11) => c_state_mul_11_port, A(10) => 
                           c_state_mul_10_port, A(9) => c_state_mul_9_port, 
                           A(8) => c_state_mul_8_port, A(7) => 
                           c_state_mul_7_port, A(6) => c_state_mul_6_port, A(5)
                           => c_state_mul_5_port, A(4) => c_state_mul_4_port, 
                           A(3) => c_state_mul_3_port, A(2) => 
                           c_state_mul_2_port, A(1) => c_state_mul_1_port, A(0)
                           => c_state_mul_0_port, SUM(31) => N224, SUM(30) => 
                           N223, SUM(29) => N222, SUM(28) => N221, SUM(27) => 
                           N220, SUM(26) => N219, SUM(25) => N218, SUM(24) => 
                           N217, SUM(23) => N216, SUM(22) => N215, SUM(21) => 
                           N214, SUM(20) => N213, SUM(19) => N212, SUM(18) => 
                           N211, SUM(17) => N210, SUM(16) => N209, SUM(15) => 
                           N208, SUM(14) => N207, SUM(13) => N206, SUM(12) => 
                           N205, SUM(11) => N204, SUM(10) => N203, SUM(9) => 
                           N202, SUM(8) => N201, SUM(7) => N200, SUM(6) => N199
                           , SUM(5) => N198, SUM(4) => N197, SUM(3) => N196, 
                           SUM(2) => N195, SUM(1) => N194, SUM(0) => N193);
   add_109 : StallGenerator_CWRD_SIZE20_DW01_inc_4 port map( A(31) => 
                           c_state_bpw_31_port, A(30) => c_state_bpw_30_port, 
                           A(29) => c_state_bpw_29_port, A(28) => 
                           c_state_bpw_28_port, A(27) => c_state_bpw_27_port, 
                           A(26) => c_state_bpw_26_port, A(25) => 
                           c_state_bpw_25_port, A(24) => c_state_bpw_24_port, 
                           A(23) => c_state_bpw_23_port, A(22) => 
                           c_state_bpw_22_port, A(21) => c_state_bpw_21_port, 
                           A(20) => c_state_bpw_20_port, A(19) => 
                           c_state_bpw_19_port, A(18) => c_state_bpw_18_port, 
                           A(17) => c_state_bpw_17_port, A(16) => 
                           c_state_bpw_16_port, A(15) => c_state_bpw_15_port, 
                           A(14) => c_state_bpw_14_port, A(13) => 
                           c_state_bpw_13_port, A(12) => c_state_bpw_12_port, 
                           A(11) => c_state_bpw_11_port, A(10) => 
                           c_state_bpw_10_port, A(9) => c_state_bpw_9_port, 
                           A(8) => c_state_bpw_8_port, A(7) => 
                           c_state_bpw_7_port, A(6) => c_state_bpw_6_port, A(5)
                           => c_state_bpw_5_port, A(4) => c_state_bpw_4_port, 
                           A(3) => c_state_bpw_3_port, A(2) => 
                           c_state_bpw_2_port, A(1) => c_state_bpw_1_port, A(0)
                           => c_state_bpw_0_port, SUM(31) => N150, SUM(30) => 
                           N149, SUM(29) => N148, SUM(28) => N147, SUM(27) => 
                           N146, SUM(26) => N145, SUM(25) => N144, SUM(24) => 
                           N143, SUM(23) => N142, SUM(22) => N141, SUM(21) => 
                           N140, SUM(20) => N139, SUM(19) => N138, SUM(18) => 
                           N137, SUM(17) => N136, SUM(16) => N135, SUM(15) => 
                           N134, SUM(14) => N133, SUM(13) => N132, SUM(12) => 
                           N131, SUM(11) => N130, SUM(10) => N129, SUM(9) => 
                           N128, SUM(8) => N127, SUM(7) => N126, SUM(6) => N125
                           , SUM(5) => N124, SUM(4) => N123, SUM(3) => N122, 
                           SUM(2) => N121, SUM(1) => N120, SUM(0) => N119);
   add_69 : StallGenerator_CWRD_SIZE20_DW01_inc_5 port map( A(31) => 
                           c_state_ral_31_port, A(30) => c_state_ral_30_port, 
                           A(29) => c_state_ral_29_port, A(28) => 
                           c_state_ral_28_port, A(27) => c_state_ral_27_port, 
                           A(26) => c_state_ral_26_port, A(25) => 
                           c_state_ral_25_port, A(24) => c_state_ral_24_port, 
                           A(23) => c_state_ral_23_port, A(22) => 
                           c_state_ral_22_port, A(21) => c_state_ral_21_port, 
                           A(20) => c_state_ral_20_port, A(19) => 
                           c_state_ral_19_port, A(18) => c_state_ral_18_port, 
                           A(17) => c_state_ral_17_port, A(16) => 
                           c_state_ral_16_port, A(15) => c_state_ral_15_port, 
                           A(14) => c_state_ral_14_port, A(13) => 
                           c_state_ral_13_port, A(12) => c_state_ral_12_port, 
                           A(11) => c_state_ral_11_port, A(10) => 
                           c_state_ral_10_port, A(9) => c_state_ral_9_port, 
                           A(8) => c_state_ral_8_port, A(7) => 
                           c_state_ral_7_port, A(6) => c_state_ral_6_port, A(5)
                           => c_state_ral_5_port, A(4) => c_state_ral_4_port, 
                           A(3) => c_state_ral_3_port, A(2) => 
                           c_state_ral_2_port, A(1) => c_state_ral_1_port, A(0)
                           => c_state_ral_0_port, SUM(31) => N77, SUM(30) => 
                           N76, SUM(29) => N75, SUM(28) => N74, SUM(27) => N73,
                           SUM(26) => N72, SUM(25) => N71, SUM(24) => N70, 
                           SUM(23) => N69, SUM(22) => N68, SUM(21) => N67, 
                           SUM(20) => N66, SUM(19) => N65, SUM(18) => N64, 
                           SUM(17) => N63, SUM(16) => N62, SUM(15) => N61, 
                           SUM(14) => N60, SUM(13) => N59, SUM(12) => N58, 
                           SUM(11) => N57, SUM(10) => N56, SUM(9) => N55, 
                           SUM(8) => N54, SUM(7) => N53, SUM(6) => N52, SUM(5) 
                           => N51, SUM(4) => N50, SUM(3) => N49, SUM(2) => N48,
                           SUM(1) => N47, SUM(0) => N46);
   U3 : OAI21_X4 port map( B1 => n67_port, B2 => n50_port, A => n228, ZN => 
                           n65_port);
   U4 : OR2_X1 port map( A1 => sig_jral, A2 => n1, ZN => stall_flag_3_port);
   U5 : NAND3_X1 port map( A1 => n2, A2 => n3, A3 => n4, ZN => 
                           stall_flag_2_port);
   U6 : INV_X1 port map( A => n1, ZN => n4);
   U7 : NAND3_X1 port map( A1 => n5, A2 => n6, A3 => n7, ZN => n1);
   U8 : AND3_X1 port map( A1 => n8, A2 => n9, A3 => n10, ZN => n7);
   U9 : INV_X1 port map( A => n11, ZN => n5);
   U10 : NAND4_X1 port map( A1 => n12, A2 => n2, A3 => n13, A4 => n14, ZN => 
                           stall_flag_1_port);
   U11 : AOI211_X1 port map( C1 => n15, C2 => c_state_div_0_port, A => n16, B 
                           => n11, ZN => n14);
   U12 : OAI221_X1 port map( B1 => n17, B2 => n18, C1 => n2, C2 => 
                           c_state_stu_0_port, A => n19, ZN => n11);
   U13 : AOI22_X1 port map( A1 => n20, A2 => n21, B1 => n22, B2 => n23, ZN => 
                           n19);
   U14 : OAI21_X1 port map( B1 => n24, B2 => c_state_mul_3_port, A => n25, ZN 
                           => n22);
   U15 : OAI21_X1 port map( B1 => n26, B2 => c_state_sqrt_4_port, A => n27, ZN 
                           => n20);
   U16 : INV_X1 port map( A => n28, ZN => n27);
   U17 : AOI21_X1 port map( B1 => n230, B2 => n15, A => n29, ZN => n18);
   U18 : OAI22_X1 port map( A1 => n294_port, A2 => n24, B1 => n247, B2 => n26, 
                           ZN => n16);
   U19 : INV_X1 port map( A => n30, ZN => n24);
   U20 : AOI22_X1 port map( A1 => n31, A2 => n232, B1 => n192, B2 => n32, ZN =>
                           n13);
   U21 : NOR2_X1 port map( A1 => n197_port, A2 => n33, ZN => n31);
   U22 : NAND2_X1 port map( A1 => n194_port, A2 => n32, ZN => n2);
   U23 : OR3_X1 port map( A1 => n34, A2 => n195_port, A3 => c_state_ral_1_port,
                           ZN => n12);
   U24 : NAND4_X1 port map( A1 => n35, A2 => n36, A3 => n37, A4 => n38, ZN => 
                           stall_flag_0_port);
   U25 : NOR3_X1 port map( A1 => n39, A2 => n40, A3 => n41, ZN => n38);
   U26 : NOR3_X1 port map( A1 => n29, A2 => n32, A3 => n42, ZN => n37);
   U27 : INV_X1 port map( A => n25, ZN => n42);
   U28 : NAND3_X1 port map( A1 => n312, A2 => n43, A3 => n44, ZN => n25);
   U29 : MUX2_X1 port map( A => n45, B => n46_port, S => c_state_mul_3_port, Z 
                           => n44);
   U30 : AND2_X1 port map( A1 => n294_port, A2 => n47_port, ZN => n46_port);
   U31 : INV_X1 port map( A => n48_port, ZN => n43);
   U32 : AND3_X1 port map( A1 => n214_port, A2 => n49_port, A3 => n228, ZN => 
                           n32);
   U33 : INV_X1 port map( A => n50_port, ZN => n49_port);
   U34 : AND2_X1 port map( A1 => n51_port, A2 => n52_port, ZN => n29);
   U35 : MUX2_X1 port map( A => n53_port, B => n54_port, S => 
                           c_state_div_5_port, Z => n51_port);
   U36 : NOR2_X1 port map( A1 => c_state_div_0_port, A2 => n53_port, ZN => 
                           n54_port);
   U37 : AOI221_X1 port map( B1 => n55_port, B2 => n197_port, C1 => n56_port, 
                           C2 => n195_port, A => n28, ZN => n36);
   U38 : NOR3_X1 port map( A1 => c_state_sqrt_31_port, A2 => n57_port, A3 => 
                           n58_port, ZN => n28);
   U39 : INV_X1 port map( A => n59_port, ZN => n58_port);
   U40 : MUX2_X1 port map( A => n60_port, B => n61_port, S => 
                           c_state_sqrt_4_port, Z => n59_port);
   U41 : NOR2_X1 port map( A1 => c_state_sqrt_0_port, A2 => n60_port, ZN => 
                           n61_port);
   U42 : NOR2_X1 port map( A1 => n231, A2 => n34, ZN => n56_port);
   U43 : INV_X1 port map( A => n62_port, ZN => n34);
   U44 : NOR2_X1 port map( A1 => n232, A2 => n33, ZN => n55_port);
   U45 : INV_X1 port map( A => n63_port, ZN => n33);
   U46 : AOI222_X1 port map( A1 => n15, A2 => c_state_div_5_port, B1 => 
                           n64_port, B2 => c_state_sqrt_4_port, C1 => n30, C2 
                           => c_state_mul_3_port, ZN => n35);
   U47 : AND2_X1 port map( A1 => N453, A2 => n65_port, ZN => n_state_stu_9_port
                           );
   U48 : AND2_X1 port map( A1 => N452, A2 => n65_port, ZN => n_state_stu_8_port
                           );
   U49 : AND2_X1 port map( A1 => N451, A2 => n65_port, ZN => n_state_stu_7_port
                           );
   U50 : AND2_X1 port map( A1 => N450, A2 => n65_port, ZN => n_state_stu_6_port
                           );
   U51 : AND2_X1 port map( A1 => N449, A2 => n65_port, ZN => n_state_stu_5_port
                           );
   U52 : AND2_X1 port map( A1 => N448, A2 => n65_port, ZN => n_state_stu_4_port
                           );
   U53 : AND2_X1 port map( A1 => N447, A2 => n65_port, ZN => n_state_stu_3_port
                           );
   U54 : AND2_X1 port map( A1 => N475, A2 => n65_port, ZN => 
                           n_state_stu_31_port);
   U55 : AND2_X1 port map( A1 => N474, A2 => n65_port, ZN => 
                           n_state_stu_30_port);
   U56 : OR2_X1 port map( A1 => n66_port, A2 => N446, ZN => n_state_stu_2_port)
                           ;
   U57 : AND2_X1 port map( A1 => N473, A2 => n65_port, ZN => 
                           n_state_stu_29_port);
   U58 : AND2_X1 port map( A1 => N472, A2 => n65_port, ZN => 
                           n_state_stu_28_port);
   U59 : AND2_X1 port map( A1 => N471, A2 => n65_port, ZN => 
                           n_state_stu_27_port);
   U60 : AND2_X1 port map( A1 => N470, A2 => n65_port, ZN => 
                           n_state_stu_26_port);
   U61 : AND2_X1 port map( A1 => N469, A2 => n65_port, ZN => 
                           n_state_stu_25_port);
   U62 : AND2_X1 port map( A1 => N468, A2 => n65_port, ZN => 
                           n_state_stu_24_port);
   U63 : AND2_X1 port map( A1 => N467, A2 => n65_port, ZN => 
                           n_state_stu_23_port);
   U64 : AND2_X1 port map( A1 => N466, A2 => n65_port, ZN => 
                           n_state_stu_22_port);
   U65 : AND2_X1 port map( A1 => N465, A2 => n65_port, ZN => 
                           n_state_stu_21_port);
   U66 : AND2_X1 port map( A1 => N464, A2 => n65_port, ZN => 
                           n_state_stu_20_port);
   U67 : AND2_X1 port map( A1 => N445, A2 => n65_port, ZN => n_state_stu_1_port
                           );
   U68 : AND2_X1 port map( A1 => N463, A2 => n65_port, ZN => 
                           n_state_stu_19_port);
   U69 : AND2_X1 port map( A1 => N462, A2 => n65_port, ZN => 
                           n_state_stu_18_port);
   U70 : AND2_X1 port map( A1 => N461, A2 => n65_port, ZN => 
                           n_state_stu_17_port);
   U71 : AND2_X1 port map( A1 => N460, A2 => n65_port, ZN => 
                           n_state_stu_16_port);
   U72 : AND2_X1 port map( A1 => N459, A2 => n65_port, ZN => 
                           n_state_stu_15_port);
   U73 : AND2_X1 port map( A1 => N458, A2 => n65_port, ZN => 
                           n_state_stu_14_port);
   U74 : AND2_X1 port map( A1 => N457, A2 => n65_port, ZN => 
                           n_state_stu_13_port);
   U75 : AND2_X1 port map( A1 => N456, A2 => n65_port, ZN => 
                           n_state_stu_12_port);
   U76 : AND2_X1 port map( A1 => N455, A2 => n65_port, ZN => 
                           n_state_stu_11_port);
   U77 : AND2_X1 port map( A1 => N454, A2 => n65_port, ZN => 
                           n_state_stu_10_port);
   U78 : OR2_X1 port map( A1 => n66_port, A2 => N444, ZN => n_state_stu_0_port)
                           ;
   U79 : INV_X1 port map( A => n65_port, ZN => n66_port);
   U80 : NAND4_X1 port map( A1 => n68_port, A2 => n69_port, A3 => n70_port, A4 
                           => n71_port, ZN => n50_port);
   U81 : NOR4_X1 port map( A1 => n72_port, A2 => c_state_stu_16_port, A3 => 
                           c_state_stu_14_port, A4 => c_state_stu_15_port, ZN 
                           => n71_port);
   U82 : NAND4_X1 port map( A1 => n213_port, A2 => n212_port, A3 => n211_port, 
                           A4 => n210_port, ZN => n72_port);
   U83 : NOR4_X1 port map( A1 => n73_port, A2 => c_state_stu_23_port, A3 => 
                           c_state_stu_21_port, A4 => c_state_stu_22_port, ZN 
                           => n70_port);
   U84 : NAND4_X1 port map( A1 => n218_port, A2 => n217_port, A3 => n216_port, 
                           A4 => n215_port, ZN => n73_port);
   U85 : NOR4_X1 port map( A1 => n74_port, A2 => c_state_stu_30_port, A3 => 
                           c_state_stu_28_port, A4 => c_state_stu_29_port, ZN 
                           => n69_port);
   U86 : NAND4_X1 port map( A1 => n223_port, A2 => n221_port, A3 => n220_port, 
                           A4 => n219_port, ZN => n74_port);
   U87 : NOR4_X1 port map( A1 => n75_port, A2 => c_state_stu_9_port, A3 => 
                           c_state_stu_7_port, A4 => c_state_stu_8_port, ZN => 
                           n68_port);
   U88 : NAND4_X1 port map( A1 => n227, A2 => n226, A3 => n225, A4 => n224_port
                           , ZN => n75_port);
   U89 : AOI21_X1 port map( B1 => n192, B2 => n194_port, A => n214_port, ZN => 
                           n67_port);
   U90 : AND2_X1 port map( A1 => N372, A2 => n76_port, ZN => 
                           n_state_sqrt_9_port);
   U91 : AND2_X1 port map( A1 => N371, A2 => n76_port, ZN => 
                           n_state_sqrt_8_port);
   U92 : AND2_X1 port map( A1 => N370, A2 => n76_port, ZN => 
                           n_state_sqrt_7_port);
   U93 : AND2_X1 port map( A1 => N369, A2 => n76_port, ZN => 
                           n_state_sqrt_6_port);
   U94 : AND2_X1 port map( A1 => N368, A2 => n76_port, ZN => 
                           n_state_sqrt_5_port);
   U95 : AND2_X1 port map( A1 => N367, A2 => n76_port, ZN => 
                           n_state_sqrt_4_port);
   U96 : AND2_X1 port map( A1 => N366, A2 => n76_port, ZN => 
                           n_state_sqrt_3_port);
   U97 : AND2_X1 port map( A1 => N394, A2 => n76_port, ZN => 
                           n_state_sqrt_31_port);
   U98 : AND2_X1 port map( A1 => N393, A2 => n76_port, ZN => 
                           n_state_sqrt_30_port);
   U99 : AND2_X1 port map( A1 => N365, A2 => n76_port, ZN => 
                           n_state_sqrt_2_port);
   U100 : AND2_X1 port map( A1 => N392, A2 => n76_port, ZN => 
                           n_state_sqrt_29_port);
   U101 : AND2_X1 port map( A1 => N391, A2 => n76_port, ZN => 
                           n_state_sqrt_28_port);
   U102 : AND2_X1 port map( A1 => N390, A2 => n76_port, ZN => 
                           n_state_sqrt_27_port);
   U103 : AND2_X1 port map( A1 => N389, A2 => n76_port, ZN => 
                           n_state_sqrt_26_port);
   U104 : AND2_X1 port map( A1 => N388, A2 => n76_port, ZN => 
                           n_state_sqrt_25_port);
   U105 : AND2_X1 port map( A1 => N387, A2 => n76_port, ZN => 
                           n_state_sqrt_24_port);
   U106 : AND2_X1 port map( A1 => N386, A2 => n76_port, ZN => 
                           n_state_sqrt_23_port);
   U107 : AND2_X1 port map( A1 => N385, A2 => n76_port, ZN => 
                           n_state_sqrt_22_port);
   U108 : AND2_X1 port map( A1 => N384, A2 => n76_port, ZN => 
                           n_state_sqrt_21_port);
   U109 : AND2_X1 port map( A1 => N383, A2 => n76_port, ZN => 
                           n_state_sqrt_20_port);
   U110 : AND2_X1 port map( A1 => N364, A2 => n76_port, ZN => 
                           n_state_sqrt_1_port);
   U111 : AND2_X1 port map( A1 => N382, A2 => n76_port, ZN => 
                           n_state_sqrt_19_port);
   U112 : AND2_X1 port map( A1 => N381, A2 => n76_port, ZN => 
                           n_state_sqrt_18_port);
   U113 : AND2_X1 port map( A1 => N380, A2 => n76_port, ZN => 
                           n_state_sqrt_17_port);
   U114 : AND2_X1 port map( A1 => N379, A2 => n76_port, ZN => 
                           n_state_sqrt_16_port);
   U115 : AND2_X1 port map( A1 => N378, A2 => n76_port, ZN => 
                           n_state_sqrt_15_port);
   U116 : AND2_X1 port map( A1 => N377, A2 => n76_port, ZN => 
                           n_state_sqrt_14_port);
   U117 : AND2_X1 port map( A1 => N376, A2 => n76_port, ZN => 
                           n_state_sqrt_13_port);
   U118 : AND2_X1 port map( A1 => N375, A2 => n76_port, ZN => 
                           n_state_sqrt_12_port);
   U119 : AND2_X1 port map( A1 => N374, A2 => n76_port, ZN => 
                           n_state_sqrt_11_port);
   U120 : AND2_X1 port map( A1 => N373, A2 => n76_port, ZN => 
                           n_state_sqrt_10_port);
   U121 : INV_X1 port map( A => n77_port, ZN => n76_port);
   U122 : OAI21_X1 port map( B1 => n77_port, B2 => n78, A => n6, ZN => 
                           n_state_sqrt_0_port);
   U123 : OAI211_X1 port map( C1 => n39, C2 => n79, A => n9, B => sig_sqrt, ZN 
                           => n6);
   U124 : AND4_X1 port map( A1 => c_state_sqrt_4_port, A2 => 
                           c_state_sqrt_1_port, A3 => n80, A4 => n81, ZN => n39
                           );
   U125 : NOR3_X1 port map( A1 => c_state_sqrt_31_port, A2 => n57_port, A3 => 
                           c_state_sqrt_0_port, ZN => n81);
   U126 : INV_X1 port map( A => N363, ZN => n78);
   U127 : OAI21_X1 port map( B1 => n82, B2 => c_state_sqrt_31_port, A => n21, 
                           ZN => n77_port);
   U128 : INV_X1 port map( A => n79, ZN => n21);
   U129 : NOR3_X1 port map( A1 => n26, A2 => c_state_sqrt_0_port, A3 => 
                           c_state_sqrt_4_port, ZN => n79);
   U130 : INV_X1 port map( A => n64_port, ZN => n26);
   U131 : NOR3_X1 port map( A1 => c_state_sqrt_31_port, A2 => n57_port, A3 => 
                           n60_port, ZN => n64_port);
   U132 : AOI21_X1 port map( B1 => c_state_sqrt_4_port, B2 => n60_port, A => 
                           n57_port, ZN => n82);
   U133 : NAND4_X1 port map( A1 => n83, A2 => n84, A3 => n85, A4 => n86, ZN => 
                           n57_port);
   U134 : NOR4_X1 port map( A1 => n87, A2 => c_state_sqrt_16_port, A3 => 
                           c_state_sqrt_18_port, A4 => c_state_sqrt_17_port, ZN
                           => n86);
   U135 : NAND4_X1 port map( A1 => n236, A2 => n235, A3 => n234, A4 => n276, ZN
                           => n87);
   U136 : NOR4_X1 port map( A1 => n88, A2 => c_state_sqrt_27_port, A3 => 
                           c_state_sqrt_12_port, A4 => c_state_sqrt_11_port, ZN
                           => n85);
   U137 : NAND3_X1 port map( A1 => n238, A2 => n237, A3 => n239, ZN => n88);
   U138 : NOR4_X1 port map( A1 => n89, A2 => c_state_sqrt_8_port, A3 => 
                           c_state_sqrt_6_port, A4 => c_state_sqrt_7_port, ZN 
                           => n84);
   U139 : NAND4_X1 port map( A1 => n267, A2 => n264, A3 => n262, A4 => n261, ZN
                           => n89);
   U140 : NOR4_X1 port map( A1 => n90, A2 => c_state_sqrt_22_port, A3 => 
                           c_state_sqrt_24_port, A4 => c_state_sqrt_23_port, ZN
                           => n83);
   U141 : NAND3_X1 port map( A1 => n229, A2 => n271, A3 => n233, ZN => n90);
   U142 : NAND2_X1 port map( A1 => n240, A2 => n80, ZN => n60_port);
   U143 : AND2_X1 port map( A1 => n266, A2 => n263, ZN => n80);
   U144 : AND2_X1 port map( A1 => N55, A2 => n91, ZN => n_state_ral_9_port);
   U145 : AND2_X1 port map( A1 => N54, A2 => n91, ZN => n_state_ral_8_port);
   U146 : AND2_X1 port map( A1 => N53, A2 => n91, ZN => n_state_ral_7_port);
   U147 : AND2_X1 port map( A1 => N52, A2 => n91, ZN => n_state_ral_6_port);
   U148 : AND2_X1 port map( A1 => N51, A2 => n91, ZN => n_state_ral_5_port);
   U149 : AND2_X1 port map( A1 => N50, A2 => n91, ZN => n_state_ral_4_port);
   U150 : AND2_X1 port map( A1 => N49, A2 => n91, ZN => n_state_ral_3_port);
   U151 : AND2_X1 port map( A1 => N77, A2 => n91, ZN => n_state_ral_31_port);
   U152 : AND2_X1 port map( A1 => N76, A2 => n91, ZN => n_state_ral_30_port);
   U153 : AND2_X1 port map( A1 => N48, A2 => n91, ZN => n_state_ral_2_port);
   U154 : AND2_X1 port map( A1 => N75, A2 => n91, ZN => n_state_ral_29_port);
   U155 : AND2_X1 port map( A1 => N74, A2 => n91, ZN => n_state_ral_28_port);
   U156 : AND2_X1 port map( A1 => N73, A2 => n91, ZN => n_state_ral_27_port);
   U157 : AND2_X1 port map( A1 => N72, A2 => n91, ZN => n_state_ral_26_port);
   U158 : AND2_X1 port map( A1 => N71, A2 => n91, ZN => n_state_ral_25_port);
   U159 : AND2_X1 port map( A1 => N70, A2 => n91, ZN => n_state_ral_24_port);
   U160 : AND2_X1 port map( A1 => N69, A2 => n91, ZN => n_state_ral_23_port);
   U161 : AND2_X1 port map( A1 => N68, A2 => n91, ZN => n_state_ral_22_port);
   U162 : AND2_X1 port map( A1 => N67, A2 => n91, ZN => n_state_ral_21_port);
   U163 : AND2_X1 port map( A1 => N66, A2 => n91, ZN => n_state_ral_20_port);
   U164 : AND2_X1 port map( A1 => N47, A2 => n91, ZN => n_state_ral_1_port);
   U165 : AND2_X1 port map( A1 => N65, A2 => n91, ZN => n_state_ral_19_port);
   U166 : AND2_X1 port map( A1 => N64, A2 => n91, ZN => n_state_ral_18_port);
   U167 : AND2_X1 port map( A1 => N63, A2 => n91, ZN => n_state_ral_17_port);
   U168 : AND2_X1 port map( A1 => N62, A2 => n91, ZN => n_state_ral_16_port);
   U169 : AND2_X1 port map( A1 => N61, A2 => n91, ZN => n_state_ral_15_port);
   U170 : AND2_X1 port map( A1 => N60, A2 => n91, ZN => n_state_ral_14_port);
   U171 : AND2_X1 port map( A1 => N59, A2 => n91, ZN => n_state_ral_13_port);
   U172 : AND2_X1 port map( A1 => N58, A2 => n91, ZN => n_state_ral_12_port);
   U173 : AND2_X1 port map( A1 => N57, A2 => n91, ZN => n_state_ral_11_port);
   U174 : AND2_X1 port map( A1 => N56, A2 => n91, ZN => n_state_ral_10_port);
   U175 : AND3_X1 port map( A1 => n92, A2 => n9, A3 => n93, ZN => n91);
   U176 : NAND2_X1 port map( A1 => n9, A2 => n94, ZN => n_state_ral_0_port);
   U177 : NAND3_X1 port map( A1 => n93, A2 => n92, A3 => N46, ZN => n94);
   U178 : OAI21_X1 port map( B1 => n95, B2 => c_state_ral_1_port, A => n185, ZN
                           => n92);
   U179 : NAND2_X1 port map( A1 => n195_port, A2 => n62_port, ZN => n93);
   U180 : NOR2_X1 port map( A1 => c_state_ral_31_port, A2 => n95, ZN => 
                           n62_port);
   U181 : NAND4_X1 port map( A1 => n96, A2 => n97, A3 => n98, A4 => n99, ZN => 
                           n95);
   U182 : NOR2_X1 port map( A1 => n100, A2 => n101, ZN => n99);
   U183 : NAND4_X1 port map( A1 => n196_port, A2 => n193_port, A3 => n191, A4 
                           => n190, ZN => n101);
   U184 : NAND4_X1 port map( A1 => n189, A2 => n188, A3 => n187, A4 => n186, ZN
                           => n100);
   U185 : NOR4_X1 port map( A1 => n102, A2 => c_state_ral_16_port, A3 => 
                           c_state_ral_18_port, A4 => c_state_ral_17_port, ZN 
                           => n98);
   U186 : NAND4_X1 port map( A1 => n201_port, A2 => n200_port, A3 => n199_port,
                           A4 => n198_port, ZN => n102);
   U187 : NOR4_X1 port map( A1 => n103, A2 => c_state_ral_8_port, A3 => 
                           c_state_ral_11_port, A4 => c_state_ral_9_port, ZN =>
                           n97);
   U188 : NAND4_X1 port map( A1 => n205_port, A2 => n204_port, A3 => n203_port,
                           A4 => n202_port, ZN => n103);
   U189 : NOR4_X1 port map( A1 => n104, A2 => c_state_ral_10_port, A3 => 
                           c_state_ral_3_port, A4 => c_state_ral_2_port, ZN => 
                           n96);
   U190 : NAND4_X1 port map( A1 => n209_port, A2 => n208_port, A3 => n207_port,
                           A4 => n206_port, ZN => n104);
   U191 : AND2_X1 port map( A1 => N202, A2 => n105, ZN => n_state_mul_9_port);
   U192 : AND2_X1 port map( A1 => N201, A2 => n105, ZN => n_state_mul_8_port);
   U193 : AND2_X1 port map( A1 => N200, A2 => n105, ZN => n_state_mul_7_port);
   U194 : AND2_X1 port map( A1 => N199, A2 => n105, ZN => n_state_mul_6_port);
   U195 : AND2_X1 port map( A1 => N198, A2 => n105, ZN => n_state_mul_5_port);
   U196 : AND2_X1 port map( A1 => N197, A2 => n105, ZN => n_state_mul_4_port);
   U197 : AND2_X1 port map( A1 => N196, A2 => n105, ZN => n_state_mul_3_port);
   U198 : AND2_X1 port map( A1 => N224, A2 => n105, ZN => n_state_mul_31_port);
   U199 : AND2_X1 port map( A1 => N223, A2 => n105, ZN => n_state_mul_30_port);
   U200 : AND2_X1 port map( A1 => N195, A2 => n105, ZN => n_state_mul_2_port);
   U201 : AND2_X1 port map( A1 => N222, A2 => n105, ZN => n_state_mul_29_port);
   U202 : AND2_X1 port map( A1 => N221, A2 => n105, ZN => n_state_mul_28_port);
   U203 : AND2_X1 port map( A1 => N220, A2 => n105, ZN => n_state_mul_27_port);
   U204 : AND2_X1 port map( A1 => N219, A2 => n105, ZN => n_state_mul_26_port);
   U205 : AND2_X1 port map( A1 => N218, A2 => n105, ZN => n_state_mul_25_port);
   U206 : AND2_X1 port map( A1 => N217, A2 => n105, ZN => n_state_mul_24_port);
   U207 : AND2_X1 port map( A1 => N216, A2 => n105, ZN => n_state_mul_23_port);
   U208 : AND2_X1 port map( A1 => N215, A2 => n105, ZN => n_state_mul_22_port);
   U209 : AND2_X1 port map( A1 => N214, A2 => n105, ZN => n_state_mul_21_port);
   U210 : AND2_X1 port map( A1 => N213, A2 => n105, ZN => n_state_mul_20_port);
   U211 : AND2_X1 port map( A1 => N194, A2 => n105, ZN => n_state_mul_1_port);
   U212 : AND2_X1 port map( A1 => N212, A2 => n105, ZN => n_state_mul_19_port);
   U213 : AND2_X1 port map( A1 => N211, A2 => n105, ZN => n_state_mul_18_port);
   U214 : AND2_X1 port map( A1 => N210, A2 => n105, ZN => n_state_mul_17_port);
   U215 : AND2_X1 port map( A1 => N209, A2 => n105, ZN => n_state_mul_16_port);
   U216 : AND2_X1 port map( A1 => N208, A2 => n105, ZN => n_state_mul_15_port);
   U217 : AND2_X1 port map( A1 => N207, A2 => n105, ZN => n_state_mul_14_port);
   U218 : AND2_X1 port map( A1 => N206, A2 => n105, ZN => n_state_mul_13_port);
   U219 : AND2_X1 port map( A1 => N205, A2 => n105, ZN => n_state_mul_12_port);
   U220 : AND2_X1 port map( A1 => N204, A2 => n105, ZN => n_state_mul_11_port);
   U221 : AND2_X1 port map( A1 => N203, A2 => n105, ZN => n_state_mul_10_port);
   U222 : INV_X1 port map( A => n106, ZN => n105);
   U223 : OAI21_X1 port map( B1 => n106, B2 => n107, A => n8, ZN => 
                           n_state_mul_0_port);
   U224 : OAI211_X1 port map( C1 => n41, C2 => n108, A => n9, B => sig_mul, ZN 
                           => n8);
   U225 : INV_X1 port map( A => n23, ZN => n108);
   U226 : NOR4_X1 port map( A1 => n222_port, A2 => n163, A3 => n48_port, A4 => 
                           n109, ZN => n41);
   U227 : NAND3_X1 port map( A1 => n312, A2 => n294_port, A3 => n310, ZN => 
                           n109);
   U228 : INV_X1 port map( A => N193, ZN => n107);
   U229 : OAI21_X1 port map( B1 => n110, B2 => c_state_mul_31_port, A => n23, 
                           ZN => n106);
   U230 : NAND3_X1 port map( A1 => n30, A2 => n294_port, A3 => n222_port, ZN =>
                           n23);
   U231 : NOR3_X1 port map( A1 => c_state_mul_31_port, A2 => n111, A3 => n45, 
                           ZN => n30);
   U232 : NAND3_X1 port map( A1 => n156, A2 => n112, A3 => n47_port, ZN => n45)
                           ;
   U233 : INV_X1 port map( A => n113, ZN => n47_port);
   U234 : AOI21_X1 port map( B1 => n113, B2 => c_state_mul_3_port, A => 
                           n48_port, ZN => n110);
   U235 : NAND3_X1 port map( A1 => n114, A2 => n112, A3 => n156, ZN => n48_port
                           );
   U236 : AND2_X1 port map( A1 => n115, A2 => n116, ZN => n112);
   U237 : NOR4_X1 port map( A1 => n117, A2 => c_state_mul_17_port, A3 => 
                           c_state_mul_19_port, A4 => c_state_mul_18_port, ZN 
                           => n116);
   U238 : NAND4_X1 port map( A1 => n159, A2 => n158, A3 => n157, A4 => n323, ZN
                           => n117);
   U239 : NOR4_X1 port map( A1 => n118, A2 => c_state_mul_11_port, A3 => 
                           c_state_mul_13_port, A4 => c_state_mul_12_port, ZN 
                           => n115);
   U240 : NAND3_X1 port map( A1 => n161, A2 => n160, A3 => n162, ZN => n118);
   U241 : INV_X1 port map( A => n111, ZN => n114);
   U242 : NAND2_X1 port map( A1 => n119_port, A2 => n120_port, ZN => n111);
   U243 : NOR4_X1 port map( A1 => n121_port, A2 => c_state_mul_6_port, A3 => 
                           c_state_mul_4_port, A4 => c_state_mul_5_port, ZN => 
                           n120_port);
   U244 : NAND4_X1 port map( A1 => n311, A2 => n309_port, A3 => n308_port, A4 
                           => n307_port, ZN => n121_port);
   U245 : NOR4_X1 port map( A1 => n122_port, A2 => c_state_mul_24_port, A3 => 
                           c_state_mul_26_port, A4 => c_state_mul_25_port, ZN 
                           => n119_port);
   U246 : NAND3_X1 port map( A1 => n317, A2 => n316, A3 => n318, ZN => 
                           n122_port);
   U247 : NAND2_X1 port map( A1 => n163, A2 => n310, ZN => n113);
   U248 : AND2_X1 port map( A1 => N287, A2 => n123_port, ZN => 
                           n_state_div_9_port);
   U249 : AND2_X1 port map( A1 => N286, A2 => n123_port, ZN => 
                           n_state_div_8_port);
   U250 : AND2_X1 port map( A1 => N285, A2 => n123_port, ZN => 
                           n_state_div_7_port);
   U251 : AND2_X1 port map( A1 => N284, A2 => n123_port, ZN => 
                           n_state_div_6_port);
   U252 : AND2_X1 port map( A1 => N283, A2 => n123_port, ZN => 
                           n_state_div_5_port);
   U253 : AND2_X1 port map( A1 => N282, A2 => n123_port, ZN => 
                           n_state_div_4_port);
   U254 : AND2_X1 port map( A1 => N281, A2 => n123_port, ZN => 
                           n_state_div_3_port);
   U255 : AND2_X1 port map( A1 => N309, A2 => n123_port, ZN => 
                           n_state_div_31_port);
   U256 : AND2_X1 port map( A1 => N308, A2 => n123_port, ZN => 
                           n_state_div_30_port);
   U257 : AND2_X1 port map( A1 => N280, A2 => n123_port, ZN => 
                           n_state_div_2_port);
   U258 : AND2_X1 port map( A1 => N307, A2 => n123_port, ZN => 
                           n_state_div_29_port);
   U259 : AND2_X1 port map( A1 => N306, A2 => n123_port, ZN => 
                           n_state_div_28_port);
   U260 : AND2_X1 port map( A1 => N305, A2 => n123_port, ZN => 
                           n_state_div_27_port);
   U261 : AND2_X1 port map( A1 => N304, A2 => n123_port, ZN => 
                           n_state_div_26_port);
   U262 : AND2_X1 port map( A1 => N303, A2 => n123_port, ZN => 
                           n_state_div_25_port);
   U263 : AND2_X1 port map( A1 => N302, A2 => n123_port, ZN => 
                           n_state_div_24_port);
   U264 : AND2_X1 port map( A1 => N301, A2 => n123_port, ZN => 
                           n_state_div_23_port);
   U265 : AND2_X1 port map( A1 => N300, A2 => n123_port, ZN => 
                           n_state_div_22_port);
   U266 : AND2_X1 port map( A1 => N299, A2 => n123_port, ZN => 
                           n_state_div_21_port);
   U267 : AND2_X1 port map( A1 => N298, A2 => n123_port, ZN => 
                           n_state_div_20_port);
   U268 : AND2_X1 port map( A1 => N279, A2 => n123_port, ZN => 
                           n_state_div_1_port);
   U269 : AND2_X1 port map( A1 => N297, A2 => n123_port, ZN => 
                           n_state_div_19_port);
   U270 : AND2_X1 port map( A1 => N296, A2 => n123_port, ZN => 
                           n_state_div_18_port);
   U271 : AND2_X1 port map( A1 => N295, A2 => n123_port, ZN => 
                           n_state_div_17_port);
   U272 : AND2_X1 port map( A1 => N294, A2 => n123_port, ZN => 
                           n_state_div_16_port);
   U273 : AND2_X1 port map( A1 => N293, A2 => n123_port, ZN => 
                           n_state_div_15_port);
   U274 : AND2_X1 port map( A1 => N292, A2 => n123_port, ZN => 
                           n_state_div_14_port);
   U275 : AND2_X1 port map( A1 => N291, A2 => n123_port, ZN => 
                           n_state_div_13_port);
   U276 : AND2_X1 port map( A1 => N290, A2 => n123_port, ZN => 
                           n_state_div_12_port);
   U277 : AND2_X1 port map( A1 => N289, A2 => n123_port, ZN => 
                           n_state_div_11_port);
   U278 : AND2_X1 port map( A1 => N288, A2 => n123_port, ZN => 
                           n_state_div_10_port);
   U279 : INV_X1 port map( A => n124_port, ZN => n123_port);
   U280 : OAI21_X1 port map( B1 => n124_port, B2 => n125_port, A => n10, ZN => 
                           n_state_div_0_port);
   U281 : OAI211_X1 port map( C1 => n40, C2 => n17, A => n9, B => sig_div, ZN 
                           => n10);
   U282 : INV_X1 port map( A => sig_ral, ZN => n9);
   U283 : INV_X1 port map( A => n126_port, ZN => n17);
   U284 : AND3_X1 port map( A1 => n328, A2 => n52_port, A3 => n127_port, ZN => 
                           n40);
   U285 : NOR3_X1 port map( A1 => n128_port, A2 => n155, A3 => n230, ZN => 
                           n127_port);
   U286 : INV_X1 port map( A => N278, ZN => n125_port);
   U287 : OAI21_X1 port map( B1 => n129_port, B2 => c_state_div_31_port, A => 
                           n126_port, ZN => n124_port);
   U288 : NAND3_X1 port map( A1 => n15, A2 => n328, A3 => n230, ZN => n126_port
                           );
   U289 : NOR2_X1 port map( A1 => n53_port, A2 => n130_port, ZN => n15);
   U290 : INV_X1 port map( A => n52_port, ZN => n130_port);
   U291 : NOR2_X1 port map( A1 => c_state_div_31_port, A2 => n131_port, ZN => 
                           n52_port);
   U292 : AOI21_X1 port map( B1 => c_state_div_5_port, B2 => n53_port, A => 
                           n131_port, ZN => n129_port);
   U293 : NAND4_X1 port map( A1 => n132_port, A2 => n133_port, A3 => n134_port,
                           A4 => n135_port, ZN => n131_port);
   U294 : NOR4_X1 port map( A1 => n136_port, A2 => c_state_div_16_port, A3 => 
                           c_state_div_18_port, A4 => c_state_div_17_port, ZN 
                           => n135_port);
   U295 : NAND4_X1 port map( A1 => n245, A2 => n244, A3 => n243, A4 => n357, ZN
                           => n136_port);
   U296 : NOR4_X1 port map( A1 => n137_port, A2 => c_state_div_27_port, A3 => 
                           c_state_div_12_port, A4 => c_state_div_11_port, ZN 
                           => n134_port);
   U297 : NAND3_X1 port map( A1 => n248, A2 => n246, A3 => n249, ZN => 
                           n137_port);
   U298 : NOR4_X1 port map( A1 => n138_port, A2 => c_state_div_8_port, A3 => 
                           c_state_div_6_port, A4 => c_state_div_7_port, ZN => 
                           n133_port);
   U299 : NAND3_X1 port map( A1 => n343, A2 => n342, A3 => n345, ZN => 
                           n138_port);
   U300 : NOR4_X1 port map( A1 => n139_port, A2 => c_state_div_22_port, A3 => 
                           c_state_div_24_port, A4 => c_state_div_23_port, ZN 
                           => n132_port);
   U301 : NAND3_X1 port map( A1 => n241, A2 => n352, A3 => n242, ZN => 
                           n139_port);
   U302 : NAND2_X1 port map( A1 => n155, A2 => n140_port, ZN => n53_port);
   U303 : INV_X1 port map( A => n128_port, ZN => n140_port);
   U304 : NAND3_X1 port map( A1 => n347, A2 => n344, A3 => n348, ZN => 
                           n128_port);
   U305 : AND2_X1 port map( A1 => N128, A2 => n141_port, ZN => 
                           n_state_bpw_9_port);
   U306 : AND2_X1 port map( A1 => N127, A2 => n141_port, ZN => 
                           n_state_bpw_8_port);
   U307 : AND2_X1 port map( A1 => N126, A2 => n141_port, ZN => 
                           n_state_bpw_7_port);
   U308 : AND2_X1 port map( A1 => N125, A2 => n141_port, ZN => 
                           n_state_bpw_6_port);
   U309 : AND2_X1 port map( A1 => N124, A2 => n141_port, ZN => 
                           n_state_bpw_5_port);
   U310 : AND2_X1 port map( A1 => N123, A2 => n141_port, ZN => 
                           n_state_bpw_4_port);
   U311 : AND2_X1 port map( A1 => N122, A2 => n141_port, ZN => 
                           n_state_bpw_3_port);
   U312 : AND2_X1 port map( A1 => N150, A2 => n141_port, ZN => 
                           n_state_bpw_31_port);
   U313 : AND2_X1 port map( A1 => N149, A2 => n141_port, ZN => 
                           n_state_bpw_30_port);
   U314 : AND2_X1 port map( A1 => N121, A2 => n141_port, ZN => 
                           n_state_bpw_2_port);
   U315 : AND2_X1 port map( A1 => N148, A2 => n141_port, ZN => 
                           n_state_bpw_29_port);
   U316 : AND2_X1 port map( A1 => N147, A2 => n141_port, ZN => 
                           n_state_bpw_28_port);
   U317 : AND2_X1 port map( A1 => N146, A2 => n141_port, ZN => 
                           n_state_bpw_27_port);
   U318 : AND2_X1 port map( A1 => N145, A2 => n141_port, ZN => 
                           n_state_bpw_26_port);
   U319 : AND2_X1 port map( A1 => N144, A2 => n141_port, ZN => 
                           n_state_bpw_25_port);
   U320 : AND2_X1 port map( A1 => N143, A2 => n141_port, ZN => 
                           n_state_bpw_24_port);
   U321 : AND2_X1 port map( A1 => N142, A2 => n141_port, ZN => 
                           n_state_bpw_23_port);
   U322 : AND2_X1 port map( A1 => N141, A2 => n141_port, ZN => 
                           n_state_bpw_22_port);
   U323 : AND2_X1 port map( A1 => N140, A2 => n141_port, ZN => 
                           n_state_bpw_21_port);
   U324 : AND2_X1 port map( A1 => N139, A2 => n141_port, ZN => 
                           n_state_bpw_20_port);
   U325 : AND2_X1 port map( A1 => N120, A2 => n141_port, ZN => 
                           n_state_bpw_1_port);
   U326 : AND2_X1 port map( A1 => N138, A2 => n141_port, ZN => 
                           n_state_bpw_19_port);
   U327 : AND2_X1 port map( A1 => N137, A2 => n141_port, ZN => 
                           n_state_bpw_18_port);
   U328 : AND2_X1 port map( A1 => N136, A2 => n141_port, ZN => 
                           n_state_bpw_17_port);
   U329 : AND2_X1 port map( A1 => N135, A2 => n141_port, ZN => 
                           n_state_bpw_16_port);
   U330 : AND2_X1 port map( A1 => N134, A2 => n141_port, ZN => 
                           n_state_bpw_15_port);
   U331 : AND2_X1 port map( A1 => N133, A2 => n141_port, ZN => 
                           n_state_bpw_14_port);
   U332 : AND2_X1 port map( A1 => N132, A2 => n141_port, ZN => 
                           n_state_bpw_13_port);
   U333 : AND2_X1 port map( A1 => N131, A2 => n141_port, ZN => 
                           n_state_bpw_12_port);
   U334 : AND2_X1 port map( A1 => N130, A2 => n141_port, ZN => 
                           n_state_bpw_11_port);
   U335 : AND2_X1 port map( A1 => N129, A2 => n141_port, ZN => 
                           n_state_bpw_10_port);
   U336 : AND3_X1 port map( A1 => n142_port, A2 => n3, A3 => n143_port, ZN => 
                           n141_port);
   U337 : NAND2_X1 port map( A1 => n3, A2 => n144_port, ZN => 
                           n_state_bpw_0_port);
   U338 : NAND3_X1 port map( A1 => n143_port, A2 => n142_port, A3 => N119, ZN 
                           => n144_port);
   U339 : OAI21_X1 port map( B1 => n145_port, B2 => c_state_bpw_1_port, A => 
                           n164, ZN => n142_port);
   U340 : NAND2_X1 port map( A1 => n197_port, A2 => n63_port, ZN => n143_port);
   U341 : NOR2_X1 port map( A1 => c_state_bpw_31_port, A2 => n145_port, ZN => 
                           n63_port);
   U342 : NAND4_X1 port map( A1 => n146_port, A2 => n147_port, A3 => n148_port,
                           A4 => n149_port, ZN => n145_port);
   U343 : NOR2_X1 port map( A1 => n150_port, A2 => n151, ZN => n149_port);
   U344 : NAND4_X1 port map( A1 => n172, A2 => n171, A3 => n170, A4 => n169, ZN
                           => n151);
   U345 : NAND4_X1 port map( A1 => n168, A2 => n167, A3 => n166, A4 => n165, ZN
                           => n150_port);
   U346 : NOR4_X1 port map( A1 => n152, A2 => c_state_bpw_16_port, A3 => 
                           c_state_bpw_18_port, A4 => c_state_bpw_17_port, ZN 
                           => n148_port);
   U347 : NAND4_X1 port map( A1 => n176, A2 => n175, A3 => n174, A4 => n173, ZN
                           => n152);
   U348 : NOR4_X1 port map( A1 => n153, A2 => c_state_bpw_8_port, A3 => 
                           c_state_bpw_11_port, A4 => c_state_bpw_9_port, ZN =>
                           n147_port);
   U349 : NAND4_X1 port map( A1 => n180, A2 => n179, A3 => n178, A4 => n177, ZN
                           => n153);
   U350 : NOR4_X1 port map( A1 => n154, A2 => c_state_bpw_10_port, A3 => 
                           c_state_bpw_3_port, A4 => c_state_bpw_2_port, ZN => 
                           n146_port);
   U351 : NAND4_X1 port map( A1 => n184, A2 => n183, A3 => n182, A4 => n181, ZN
                           => n154);
   U352 : INV_X1 port map( A => sig_bpw, ZN => n3);

end SYN_stall_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity CwGenerator_DATA_SIZE32_OPCD_SIZE6_FUNC_SIZE11_CWRD_SIZE20_CALU_SIZE5 is

   port( clk, rst : in std_logic;  opcd : in std_logic_vector (5 downto 0);  
         func : in std_logic_vector (10 downto 0);  stall_flag : in 
         std_logic_vector (4 downto 0);  taken : in std_logic;  cw : out 
         std_logic_vector (19 downto 0);  calu : out std_logic_vector (4 downto
         0));

end CwGenerator_DATA_SIZE32_OPCD_SIZE6_FUNC_SIZE11_CWRD_SIZE20_CALU_SIZE5;

architecture SYN_cw_generator_arch of 
   CwGenerator_DATA_SIZE32_OPCD_SIZE6_FUNC_SIZE11_CWRD_SIZE20_CALU_SIZE5 is

   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X2
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal n4, cw_0_port, calu_4_port, calu_3_port, calu_2_port, calu_1_port, 
      calu_0_port, cw_2_port, cw_1_port, n2, n3, net107991, net107992, 
      net107993, net107994 : std_logic;

begin
   cw <= ( cw_2_port, cw_2_port, cw_2_port, cw_2_port, cw_2_port, cw_2_port, 
      cw_2_port, cw_2_port, cw_2_port, cw_2_port, cw_2_port, cw_2_port, 
      cw_2_port, cw_2_port, cw_2_port, cw_2_port, cw_2_port, cw_2_port, 
      cw_1_port, cw_0_port );
   calu <= ( calu_4_port, calu_3_port, calu_2_port, calu_1_port, calu_0_port );
   
   calu_reg_3_inst : DFF_X1 port map( D => calu_3_port, CK => clk, Q => 
                           calu_3_port, QN => net107994);
   calu_reg_2_inst : DFF_X1 port map( D => calu_2_port, CK => clk, Q => 
                           calu_2_port, QN => net107993);
   calu_reg_1_inst : DFF_X1 port map( D => calu_1_port, CK => clk, Q => 
                           calu_1_port, QN => net107992);
   calu_reg_0_inst : DFF_X1 port map( D => calu_0_port, CK => clk, Q => 
                           calu_0_port, QN => net107991);
   cw_2_port <= '0';
   calu_reg_4_inst : DFF_X2 port map( D => calu_4_port, CK => clk, Q => 
                           calu_4_port, QN => n2);
   U3 : NOR2_X1 port map( A1 => stall_flag(3), A2 => n3, ZN => n4);
   U4 : INV_X1 port map( A => taken, ZN => n3);
   U5 : CLKBUF_X3 port map( A => n4, Z => cw_1_port);
   U7 : INV_X4 port map( A => stall_flag(4), ZN => cw_0_port);

end SYN_cw_generator_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity 
   DataPath_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_OPCD_SIZE6_IMME_SIZE16_CWRD_SIZE20_CALU_SIZE5_DRCW_SIZE4 
   is

   port( clk, rst : in std_logic;  istr_addr : out std_logic_vector (31 downto 
         0);  istr_val : in std_logic_vector (31 downto 0);  ir_out, pc_out, 
         reg_a_out, ld_a_out, data_addr : out std_logic_vector (31 downto 0);  
         data_i_val : in std_logic_vector (31 downto 0);  data_o_val : out 
         std_logic_vector (31 downto 0);  cw : in std_logic_vector (19 downto 
         0);  dr_cw : out std_logic_vector (3 downto 0);  calu : in 
         std_logic_vector (4 downto 0);  sig_bal : out std_logic;  sig_bpw : in
         std_logic;  sig_jral, sig_ral, sig_mul, sig_div, sig_sqrt : out 
         std_logic);

end 
   DataPath_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_OPCD_SIZE6_IMME_SIZE16_CWRD_SIZE20_CALU_SIZE5_DRCW_SIZE4;

architecture SYN_data_path_arch of 
   DataPath_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_OPCD_SIZE6_IMME_SIZE16_CWRD_SIZE20_CALU_SIZE5_DRCW_SIZE4 
   is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X2
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component Reg_DATA_SIZE5_1
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 
            0);  dout : out std_logic_vector (4 downto 0));
   end component;
   
   component Reg_DATA_SIZE32_2
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 
            0);  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Reg_DATA_SIZE5_2
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 
            0);  dout : out std_logic_vector (4 downto 0));
   end component;
   
   component Reg_DATA_SIZE32_3
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 
            0);  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Mux_DATA_SIZE32_2
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0)
            ;  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_1
      port( reg_c, reg_f, reg_ff : in std_logic_vector (31 downto 0);  addr_c, 
            addr_f, addr_ff : in std_logic_vector (4 downto 0);  valid_f, 
            valid_ff, dirty_f, dirty_ff, en : in std_logic;  output : out 
            std_logic_vector (31 downto 0);  match_dirty_f, match_dirty_ff : 
            out std_logic);
   end component;
   
   component Reg_DATA_SIZE32_4
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 
            0);  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Reg_DATA_SIZE32_5
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 
            0);  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Reg_DATA_SIZE5_3
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 
            0);  dout : out std_logic_vector (4 downto 0));
   end component;
   
   component Reg_DATA_SIZE5_4
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 
            0);  dout : out std_logic_vector (4 downto 0));
   end component;
   
   component Reg_DATA_SIZE32_6
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 
            0);  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Reg_DATA_SIZE32_7
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 
            0);  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Mux4_DATA_SIZE32
      port( sel : in std_logic_vector (1 downto 0);  din0, din1, din2, din3 : 
            in std_logic_vector (31 downto 0);  dout : out std_logic_vector (31
            downto 0));
   end component;
   
   component Div_DATA_SIZE32_DIV_STAGE34_SQRT_STAGE18
      port( rst, clk, en, lock, sign, func : in std_logic;  a, b : in 
            std_logic_vector (31 downto 0);  o : out std_logic_vector (31 
            downto 0));
   end component;
   
   component Mul_DATA_SIZE16_STAGE10
      port( rst, clk, en, lock, sign : in std_logic;  a, b : in 
            std_logic_vector (15 downto 0);  o : out std_logic_vector (31 
            downto 0));
   end component;
   
   component Alu_DATA_SIZE32
      port( f : in std_logic_vector (4 downto 0);  a, b : in std_logic_vector 
            (31 downto 0);  o : out std_logic_vector (31 downto 0));
   end component;
   
   component Mux_DATA_SIZE32_3
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0)
            ;  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_2
      port( reg_c, reg_f, reg_ff : in std_logic_vector (31 downto 0);  addr_c, 
            addr_f, addr_ff : in std_logic_vector (4 downto 0);  valid_f, 
            valid_ff, dirty_f, dirty_ff, en : in std_logic;  output : out 
            std_logic_vector (31 downto 0);  match_dirty_f, match_dirty_ff : 
            out std_logic);
   end component;
   
   component FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_3
      port( reg_c, reg_f, reg_ff : in std_logic_vector (31 downto 0);  addr_c, 
            addr_f, addr_ff : in std_logic_vector (4 downto 0);  valid_f, 
            valid_ff, dirty_f, dirty_ff, en : in std_logic;  output : out 
            std_logic_vector (31 downto 0);  match_dirty_f, match_dirty_ff : 
            out std_logic);
   end component;
   
   component Mux_DATA_SIZE32_4
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0)
            ;  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Mux_DATA_SIZE32_5
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0)
            ;  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Reg_DATA_SIZE32_8
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 
            0);  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Reg_DATA_SIZE5_5
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 
            0);  dout : out std_logic_vector (4 downto 0));
   end component;
   
   component Reg_DATA_SIZE5_6
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 
            0);  dout : out std_logic_vector (4 downto 0));
   end component;
   
   component Reg_DATA_SIZE5_0
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (4 downto 
            0);  dout : out std_logic_vector (4 downto 0));
   end component;
   
   component Reg_DATA_SIZE32_9
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 
            0);  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Reg_DATA_SIZE32_10
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 
            0);  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Reg_DATA_SIZE32_11
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 
            0);  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_4
      port( reg_c, reg_f, reg_ff : in std_logic_vector (31 downto 0);  addr_c, 
            addr_f, addr_ff : in std_logic_vector (4 downto 0);  valid_f, 
            valid_ff, dirty_f, dirty_ff, en : in std_logic;  output : out 
            std_logic_vector (31 downto 0);  match_dirty_f, match_dirty_ff : 
            out std_logic);
   end component;
   
   component FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_0
      port( reg_c, reg_f, reg_ff : in std_logic_vector (31 downto 0);  addr_c, 
            addr_f, addr_ff : in std_logic_vector (4 downto 0);  valid_f, 
            valid_ff, dirty_f, dirty_ff, en : in std_logic;  output : out 
            std_logic_vector (31 downto 0);  match_dirty_f, match_dirty_ff : 
            out std_logic);
   end component;
   
   component Mux_DATA_SIZE32_6
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0)
            ;  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Adder_DATA_SIZE32_7
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;
   
   component Mux_DATA_SIZE32_7
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0)
            ;  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component RegisterFile_DATA_SIZE32_REG_NUM32
      port( clk, rst, en, rd1_en, rd2_en, wr_en, link_en : in std_logic;  
            rd1_addr, rd2_addr, wr_addr : in std_logic_vector (4 downto 0);  
            d_out1, d_out2 : out std_logic_vector (31 downto 0);  d_in, d_link 
            : in std_logic_vector (31 downto 0));
   end component;
   
   component Extender_SRC_SIZE26_DEST_SIZE32
      port( s : in std_logic;  i : in std_logic_vector (25 downto 0);  o : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component Extender_SRC_SIZE16_DEST_SIZE32
      port( s : in std_logic;  i : in std_logic_vector (15 downto 0);  o : out 
            std_logic_vector (31 downto 0));
   end component;
   
   component Mux_DATA_SIZE5
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (4 downto 0);
            dout : out std_logic_vector (4 downto 0));
   end component;
   
   component Mux_DATA_SIZE32_8
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0)
            ;  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Mux_DATA_SIZE32_9
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0)
            ;  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Reg_DATA_SIZE32_12
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 
            0);  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Reg_DATA_SIZE32_0
      port( rst, en, clk : in std_logic;  din : in std_logic_vector (31 downto 
            0);  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Mux_DATA_SIZE32_0
      port( sel : in std_logic;  din0, din1 : in std_logic_vector (31 downto 0)
            ;  dout : out std_logic_vector (31 downto 0));
   end component;
   
   component Adder_DATA_SIZE32_0
      port( cin : in std_logic;  a, b : in std_logic_vector (31 downto 0);  s :
            out std_logic_vector (31 downto 0);  cout : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, istr_addr_31_port, istr_addr_30_port, 
      istr_addr_29_port, istr_addr_28_port, istr_addr_27_port, 
      istr_addr_26_port, istr_addr_25_port, istr_addr_24_port, 
      istr_addr_23_port, istr_addr_22_port, istr_addr_21_port, 
      istr_addr_20_port, istr_addr_19_port, istr_addr_18_port, 
      istr_addr_17_port, istr_addr_16_port, istr_addr_15_port, 
      istr_addr_14_port, istr_addr_13_port, istr_addr_12_port, 
      istr_addr_11_port, istr_addr_10_port, istr_addr_9_port, istr_addr_8_port,
      istr_addr_7_port, istr_addr_6_port, istr_addr_5_port, istr_addr_4_port, 
      istr_addr_3_port, istr_addr_2_port, istr_addr_1_port, istr_addr_0_port, 
      data_addr_31_port, data_addr_30_port, data_addr_29_port, 
      data_addr_28_port, data_addr_27_port, data_addr_26_port, 
      data_addr_25_port, data_addr_24_port, data_addr_23_port, 
      data_addr_22_port, data_addr_21_port, data_addr_20_port, 
      data_addr_19_port, data_addr_18_port, data_addr_17_port, 
      data_addr_16_port, data_addr_15_port, data_addr_14_port, 
      data_addr_13_port, data_addr_12_port, data_addr_11_port, 
      data_addr_10_port, data_addr_9_port, data_addr_8_port, data_addr_7_port, 
      data_addr_6_port, data_addr_5_port, data_addr_4_port, data_addr_3_port, 
      data_addr_2_port, data_addr_1_port, data_addr_0_port, sig_ral_port, 
      sig_mul_port, sig_sqrt_port, s1_npc_31_port, s1_npc_30_port, 
      s1_npc_29_port, s1_npc_28_port, s1_npc_27_port, s1_npc_26_port, 
      s1_npc_25_port, s1_npc_24_port, s1_npc_23_port, s1_npc_22_port, 
      s1_npc_21_port, s1_npc_20_port, s1_npc_19_port, s1_npc_18_port, 
      s1_npc_17_port, s1_npc_16_port, s1_npc_15_port, s1_npc_14_port, 
      s1_npc_13_port, s1_npc_12_port, s1_npc_11_port, s1_npc_10_port, 
      s1_npc_9_port, s1_npc_8_port, s1_npc_7_port, s1_npc_6_port, s1_npc_5_port
      , s1_npc_4_port, s1_npc_3_port, s1_npc_2_port, s1_npc_1_port, 
      s1_npc_0_port, s2_pc_sel_31_port, s2_pc_sel_30_port, s2_pc_sel_29_port, 
      s2_pc_sel_28_port, s2_pc_sel_27_port, s2_pc_sel_26_port, 
      s2_pc_sel_25_port, s2_pc_sel_24_port, s2_pc_sel_23_port, 
      s2_pc_sel_22_port, s2_pc_sel_21_port, s2_pc_sel_20_port, 
      s2_pc_sel_19_port, s2_pc_sel_18_port, s2_pc_sel_17_port, 
      s2_pc_sel_16_port, s2_pc_sel_15_port, s2_pc_sel_14_port, 
      s2_pc_sel_13_port, s2_pc_sel_12_port, s2_pc_sel_11_port, 
      s2_pc_sel_10_port, s2_pc_sel_9_port, s2_pc_sel_8_port, s2_pc_sel_7_port, 
      s2_pc_sel_6_port, s2_pc_sel_5_port, s2_pc_sel_4_port, s2_pc_sel_3_port, 
      s2_pc_sel_2_port, s2_pc_sel_1_port, s2_pc_sel_0_port, 
      s3_pc_notsel_31_port, s3_pc_notsel_30_port, s3_pc_notsel_29_port, 
      s3_pc_notsel_28_port, s3_pc_notsel_27_port, s3_pc_notsel_26_port, 
      s3_pc_notsel_25_port, s3_pc_notsel_24_port, s3_pc_notsel_23_port, 
      s3_pc_notsel_22_port, s3_pc_notsel_21_port, s3_pc_notsel_20_port, 
      s3_pc_notsel_19_port, s3_pc_notsel_18_port, s3_pc_notsel_17_port, 
      s3_pc_notsel_16_port, s3_pc_notsel_15_port, s3_pc_notsel_14_port, 
      s3_pc_notsel_13_port, s3_pc_notsel_12_port, s3_pc_notsel_11_port, 
      s3_pc_notsel_10_port, s3_pc_notsel_9_port, s3_pc_notsel_8_port, 
      s3_pc_notsel_7_port, s3_pc_notsel_6_port, s3_pc_notsel_5_port, 
      s3_pc_notsel_4_port, s3_pc_notsel_3_port, s3_pc_notsel_2_port, 
      s3_pc_notsel_1_port, s3_pc_notsel_0_port, s2_npc_31_port, s2_npc_30_port,
      s2_npc_29_port, s2_npc_28_port, s2_npc_27_port, s2_npc_26_port, 
      s2_npc_25_port, s2_npc_24_port, s2_npc_23_port, s2_npc_22_port, 
      s2_npc_21_port, s2_npc_20_port, s2_npc_19_port, s2_npc_18_port, 
      s2_npc_17_port, s2_npc_16_port, s2_npc_15_port, s2_npc_14_port, 
      s2_npc_13_port, s2_npc_12_port, s2_npc_11_port, s2_npc_10_port, 
      s2_npc_9_port, s2_npc_8_port, s2_npc_7_port, s2_npc_6_port, s2_npc_5_port
      , s2_npc_4_port, s2_npc_3_port, s2_npc_2_port, s2_npc_1_port, 
      s2_npc_0_port, s2_jpc_30_port, s2_jpc_29_port, s2_jpc_28_port, 
      s2_jpc_27_port, s2_jpc_26_port, s2_jpc_25_port, s2_jpc_24_port, 
      s2_jpc_23_port, s2_jpc_22_port, s2_jpc_21_port, s2_jpc_20_port, 
      s2_jpc_19_port, s2_jpc_18_port, s2_jpc_17_port, s2_jpc_16_port, 
      s2_jpc_15_port, s2_jpc_14_port, s2_jpc_13_port, s2_jpc_12_port, 
      s2_jpc_11_port, s2_jpc_10_port, s2_jpc_9_port, s2_jpc_8_port, 
      s2_jpc_7_port, s2_jpc_6_port, s2_jpc_5_port, s2_jpc_4_port, s2_jpc_3_port
      , s2_jpc_2_port, s2_jpc_1_port, s2_jpc_0_port, s2_pc_notsel_31_port, 
      s2_pc_notsel_30_port, s2_pc_notsel_29_port, s2_pc_notsel_28_port, 
      s2_pc_notsel_27_port, s2_pc_notsel_26_port, s2_pc_notsel_25_port, 
      s2_pc_notsel_24_port, s2_pc_notsel_23_port, s2_pc_notsel_22_port, 
      s2_pc_notsel_21_port, s2_pc_notsel_20_port, s2_pc_notsel_19_port, 
      s2_pc_notsel_18_port, s2_pc_notsel_17_port, s2_pc_notsel_16_port, 
      s2_pc_notsel_15_port, s2_pc_notsel_14_port, s2_pc_notsel_13_port, 
      s2_pc_notsel_12_port, s2_pc_notsel_11_port, s2_pc_notsel_10_port, 
      s2_pc_notsel_9_port, s2_pc_notsel_8_port, s2_pc_notsel_7_port, 
      s2_pc_notsel_6_port, s2_pc_notsel_5_port, s2_pc_notsel_4_port, 
      s2_pc_notsel_3_port, s2_pc_notsel_2_port, s2_pc_notsel_1_port, 
      s2_pc_notsel_0_port, s2_wr_addr_sel, s2_wr_addr_4_port, s2_wr_addr_3_port
      , s2_wr_addr_2_port, s2_wr_addr_1_port, s2_wr_addr_0_port, 
      s2_imm_l_ext_31_port, s2_imm_l_ext_15_port, s2_imm_l_ext_14_port, 
      s2_imm_l_ext_13_port, s2_imm_l_ext_12_port, s2_imm_l_ext_11_port, 
      s2_imm_l_ext_10_port, s2_imm_l_ext_9_port, s2_imm_l_ext_8_port, 
      s2_imm_l_ext_7_port, s2_imm_l_ext_6_port, s2_imm_l_ext_5_port, 
      s2_imm_l_ext_4_port, s2_imm_l_ext_3_port, s2_imm_l_ext_2_port, 
      s2_imm_l_ext_1_port, s2_imm_l_ext_0_port, s2_imm_j_ext_31_port, 
      s2_imm_j_ext_30_port, s2_imm_j_ext_29_port, s2_imm_j_ext_28_port, 
      s2_imm_j_ext_27_port, s2_imm_j_ext_26_port, s2_imm_j_ext_25_port, 
      s2_imm_j_ext_24_port, s2_imm_j_ext_23_port, s2_imm_j_ext_22_port, 
      s2_imm_j_ext_21_port, s2_imm_j_ext_20_port, s2_imm_j_ext_19_port, 
      s2_imm_j_ext_18_port, s2_imm_j_ext_17_port, s2_imm_j_ext_16_port, 
      s2_imm_j_ext_15_port, s2_imm_j_ext_14_port, s2_imm_j_ext_13_port, 
      s2_imm_j_ext_12_port, s2_imm_j_ext_11_port, s2_imm_j_ext_10_port, 
      s2_imm_j_ext_9_port, s2_imm_j_ext_8_port, s2_imm_j_ext_7_port, 
      s2_imm_j_ext_6_port, s2_imm_j_ext_5_port, s2_imm_j_ext_4_port, 
      s2_imm_j_ext_3_port, s2_imm_j_ext_2_port, s2_imm_j_ext_1_port, 
      s2_imm_j_ext_0_port, s2_imm_i_ext_31_port, s2_imm_i_ext_30_port, 
      s2_imm_i_ext_29_port, s2_imm_i_ext_28_port, s2_imm_i_ext_27_port, 
      s2_imm_i_ext_26_port, s2_imm_i_ext_25_port, s2_imm_i_ext_24_port, 
      s2_imm_i_ext_23_port, s2_imm_i_ext_22_port, s2_imm_i_ext_21_port, 
      s2_imm_i_ext_20_port, s2_imm_i_ext_19_port, s2_imm_i_ext_18_port, 
      s2_imm_i_ext_17_port, s2_imm_i_ext_16_port, s2_imm_i_ext_15_port, 
      s2_imm_i_ext_14_port, s2_imm_i_ext_13_port, s2_imm_i_ext_12_port, 
      s2_imm_i_ext_11_port, s2_imm_i_ext_10_port, s2_imm_i_ext_9_port, 
      s2_imm_i_ext_8_port, s2_imm_i_ext_7_port, s2_imm_i_ext_6_port, 
      s2_imm_i_ext_5_port, s2_imm_i_ext_4_port, s2_imm_i_ext_3_port, 
      s2_imm_i_ext_2_port, s2_imm_i_ext_1_port, s2_imm_i_ext_0_port, s2_rf_en, 
      s5_wr_addr_4_port, s5_wr_addr_3_port, s5_wr_addr_2_port, 
      s5_wr_addr_1_port, s5_wr_addr_0_port, s2_a_31_port, s2_a_30_port, 
      s2_a_29_port, s2_a_28_port, s2_a_27_port, s2_a_26_port, s2_a_25_port, 
      s2_a_24_port, s2_a_23_port, s2_a_22_port, s2_a_21_port, s2_a_20_port, 
      s2_a_19_port, s2_a_18_port, s2_a_17_port, s2_a_16_port, s2_a_15_port, 
      s2_a_14_port, s2_a_13_port, s2_a_12_port, s2_a_11_port, s2_a_10_port, 
      s2_a_9_port, s2_a_8_port, s2_a_7_port, s2_a_6_port, s2_a_5_port, 
      s2_a_4_port, s2_a_3_port, s2_a_2_port, s2_a_1_port, s2_a_0_port, 
      s2_b_31_port, s2_b_30_port, s2_b_29_port, s2_b_28_port, s2_b_27_port, 
      s2_b_26_port, s2_b_25_port, s2_b_24_port, s2_b_23_port, s2_b_22_port, 
      s2_b_21_port, s2_b_20_port, s2_b_19_port, s2_b_18_port, s2_b_17_port, 
      s2_b_16_port, s2_b_15_port, s2_b_14_port, s2_b_13_port, s2_b_12_port, 
      s2_b_11_port, s2_b_10_port, s2_b_9_port, s2_b_8_port, s2_b_7_port, 
      s2_b_6_port, s2_b_5_port, s2_b_4_port, s2_b_3_port, s2_b_2_port, 
      s2_b_1_port, s2_b_0_port, s5_result_31_port, s5_result_30_port, 
      s5_result_29_port, s5_result_28_port, s5_result_27_port, 
      s5_result_26_port, s5_result_25_port, s5_result_24_port, 
      s5_result_23_port, s5_result_22_port, s5_result_21_port, 
      s5_result_20_port, s5_result_19_port, s5_result_18_port, 
      s5_result_17_port, s5_result_16_port, s5_result_15_port, 
      s5_result_14_port, s5_result_13_port, s5_result_12_port, 
      s5_result_11_port, s5_result_10_port, s5_result_9_port, s5_result_8_port,
      s5_result_7_port, s5_result_6_port, s5_result_5_port, s5_result_4_port, 
      s5_result_3_port, s5_result_2_port, s5_result_1_port, s5_result_0_port, 
      s2_jump_addr_imm_31_port, s2_jump_addr_imm_30_port, 
      s2_jump_addr_imm_29_port, s2_jump_addr_imm_28_port, 
      s2_jump_addr_imm_27_port, s2_jump_addr_imm_26_port, 
      s2_jump_addr_imm_25_port, s2_jump_addr_imm_24_port, 
      s2_jump_addr_imm_23_port, s2_jump_addr_imm_22_port, 
      s2_jump_addr_imm_21_port, s2_jump_addr_imm_20_port, 
      s2_jump_addr_imm_19_port, s2_jump_addr_imm_18_port, 
      s2_jump_addr_imm_17_port, s2_jump_addr_imm_16_port, 
      s2_jump_addr_imm_15_port, s2_jump_addr_imm_14_port, 
      s2_jump_addr_imm_13_port, s2_jump_addr_imm_12_port, 
      s2_jump_addr_imm_11_port, s2_jump_addr_imm_10_port, 
      s2_jump_addr_imm_9_port, s2_jump_addr_imm_8_port, s2_jump_addr_imm_7_port
      , s2_jump_addr_imm_6_port, s2_jump_addr_imm_5_port, 
      s2_jump_addr_imm_4_port, s2_jump_addr_imm_3_port, s2_jump_addr_imm_2_port
      , s2_jump_addr_imm_1_port, s2_jump_addr_imm_0_port, 
      s2_jump_addr_rel_31_port, s2_jump_addr_rel_30_port, 
      s2_jump_addr_rel_29_port, s2_jump_addr_rel_28_port, 
      s2_jump_addr_rel_27_port, s2_jump_addr_rel_26_port, 
      s2_jump_addr_rel_25_port, s2_jump_addr_rel_24_port, 
      s2_jump_addr_rel_23_port, s2_jump_addr_rel_22_port, 
      s2_jump_addr_rel_21_port, s2_jump_addr_rel_20_port, 
      s2_jump_addr_rel_19_port, s2_jump_addr_rel_18_port, 
      s2_jump_addr_rel_17_port, s2_jump_addr_rel_16_port, 
      s2_jump_addr_rel_15_port, s2_jump_addr_rel_14_port, 
      s2_jump_addr_rel_13_port, s2_jump_addr_rel_12_port, 
      s2_jump_addr_rel_11_port, s2_jump_addr_rel_10_port, 
      s2_jump_addr_rel_9_port, s2_jump_addr_rel_8_port, s2_jump_addr_rel_7_port
      , s2_jump_addr_rel_6_port, s2_jump_addr_rel_5_port, 
      s2_jump_addr_rel_4_port, s2_jump_addr_rel_3_port, s2_jump_addr_rel_2_port
      , s2_jump_addr_rel_1_port, s2_jump_addr_rel_0_port, 
      s2_jump_addr_reg_31_port, s2_jump_addr_reg_30_port, 
      s2_jump_addr_reg_29_port, s2_jump_addr_reg_28_port, 
      s2_jump_addr_reg_27_port, s2_jump_addr_reg_26_port, 
      s2_jump_addr_reg_25_port, s2_jump_addr_reg_24_port, 
      s2_jump_addr_reg_23_port, s2_jump_addr_reg_22_port, 
      s2_jump_addr_reg_21_port, s2_jump_addr_reg_20_port, 
      s2_jump_addr_reg_19_port, s2_jump_addr_reg_18_port, 
      s2_jump_addr_reg_17_port, s2_jump_addr_reg_16_port, 
      s2_jump_addr_reg_15_port, s2_jump_addr_reg_14_port, 
      s2_jump_addr_reg_13_port, s2_jump_addr_reg_12_port, 
      s2_jump_addr_reg_11_port, s2_jump_addr_reg_10_port, 
      s2_jump_addr_reg_9_port, s2_jump_addr_reg_8_port, s2_jump_addr_reg_7_port
      , s2_jump_addr_reg_6_port, s2_jump_addr_reg_5_port, 
      s2_jump_addr_reg_4_port, s2_jump_addr_reg_3_port, s2_jump_addr_reg_2_port
      , s2_jump_addr_reg_1_port, s2_jump_addr_reg_0_port, s2_a_f_b_en, 
      s2_a_ff_b_en, s3_exe_out_31_port, s3_exe_out_30_port, s3_exe_out_29_port,
      s3_exe_out_28_port, s3_exe_out_27_port, s3_exe_out_26_port, 
      s3_exe_out_25_port, s3_exe_out_24_port, s3_exe_out_23_port, 
      s3_exe_out_22_port, s3_exe_out_21_port, s3_exe_out_20_port, 
      s3_exe_out_19_port, s3_exe_out_18_port, s3_exe_out_17_port, 
      s3_exe_out_16_port, s3_exe_out_15_port, s3_exe_out_14_port, 
      s3_exe_out_13_port, s3_exe_out_12_port, s3_exe_out_11_port, 
      s3_exe_out_10_port, s3_exe_out_9_port, s3_exe_out_8_port, 
      s3_exe_out_7_port, s3_exe_out_6_port, s3_exe_out_5_port, 
      s3_exe_out_4_port, s3_exe_out_3_port, s3_exe_out_2_port, 
      s3_exe_out_1_port, s3_exe_out_0_port, s4_result_31_port, 
      s4_result_30_port, s4_result_29_port, s4_result_28_port, 
      s4_result_27_port, s4_result_26_port, s4_result_25_port, 
      s4_result_24_port, s4_result_23_port, s4_result_22_port, 
      s4_result_21_port, s4_result_20_port, s4_result_19_port, 
      s4_result_18_port, s4_result_17_port, s4_result_16_port, 
      s4_result_15_port, s4_result_14_port, s4_result_13_port, 
      s4_result_12_port, s4_result_11_port, s4_result_10_port, s4_result_9_port
      , s4_result_8_port, s4_result_7_port, s4_result_6_port, s4_result_5_port,
      s4_result_4_port, s4_result_3_port, s4_result_2_port, s4_result_1_port, 
      s4_result_0_port, s3_wr_addr_4_port, s3_wr_addr_3_port, s3_wr_addr_2_port
      , s3_wr_addr_1_port, s3_wr_addr_0_port, s4_wr_addr_4_port, 
      s4_wr_addr_3_port, s4_wr_addr_2_port, s4_wr_addr_1_port, 
      s4_wr_addr_0_port, s2_a_f_j_en, s2_a_ff_j_en, s3_a_31_port, s3_a_30_port,
      s3_a_29_port, s3_a_28_port, s3_a_27_port, s3_a_26_port, s3_a_25_port, 
      s3_a_24_port, s3_a_23_port, s3_a_22_port, s3_a_21_port, s3_a_20_port, 
      s3_a_19_port, s3_a_18_port, s3_a_17_port, s3_a_16_port, s3_a_15_port, 
      s3_a_14_port, s3_a_13_port, s3_a_12_port, s3_a_11_port, s3_a_10_port, 
      s3_a_9_port, s3_a_8_port, s3_a_7_port, s3_a_6_port, s3_a_5_port, 
      s3_a_4_port, s3_a_3_port, s3_a_2_port, s3_a_1_port, s3_a_0_port, 
      s3_b_31_port, s3_b_30_port, s3_b_29_port, s3_b_28_port, s3_b_27_port, 
      s3_b_26_port, s3_b_25_port, s3_b_24_port, s3_b_23_port, s3_b_22_port, 
      s3_b_21_port, s3_b_20_port, s3_b_19_port, s3_b_18_port, s3_b_17_port, 
      s3_b_16_port, s3_b_15_port, s3_b_14_port, s3_b_13_port, s3_b_12_port, 
      s3_b_11_port, s3_b_10_port, s3_b_9_port, s3_b_8_port, s3_b_7_port, 
      s3_b_6_port, s3_b_5_port, s3_b_4_port, s3_b_3_port, s3_b_2_port, 
      s3_b_1_port, s3_b_0_port, s3_imm_i_ext_31_port, s3_imm_i_ext_30_port, 
      s3_imm_i_ext_29_port, s3_imm_i_ext_28_port, s3_imm_i_ext_27_port, 
      s3_imm_i_ext_26_port, s3_imm_i_ext_25_port, s3_imm_i_ext_24_port, 
      s3_imm_i_ext_23_port, s3_imm_i_ext_22_port, s3_imm_i_ext_21_port, 
      s3_imm_i_ext_20_port, s3_imm_i_ext_19_port, s3_imm_i_ext_18_port, 
      s3_imm_i_ext_17_port, s3_imm_i_ext_16_port, s3_imm_i_ext_15_port, 
      s3_imm_i_ext_14_port, s3_imm_i_ext_13_port, s3_imm_i_ext_12_port, 
      s3_imm_i_ext_11_port, s3_imm_i_ext_10_port, s3_imm_i_ext_9_port, 
      s3_imm_i_ext_8_port, s3_imm_i_ext_7_port, s3_imm_i_ext_6_port, 
      s3_imm_i_ext_5_port, s3_imm_i_ext_4_port, s3_imm_i_ext_3_port, 
      s3_imm_i_ext_2_port, s3_imm_i_ext_1_port, s3_imm_i_ext_0_port, 
      s3_rd1_addr_4_port, s3_rd1_addr_3_port, s3_rd1_addr_2_port, 
      s3_rd1_addr_1_port, s3_rd1_addr_0_port, s3_rd2_addr_4_port, 
      s3_rd2_addr_3_port, s3_rd2_addr_2_port, s3_rd2_addr_1_port, 
      s3_rd2_addr_0_port, s3_jump_flag, s4_reg_b_wait, s4_a_31_port, 
      s4_a_30_port, s4_a_29_port, s4_a_28_port, s4_a_27_port, s4_a_26_port, 
      s4_a_25_port, s4_a_24_port, s4_a_23_port, s4_a_22_port, s4_a_21_port, 
      s4_a_20_port, s4_a_19_port, s4_a_18_port, s4_a_17_port, s4_a_16_port, 
      s4_a_15_port, s4_a_14_port, s4_a_13_port, s4_a_12_port, s4_a_11_port, 
      s4_a_10_port, s4_a_9_port, s4_a_8_port, s4_a_7_port, s4_a_6_port, 
      s4_a_5_port, s4_a_4_port, s4_a_3_port, s4_a_2_port, s4_a_1_port, 
      s4_a_0_port, s3_a_keep_31_port, s3_a_keep_30_port, s3_a_keep_29_port, 
      s3_a_keep_28_port, s3_a_keep_27_port, s3_a_keep_26_port, 
      s3_a_keep_25_port, s3_a_keep_24_port, s3_a_keep_23_port, 
      s3_a_keep_22_port, s3_a_keep_21_port, s3_a_keep_20_port, 
      s3_a_keep_19_port, s3_a_keep_18_port, s3_a_keep_17_port, 
      s3_a_keep_16_port, s3_a_keep_15_port, s3_a_keep_14_port, 
      s3_a_keep_13_port, s3_a_keep_12_port, s3_a_keep_11_port, 
      s3_a_keep_10_port, s3_a_keep_9_port, s3_a_keep_8_port, s3_a_keep_7_port, 
      s3_a_keep_6_port, s3_a_keep_5_port, s3_a_keep_4_port, s3_a_keep_3_port, 
      s3_a_keep_2_port, s3_a_keep_1_port, s3_a_keep_0_port, s4_reg_a_wait, 
      s4_b_31_port, s4_b_30_port, s4_b_29_port, s4_b_28_port, s4_b_27_port, 
      s4_b_26_port, s4_b_25_port, s4_b_24_port, s4_b_23_port, s4_b_22_port, 
      s4_b_21_port, s4_b_20_port, s4_b_19_port, s4_b_18_port, s4_b_17_port, 
      s4_b_16_port, s4_b_15_port, s4_b_14_port, s4_b_13_port, s4_b_12_port, 
      s4_b_11_port, s4_b_10_port, s4_b_9_port, s4_b_8_port, s4_b_7_port, 
      s4_b_6_port, s4_b_5_port, s4_b_4_port, s4_b_3_port, s4_b_2_port, 
      s4_b_1_port, s4_b_0_port, s3_b_keep_31_port, s3_b_keep_30_port, 
      s3_b_keep_29_port, s3_b_keep_28_port, s3_b_keep_27_port, 
      s3_b_keep_26_port, s3_b_keep_25_port, s3_b_keep_24_port, 
      s3_b_keep_23_port, s3_b_keep_22_port, s3_b_keep_21_port, 
      s3_b_keep_20_port, s3_b_keep_19_port, s3_b_keep_18_port, 
      s3_b_keep_17_port, s3_b_keep_16_port, s3_b_keep_15_port, 
      s3_b_keep_14_port, s3_b_keep_13_port, s3_b_keep_12_port, 
      s3_b_keep_11_port, s3_b_keep_10_port, s3_b_keep_9_port, s3_b_keep_8_port,
      s3_b_keep_7_port, s3_b_keep_6_port, s3_b_keep_5_port, s3_b_keep_4_port, 
      s3_b_keep_3_port, s3_b_keep_2_port, s3_b_keep_1_port, s3_b_keep_0_port, 
      s3_a_sel_f_en, s3_a_sel_ff_en, s3_a_sel_31_port, s3_a_sel_30_port, 
      s3_a_sel_29_port, s3_a_sel_28_port, s3_a_sel_27_port, s3_a_sel_26_port, 
      s3_a_sel_25_port, s3_a_sel_24_port, s3_a_sel_23_port, s3_a_sel_22_port, 
      s3_a_sel_21_port, s3_a_sel_20_port, s3_a_sel_19_port, s3_a_sel_18_port, 
      s3_a_sel_17_port, s3_a_sel_16_port, s3_a_sel_15_port, s3_a_sel_14_port, 
      s3_a_sel_13_port, s3_a_sel_12_port, s3_a_sel_11_port, s3_a_sel_10_port, 
      s3_a_sel_9_port, s3_a_sel_8_port, s3_a_sel_7_port, s3_a_sel_6_port, 
      s3_a_sel_5_port, s3_a_sel_4_port, s3_a_sel_3_port, s3_a_sel_2_port, 
      s3_a_sel_1_port, s3_a_sel_0_port, s3_reg_a_wait, s3_b_sel_f_en, 
      s3_b_sel_ff_en, s3_b_fwd_31_port, s3_b_fwd_30_port, s3_b_fwd_29_port, 
      s3_b_fwd_28_port, s3_b_fwd_27_port, s3_b_fwd_26_port, s3_b_fwd_25_port, 
      s3_b_fwd_24_port, s3_b_fwd_23_port, s3_b_fwd_22_port, s3_b_fwd_21_port, 
      s3_b_fwd_20_port, s3_b_fwd_19_port, s3_b_fwd_18_port, s3_b_fwd_17_port, 
      s3_b_fwd_16_port, s3_b_fwd_15_port, s3_b_fwd_14_port, s3_b_fwd_13_port, 
      s3_b_fwd_12_port, s3_b_fwd_11_port, s3_b_fwd_10_port, s3_b_fwd_9_port, 
      s3_b_fwd_8_port, s3_b_fwd_7_port, s3_b_fwd_6_port, s3_b_fwd_5_port, 
      s3_b_fwd_4_port, s3_b_fwd_3_port, s3_b_fwd_2_port, s3_b_fwd_1_port, 
      s3_b_fwd_0_port, s3_reg_b_wait, s3_b_sel_31_port, s3_b_sel_30_port, 
      s3_b_sel_29_port, s3_b_sel_28_port, s3_b_sel_27_port, s3_b_sel_26_port, 
      s3_b_sel_25_port, s3_b_sel_24_port, s3_b_sel_23_port, s3_b_sel_22_port, 
      s3_b_sel_21_port, s3_b_sel_20_port, s3_b_sel_19_port, s3_b_sel_18_port, 
      s3_b_sel_17_port, s3_b_sel_16_port, s3_b_sel_15_port, s3_b_sel_14_port, 
      s3_b_sel_13_port, s3_b_sel_12_port, s3_b_sel_11_port, s3_b_sel_10_port, 
      s3_b_sel_9_port, s3_b_sel_8_port, s3_b_sel_7_port, s3_b_sel_6_port, 
      s3_b_sel_5_port, s3_b_sel_4_port, s3_b_sel_3_port, s3_b_sel_2_port, 
      s3_b_sel_1_port, s3_b_sel_0_port, s3_alu_out_31_port, s3_alu_out_30_port,
      s3_alu_out_29_port, s3_alu_out_28_port, s3_alu_out_27_port, 
      s3_alu_out_26_port, s3_alu_out_25_port, s3_alu_out_24_port, 
      s3_alu_out_23_port, s3_alu_out_22_port, s3_alu_out_21_port, 
      s3_alu_out_20_port, s3_alu_out_19_port, s3_alu_out_18_port, 
      s3_alu_out_17_port, s3_alu_out_16_port, s3_alu_out_15_port, 
      s3_alu_out_14_port, s3_alu_out_13_port, s3_alu_out_12_port, 
      s3_alu_out_11_port, s3_alu_out_10_port, s3_alu_out_9_port, 
      s3_alu_out_8_port, s3_alu_out_7_port, s3_alu_out_6_port, 
      s3_alu_out_5_port, s3_alu_out_4_port, s3_alu_out_3_port, 
      s3_alu_out_2_port, s3_alu_out_1_port, s3_alu_out_0_port, s3_mul_sign, 
      s3_mul_out_31_port, s3_mul_out_30_port, s3_mul_out_29_port, 
      s3_mul_out_28_port, s3_mul_out_27_port, s3_mul_out_26_port, 
      s3_mul_out_25_port, s3_mul_out_24_port, s3_mul_out_23_port, 
      s3_mul_out_22_port, s3_mul_out_21_port, s3_mul_out_20_port, 
      s3_mul_out_19_port, s3_mul_out_18_port, s3_mul_out_17_port, 
      s3_mul_out_16_port, s3_mul_out_15_port, s3_mul_out_14_port, 
      s3_mul_out_13_port, s3_mul_out_12_port, s3_mul_out_11_port, 
      s3_mul_out_10_port, s3_mul_out_9_port, s3_mul_out_8_port, 
      s3_mul_out_7_port, s3_mul_out_6_port, s3_mul_out_5_port, 
      s3_mul_out_4_port, s3_mul_out_3_port, s3_mul_out_2_port, 
      s3_mul_out_1_port, s3_mul_out_0_port, s3_div_sign, s3_div_out_31_port, 
      s3_div_out_30_port, s3_div_out_29_port, s3_div_out_28_port, 
      s3_div_out_27_port, s3_div_out_26_port, s3_div_out_25_port, 
      s3_div_out_24_port, s3_div_out_23_port, s3_div_out_22_port, 
      s3_div_out_21_port, s3_div_out_20_port, s3_div_out_19_port, 
      s3_div_out_18_port, s3_div_out_17_port, s3_div_out_16_port, 
      s3_div_out_15_port, s3_div_out_14_port, s3_div_out_13_port, 
      s3_div_out_12_port, s3_div_out_11_port, s3_div_out_10_port, 
      s3_div_out_9_port, s3_div_out_8_port, s3_div_out_7_port, 
      s3_div_out_6_port, s3_div_out_5_port, s3_div_out_4_port, 
      s3_div_out_3_port, s3_div_out_2_port, s3_div_out_1_port, 
      s3_div_out_0_port, s3_exe_sel_1_port, s4_b_fwd_31_port, s4_b_fwd_30_port,
      s4_b_fwd_29_port, s4_b_fwd_28_port, s4_b_fwd_27_port, s4_b_fwd_26_port, 
      s4_b_fwd_25_port, s4_b_fwd_24_port, s4_b_fwd_23_port, s4_b_fwd_22_port, 
      s4_b_fwd_21_port, s4_b_fwd_20_port, s4_b_fwd_19_port, s4_b_fwd_18_port, 
      s4_b_fwd_17_port, s4_b_fwd_16_port, s4_b_fwd_15_port, s4_b_fwd_14_port, 
      s4_b_fwd_13_port, s4_b_fwd_12_port, s4_b_fwd_11_port, s4_b_fwd_10_port, 
      s4_b_fwd_9_port, s4_b_fwd_8_port, s4_b_fwd_7_port, s4_b_fwd_6_port, 
      s4_b_fwd_5_port, s4_b_fwd_4_port, s4_b_fwd_3_port, s4_b_fwd_2_port, 
      s4_b_fwd_1_port, s4_b_fwd_0_port, s4_rd2_addr_4_port, s4_rd2_addr_3_port,
      s4_rd2_addr_2_port, s4_rd2_addr_1_port, s4_rd2_addr_0_port, 
      s6_result_31_port, s6_result_30_port, s6_result_29_port, 
      s6_result_28_port, s6_result_27_port, s6_result_26_port, 
      s6_result_25_port, s6_result_24_port, s6_result_23_port, 
      s6_result_22_port, s6_result_21_port, s6_result_20_port, 
      s6_result_19_port, s6_result_18_port, s6_result_17_port, 
      s6_result_16_port, s6_result_15_port, s6_result_14_port, 
      s6_result_13_port, s6_result_12_port, s6_result_11_port, 
      s6_result_10_port, s6_result_9_port, s6_result_8_port, s6_result_7_port, 
      s6_result_6_port, s6_result_5_port, s6_result_4_port, s6_result_3_port, 
      s6_result_2_port, s6_result_1_port, s6_result_0_port, s6_wr_addr_4_port, 
      s6_wr_addr_3_port, s6_wr_addr_2_port, s6_wr_addr_1_port, 
      s6_wr_addr_0_port, s6_en_wb, net1283, net1284, net1287, net1288, net1290,
      net1291, net1292, net1293, net1294, n44, n45, n48, n1, n2, n3, n4, n5, n6
      , n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
      n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36
      , n37, n38, n39, n40, n41, n42, n43, n46, net107975, net107976, net107977
      , net107978, net107979, net107980, net107981, net107982, net107983, 
      net107984, net107985, net107986, net107987, net107988, net107989, 
      net107990 : std_logic;

begin
   istr_addr <= ( istr_addr_31_port, istr_addr_30_port, istr_addr_29_port, 
      istr_addr_28_port, istr_addr_27_port, istr_addr_26_port, 
      istr_addr_25_port, istr_addr_24_port, istr_addr_23_port, 
      istr_addr_22_port, istr_addr_21_port, istr_addr_20_port, 
      istr_addr_19_port, istr_addr_18_port, istr_addr_17_port, 
      istr_addr_16_port, istr_addr_15_port, istr_addr_14_port, 
      istr_addr_13_port, istr_addr_12_port, istr_addr_11_port, 
      istr_addr_10_port, istr_addr_9_port, istr_addr_8_port, istr_addr_7_port, 
      istr_addr_6_port, istr_addr_5_port, istr_addr_4_port, istr_addr_3_port, 
      istr_addr_2_port, istr_addr_1_port, istr_addr_0_port );
   ir_out <= ( istr_val(31), istr_val(30), istr_val(29), istr_val(28), 
      istr_val(27), istr_val(26), istr_val(25), istr_val(24), istr_val(23), 
      istr_val(22), istr_val(21), istr_val(20), istr_val(19), istr_val(18), 
      istr_val(17), istr_val(16), istr_val(15), istr_val(14), istr_val(13), 
      istr_val(12), istr_val(11), istr_val(10), istr_val(9), istr_val(8), 
      istr_val(7), istr_val(6), istr_val(5), istr_val(4), istr_val(3), 
      istr_val(2), istr_val(1), istr_val(0) );
   ld_a_out <= ( data_i_val(31), data_i_val(30), data_i_val(29), data_i_val(28)
      , data_i_val(27), data_i_val(26), data_i_val(25), data_i_val(24), 
      data_i_val(23), data_i_val(22), data_i_val(21), data_i_val(20), 
      data_i_val(19), data_i_val(18), data_i_val(17), data_i_val(16), 
      data_i_val(15), data_i_val(14), data_i_val(13), data_i_val(12), 
      data_i_val(11), data_i_val(10), data_i_val(9), data_i_val(8), 
      data_i_val(7), data_i_val(6), data_i_val(5), data_i_val(4), data_i_val(3)
      , data_i_val(2), data_i_val(1), data_i_val(0) );
   data_addr <= ( data_addr_31_port, data_addr_30_port, data_addr_29_port, 
      data_addr_28_port, data_addr_27_port, data_addr_26_port, 
      data_addr_25_port, data_addr_24_port, data_addr_23_port, 
      data_addr_22_port, data_addr_21_port, data_addr_20_port, 
      data_addr_19_port, data_addr_18_port, data_addr_17_port, 
      data_addr_16_port, data_addr_15_port, data_addr_14_port, 
      data_addr_13_port, data_addr_12_port, data_addr_11_port, 
      data_addr_10_port, data_addr_9_port, data_addr_8_port, data_addr_7_port, 
      data_addr_6_port, data_addr_5_port, data_addr_4_port, data_addr_3_port, 
      data_addr_2_port, data_addr_1_port, data_addr_0_port );
   dr_cw <= ( cw(14), cw(13), cw(12), cw(11) );
   sig_ral <= sig_ral_port;
   sig_mul <= sig_mul_port;
   sig_sqrt <= sig_sqrt_port;
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   s3_jump_flag_reg : DFF_X1 port map( D => n48, CK => clk, Q => s3_jump_flag, 
                           QN => net107990);
   s6_en_wb_reg : DFFR_X1 port map( D => n45, CK => clk, RN => rst, Q => 
                           s6_en_wb, QN => n44);
   ADD_4 : Adder_DATA_SIZE32_0 port map( cin => X_Logic0_port, a(31) => 
                           istr_addr_31_port, a(30) => istr_addr_30_port, a(29)
                           => istr_addr_29_port, a(28) => istr_addr_28_port, 
                           a(27) => istr_addr_27_port, a(26) => 
                           istr_addr_26_port, a(25) => istr_addr_25_port, a(24)
                           => istr_addr_24_port, a(23) => istr_addr_23_port, 
                           a(22) => istr_addr_22_port, a(21) => 
                           istr_addr_21_port, a(20) => istr_addr_20_port, a(19)
                           => istr_addr_19_port, a(18) => istr_addr_18_port, 
                           a(17) => istr_addr_17_port, a(16) => 
                           istr_addr_16_port, a(15) => istr_addr_15_port, a(14)
                           => istr_addr_14_port, a(13) => istr_addr_13_port, 
                           a(12) => istr_addr_12_port, a(11) => 
                           istr_addr_11_port, a(10) => istr_addr_10_port, a(9) 
                           => istr_addr_9_port, a(8) => istr_addr_8_port, a(7) 
                           => istr_addr_7_port, a(6) => istr_addr_6_port, a(5) 
                           => istr_addr_5_port, a(4) => istr_addr_4_port, a(3) 
                           => istr_addr_3_port, a(2) => istr_addr_2_port, a(1) 
                           => istr_addr_1_port, a(0) => istr_addr_0_port, b(31)
                           => X_Logic0_port, b(30) => X_Logic0_port, b(29) => 
                           X_Logic0_port, b(28) => X_Logic0_port, b(27) => 
                           X_Logic0_port, b(26) => X_Logic0_port, b(25) => 
                           X_Logic0_port, b(24) => X_Logic0_port, b(23) => 
                           X_Logic0_port, b(22) => X_Logic0_port, b(21) => 
                           X_Logic0_port, b(20) => X_Logic0_port, b(19) => 
                           X_Logic0_port, b(18) => X_Logic0_port, b(17) => 
                           X_Logic0_port, b(16) => X_Logic0_port, b(15) => 
                           X_Logic0_port, b(14) => X_Logic0_port, b(13) => 
                           X_Logic0_port, b(12) => X_Logic0_port, b(11) => 
                           X_Logic0_port, b(10) => X_Logic0_port, b(9) => 
                           X_Logic0_port, b(8) => X_Logic0_port, b(7) => 
                           X_Logic0_port, b(6) => X_Logic0_port, b(5) => 
                           X_Logic0_port, b(4) => X_Logic0_port, b(3) => 
                           X_Logic0_port, b(2) => X_Logic0_port, b(1) => 
                           X_Logic0_port, b(0) => X_Logic0_port, s(31) => 
                           s1_npc_31_port, s(30) => s1_npc_30_port, s(29) => 
                           s1_npc_29_port, s(28) => s1_npc_28_port, s(27) => 
                           s1_npc_27_port, s(26) => s1_npc_26_port, s(25) => 
                           s1_npc_25_port, s(24) => s1_npc_24_port, s(23) => 
                           s1_npc_23_port, s(22) => s1_npc_22_port, s(21) => 
                           s1_npc_21_port, s(20) => s1_npc_20_port, s(19) => 
                           s1_npc_19_port, s(18) => s1_npc_18_port, s(17) => 
                           s1_npc_17_port, s(16) => s1_npc_16_port, s(15) => 
                           s1_npc_15_port, s(14) => s1_npc_14_port, s(13) => 
                           s1_npc_13_port, s(12) => s1_npc_12_port, s(11) => 
                           s1_npc_11_port, s(10) => s1_npc_10_port, s(9) => 
                           s1_npc_9_port, s(8) => s1_npc_8_port, s(7) => 
                           s1_npc_7_port, s(6) => s1_npc_6_port, s(5) => 
                           s1_npc_5_port, s(4) => s1_npc_4_port, s(3) => 
                           s1_npc_3_port, s(2) => s1_npc_2_port, s(1) => 
                           s1_npc_1_port, s(0) => s1_npc_0_port, cout => 
                           net1294);
   MUX_bpw : Mux_DATA_SIZE32_0 port map( sel => sig_bpw, din0(31) => 
                           s2_pc_sel_31_port, din0(30) => s2_pc_sel_30_port, 
                           din0(29) => s2_pc_sel_29_port, din0(28) => 
                           s2_pc_sel_28_port, din0(27) => s2_pc_sel_27_port, 
                           din0(26) => s2_pc_sel_26_port, din0(25) => 
                           s2_pc_sel_25_port, din0(24) => s2_pc_sel_24_port, 
                           din0(23) => s2_pc_sel_23_port, din0(22) => 
                           s2_pc_sel_22_port, din0(21) => s2_pc_sel_21_port, 
                           din0(20) => s2_pc_sel_20_port, din0(19) => 
                           s2_pc_sel_19_port, din0(18) => s2_pc_sel_18_port, 
                           din0(17) => s2_pc_sel_17_port, din0(16) => 
                           s2_pc_sel_16_port, din0(15) => s2_pc_sel_15_port, 
                           din0(14) => s2_pc_sel_14_port, din0(13) => 
                           s2_pc_sel_13_port, din0(12) => s2_pc_sel_12_port, 
                           din0(11) => s2_pc_sel_11_port, din0(10) => 
                           s2_pc_sel_10_port, din0(9) => s2_pc_sel_9_port, 
                           din0(8) => s2_pc_sel_8_port, din0(7) => 
                           s2_pc_sel_7_port, din0(6) => s2_pc_sel_6_port, 
                           din0(5) => s2_pc_sel_5_port, din0(4) => 
                           s2_pc_sel_4_port, din0(3) => s2_pc_sel_3_port, 
                           din0(2) => s2_pc_sel_2_port, din0(1) => 
                           s2_pc_sel_1_port, din0(0) => s2_pc_sel_0_port, 
                           din1(31) => s3_pc_notsel_31_port, din1(30) => 
                           s3_pc_notsel_30_port, din1(29) => 
                           s3_pc_notsel_29_port, din1(28) => 
                           s3_pc_notsel_28_port, din1(27) => 
                           s3_pc_notsel_27_port, din1(26) => 
                           s3_pc_notsel_26_port, din1(25) => 
                           s3_pc_notsel_25_port, din1(24) => 
                           s3_pc_notsel_24_port, din1(23) => 
                           s3_pc_notsel_23_port, din1(22) => 
                           s3_pc_notsel_22_port, din1(21) => 
                           s3_pc_notsel_21_port, din1(20) => 
                           s3_pc_notsel_20_port, din1(19) => 
                           s3_pc_notsel_19_port, din1(18) => 
                           s3_pc_notsel_18_port, din1(17) => 
                           s3_pc_notsel_17_port, din1(16) => 
                           s3_pc_notsel_16_port, din1(15) => 
                           s3_pc_notsel_15_port, din1(14) => 
                           s3_pc_notsel_14_port, din1(13) => 
                           s3_pc_notsel_13_port, din1(12) => 
                           s3_pc_notsel_12_port, din1(11) => 
                           s3_pc_notsel_11_port, din1(10) => 
                           s3_pc_notsel_10_port, din1(9) => s3_pc_notsel_9_port
                           , din1(8) => s3_pc_notsel_8_port, din1(7) => 
                           s3_pc_notsel_7_port, din1(6) => s3_pc_notsel_6_port,
                           din1(5) => s3_pc_notsel_5_port, din1(4) => 
                           s3_pc_notsel_4_port, din1(3) => s3_pc_notsel_3_port,
                           din1(2) => s3_pc_notsel_2_port, din1(1) => 
                           s3_pc_notsel_1_port, din1(0) => s3_pc_notsel_0_port,
                           dout(31) => istr_addr_31_port, dout(30) => 
                           istr_addr_30_port, dout(29) => istr_addr_29_port, 
                           dout(28) => istr_addr_28_port, dout(27) => 
                           istr_addr_27_port, dout(26) => istr_addr_26_port, 
                           dout(25) => istr_addr_25_port, dout(24) => 
                           istr_addr_24_port, dout(23) => istr_addr_23_port, 
                           dout(22) => istr_addr_22_port, dout(21) => 
                           istr_addr_21_port, dout(20) => istr_addr_20_port, 
                           dout(19) => istr_addr_19_port, dout(18) => 
                           istr_addr_18_port, dout(17) => istr_addr_17_port, 
                           dout(16) => istr_addr_16_port, dout(15) => 
                           istr_addr_15_port, dout(14) => istr_addr_14_port, 
                           dout(13) => istr_addr_13_port, dout(12) => 
                           istr_addr_12_port, dout(11) => istr_addr_11_port, 
                           dout(10) => istr_addr_10_port, dout(9) => 
                           istr_addr_9_port, dout(8) => istr_addr_8_port, 
                           dout(7) => istr_addr_7_port, dout(6) => 
                           istr_addr_6_port, dout(5) => istr_addr_5_port, 
                           dout(4) => istr_addr_4_port, dout(3) => 
                           istr_addr_3_port, dout(2) => istr_addr_2_port, 
                           dout(1) => istr_addr_1_port, dout(0) => 
                           istr_addr_0_port);
   REG_PC : Reg_DATA_SIZE32_0 port map( rst => rst, en => cw(0), clk => clk, 
                           din(31) => istr_addr_31_port, din(30) => 
                           istr_addr_30_port, din(29) => istr_addr_29_port, 
                           din(28) => istr_addr_28_port, din(27) => 
                           istr_addr_27_port, din(26) => istr_addr_26_port, 
                           din(25) => istr_addr_25_port, din(24) => 
                           istr_addr_24_port, din(23) => istr_addr_23_port, 
                           din(22) => istr_addr_22_port, din(21) => 
                           istr_addr_21_port, din(20) => istr_addr_20_port, 
                           din(19) => istr_addr_19_port, din(18) => 
                           istr_addr_18_port, din(17) => istr_addr_17_port, 
                           din(16) => istr_addr_16_port, din(15) => 
                           istr_addr_15_port, din(14) => istr_addr_14_port, 
                           din(13) => istr_addr_13_port, din(12) => 
                           istr_addr_12_port, din(11) => istr_addr_11_port, 
                           din(10) => istr_addr_10_port, din(9) => 
                           istr_addr_9_port, din(8) => istr_addr_8_port, din(7)
                           => istr_addr_7_port, din(6) => istr_addr_6_port, 
                           din(5) => istr_addr_5_port, din(4) => 
                           istr_addr_4_port, din(3) => istr_addr_3_port, din(2)
                           => istr_addr_2_port, din(1) => istr_addr_1_port, 
                           din(0) => istr_addr_0_port, dout(31) => pc_out(31), 
                           dout(30) => pc_out(30), dout(29) => pc_out(29), 
                           dout(28) => pc_out(28), dout(27) => pc_out(27), 
                           dout(26) => pc_out(26), dout(25) => pc_out(25), 
                           dout(24) => pc_out(24), dout(23) => pc_out(23), 
                           dout(22) => pc_out(22), dout(21) => pc_out(21), 
                           dout(20) => pc_out(20), dout(19) => pc_out(19), 
                           dout(18) => pc_out(18), dout(17) => pc_out(17), 
                           dout(16) => pc_out(16), dout(15) => pc_out(15), 
                           dout(14) => pc_out(14), dout(13) => pc_out(13), 
                           dout(12) => pc_out(12), dout(11) => pc_out(11), 
                           dout(10) => pc_out(10), dout(9) => pc_out(9), 
                           dout(8) => pc_out(8), dout(7) => pc_out(7), dout(6) 
                           => pc_out(6), dout(5) => pc_out(5), dout(4) => 
                           pc_out(4), dout(3) => pc_out(3), dout(2) => 
                           pc_out(2), dout(1) => pc_out(1), dout(0) => 
                           pc_out(0));
   REG_NPC : Reg_DATA_SIZE32_12 port map( rst => rst, en => cw(0), clk => clk, 
                           din(31) => s1_npc_31_port, din(30) => s1_npc_30_port
                           , din(29) => s1_npc_29_port, din(28) => 
                           s1_npc_28_port, din(27) => s1_npc_27_port, din(26) 
                           => s1_npc_26_port, din(25) => s1_npc_25_port, 
                           din(24) => s1_npc_24_port, din(23) => s1_npc_23_port
                           , din(22) => s1_npc_22_port, din(21) => 
                           s1_npc_21_port, din(20) => s1_npc_20_port, din(19) 
                           => s1_npc_19_port, din(18) => s1_npc_18_port, 
                           din(17) => s1_npc_17_port, din(16) => s1_npc_16_port
                           , din(15) => s1_npc_15_port, din(14) => 
                           s1_npc_14_port, din(13) => s1_npc_13_port, din(12) 
                           => s1_npc_12_port, din(11) => s1_npc_11_port, 
                           din(10) => s1_npc_10_port, din(9) => s1_npc_9_port, 
                           din(8) => s1_npc_8_port, din(7) => s1_npc_7_port, 
                           din(6) => s1_npc_6_port, din(5) => s1_npc_5_port, 
                           din(4) => s1_npc_4_port, din(3) => s1_npc_3_port, 
                           din(2) => s1_npc_2_port, din(1) => s1_npc_1_port, 
                           din(0) => s1_npc_0_port, dout(31) => s2_npc_31_port,
                           dout(30) => s2_npc_30_port, dout(29) => 
                           s2_npc_29_port, dout(28) => s2_npc_28_port, dout(27)
                           => s2_npc_27_port, dout(26) => s2_npc_26_port, 
                           dout(25) => s2_npc_25_port, dout(24) => 
                           s2_npc_24_port, dout(23) => s2_npc_23_port, dout(22)
                           => s2_npc_22_port, dout(21) => s2_npc_21_port, 
                           dout(20) => s2_npc_20_port, dout(19) => 
                           s2_npc_19_port, dout(18) => s2_npc_18_port, dout(17)
                           => s2_npc_17_port, dout(16) => s2_npc_16_port, 
                           dout(15) => s2_npc_15_port, dout(14) => 
                           s2_npc_14_port, dout(13) => s2_npc_13_port, dout(12)
                           => s2_npc_12_port, dout(11) => s2_npc_11_port, 
                           dout(10) => s2_npc_10_port, dout(9) => s2_npc_9_port
                           , dout(8) => s2_npc_8_port, dout(7) => s2_npc_7_port
                           , dout(6) => s2_npc_6_port, dout(5) => s2_npc_5_port
                           , dout(4) => s2_npc_4_port, dout(3) => s2_npc_3_port
                           , dout(2) => s2_npc_2_port, dout(1) => s2_npc_1_port
                           , dout(0) => s2_npc_0_port);
   MUX_PC : Mux_DATA_SIZE32_9 port map( sel => cw(1), din0(31) => 
                           s2_npc_31_port, din0(30) => s2_npc_30_port, din0(29)
                           => s2_npc_29_port, din0(28) => s2_npc_28_port, 
                           din0(27) => s2_npc_27_port, din0(26) => 
                           s2_npc_26_port, din0(25) => s2_npc_25_port, din0(24)
                           => s2_npc_24_port, din0(23) => s2_npc_23_port, 
                           din0(22) => s2_npc_22_port, din0(21) => 
                           s2_npc_21_port, din0(20) => s2_npc_20_port, din0(19)
                           => s2_npc_19_port, din0(18) => s2_npc_18_port, 
                           din0(17) => s2_npc_17_port, din0(16) => 
                           s2_npc_16_port, din0(15) => s2_npc_15_port, din0(14)
                           => s2_npc_14_port, din0(13) => s2_npc_13_port, 
                           din0(12) => s2_npc_12_port, din0(11) => 
                           s2_npc_11_port, din0(10) => s2_npc_10_port, din0(9) 
                           => s2_npc_9_port, din0(8) => s2_npc_8_port, din0(7) 
                           => s2_npc_7_port, din0(6) => s2_npc_6_port, din0(5) 
                           => s2_npc_5_port, din0(4) => s2_npc_4_port, din0(3) 
                           => s2_npc_3_port, din0(2) => s2_npc_2_port, din0(1) 
                           => s2_npc_1_port, din0(0) => s2_npc_0_port, din1(31)
                           => X_Logic0_port, din1(30) => s2_jpc_30_port, 
                           din1(29) => s2_jpc_29_port, din1(28) => 
                           s2_jpc_28_port, din1(27) => s2_jpc_27_port, din1(26)
                           => s2_jpc_26_port, din1(25) => s2_jpc_25_port, 
                           din1(24) => s2_jpc_24_port, din1(23) => 
                           s2_jpc_23_port, din1(22) => s2_jpc_22_port, din1(21)
                           => s2_jpc_21_port, din1(20) => s2_jpc_20_port, 
                           din1(19) => s2_jpc_19_port, din1(18) => 
                           s2_jpc_18_port, din1(17) => s2_jpc_17_port, din1(16)
                           => s2_jpc_16_port, din1(15) => s2_jpc_15_port, 
                           din1(14) => s2_jpc_14_port, din1(13) => 
                           s2_jpc_13_port, din1(12) => s2_jpc_12_port, din1(11)
                           => s2_jpc_11_port, din1(10) => s2_jpc_10_port, 
                           din1(9) => s2_jpc_9_port, din1(8) => s2_jpc_8_port, 
                           din1(7) => s2_jpc_7_port, din1(6) => s2_jpc_6_port, 
                           din1(5) => s2_jpc_5_port, din1(4) => s2_jpc_4_port, 
                           din1(3) => s2_jpc_3_port, din1(2) => s2_jpc_2_port, 
                           din1(1) => s2_jpc_1_port, din1(0) => s2_jpc_0_port, 
                           dout(31) => s2_pc_sel_31_port, dout(30) => 
                           s2_pc_sel_30_port, dout(29) => s2_pc_sel_29_port, 
                           dout(28) => s2_pc_sel_28_port, dout(27) => 
                           s2_pc_sel_27_port, dout(26) => s2_pc_sel_26_port, 
                           dout(25) => s2_pc_sel_25_port, dout(24) => 
                           s2_pc_sel_24_port, dout(23) => s2_pc_sel_23_port, 
                           dout(22) => s2_pc_sel_22_port, dout(21) => 
                           s2_pc_sel_21_port, dout(20) => s2_pc_sel_20_port, 
                           dout(19) => s2_pc_sel_19_port, dout(18) => 
                           s2_pc_sel_18_port, dout(17) => s2_pc_sel_17_port, 
                           dout(16) => s2_pc_sel_16_port, dout(15) => 
                           s2_pc_sel_15_port, dout(14) => s2_pc_sel_14_port, 
                           dout(13) => s2_pc_sel_13_port, dout(12) => 
                           s2_pc_sel_12_port, dout(11) => s2_pc_sel_11_port, 
                           dout(10) => s2_pc_sel_10_port, dout(9) => 
                           s2_pc_sel_9_port, dout(8) => s2_pc_sel_8_port, 
                           dout(7) => s2_pc_sel_7_port, dout(6) => 
                           s2_pc_sel_6_port, dout(5) => s2_pc_sel_5_port, 
                           dout(4) => s2_pc_sel_4_port, dout(3) => 
                           s2_pc_sel_3_port, dout(2) => s2_pc_sel_2_port, 
                           dout(1) => s2_pc_sel_1_port, dout(0) => 
                           s2_pc_sel_0_port);
   MUX_NOTPC : Mux_DATA_SIZE32_8 port map( sel => cw(1), din0(31) => 
                           X_Logic0_port, din0(30) => s2_jpc_30_port, din0(29) 
                           => s2_jpc_29_port, din0(28) => s2_jpc_28_port, 
                           din0(27) => s2_jpc_27_port, din0(26) => 
                           s2_jpc_26_port, din0(25) => s2_jpc_25_port, din0(24)
                           => s2_jpc_24_port, din0(23) => s2_jpc_23_port, 
                           din0(22) => s2_jpc_22_port, din0(21) => 
                           s2_jpc_21_port, din0(20) => s2_jpc_20_port, din0(19)
                           => s2_jpc_19_port, din0(18) => s2_jpc_18_port, 
                           din0(17) => s2_jpc_17_port, din0(16) => 
                           s2_jpc_16_port, din0(15) => s2_jpc_15_port, din0(14)
                           => s2_jpc_14_port, din0(13) => s2_jpc_13_port, 
                           din0(12) => s2_jpc_12_port, din0(11) => 
                           s2_jpc_11_port, din0(10) => s2_jpc_10_port, din0(9) 
                           => s2_jpc_9_port, din0(8) => s2_jpc_8_port, din0(7) 
                           => s2_jpc_7_port, din0(6) => s2_jpc_6_port, din0(5) 
                           => s2_jpc_5_port, din0(4) => s2_jpc_4_port, din0(3) 
                           => s2_jpc_3_port, din0(2) => s2_jpc_2_port, din0(1) 
                           => s2_jpc_1_port, din0(0) => s2_jpc_0_port, din1(31)
                           => s2_npc_31_port, din1(30) => s2_npc_30_port, 
                           din1(29) => s2_npc_29_port, din1(28) => 
                           s2_npc_28_port, din1(27) => s2_npc_27_port, din1(26)
                           => s2_npc_26_port, din1(25) => s2_npc_25_port, 
                           din1(24) => s2_npc_24_port, din1(23) => 
                           s2_npc_23_port, din1(22) => s2_npc_22_port, din1(21)
                           => s2_npc_21_port, din1(20) => s2_npc_20_port, 
                           din1(19) => s2_npc_19_port, din1(18) => 
                           s2_npc_18_port, din1(17) => s2_npc_17_port, din1(16)
                           => s2_npc_16_port, din1(15) => s2_npc_15_port, 
                           din1(14) => s2_npc_14_port, din1(13) => 
                           s2_npc_13_port, din1(12) => s2_npc_12_port, din1(11)
                           => s2_npc_11_port, din1(10) => s2_npc_10_port, 
                           din1(9) => s2_npc_9_port, din1(8) => s2_npc_8_port, 
                           din1(7) => s2_npc_7_port, din1(6) => s2_npc_6_port, 
                           din1(5) => s2_npc_5_port, din1(4) => s2_npc_4_port, 
                           din1(3) => s2_npc_3_port, din1(2) => s2_npc_2_port, 
                           din1(1) => s2_npc_1_port, din1(0) => s2_npc_0_port, 
                           dout(31) => s2_pc_notsel_31_port, dout(30) => 
                           s2_pc_notsel_30_port, dout(29) => 
                           s2_pc_notsel_29_port, dout(28) => 
                           s2_pc_notsel_28_port, dout(27) => 
                           s2_pc_notsel_27_port, dout(26) => 
                           s2_pc_notsel_26_port, dout(25) => 
                           s2_pc_notsel_25_port, dout(24) => 
                           s2_pc_notsel_24_port, dout(23) => 
                           s2_pc_notsel_23_port, dout(22) => 
                           s2_pc_notsel_22_port, dout(21) => 
                           s2_pc_notsel_21_port, dout(20) => 
                           s2_pc_notsel_20_port, dout(19) => 
                           s2_pc_notsel_19_port, dout(18) => 
                           s2_pc_notsel_18_port, dout(17) => 
                           s2_pc_notsel_17_port, dout(16) => 
                           s2_pc_notsel_16_port, dout(15) => 
                           s2_pc_notsel_15_port, dout(14) => 
                           s2_pc_notsel_14_port, dout(13) => 
                           s2_pc_notsel_13_port, dout(12) => 
                           s2_pc_notsel_12_port, dout(11) => 
                           s2_pc_notsel_11_port, dout(10) => 
                           s2_pc_notsel_10_port, dout(9) => s2_pc_notsel_9_port
                           , dout(8) => s2_pc_notsel_8_port, dout(7) => 
                           s2_pc_notsel_7_port, dout(6) => s2_pc_notsel_6_port,
                           dout(5) => s2_pc_notsel_5_port, dout(4) => 
                           s2_pc_notsel_4_port, dout(3) => s2_pc_notsel_3_port,
                           dout(2) => s2_pc_notsel_2_port, dout(1) => 
                           s2_pc_notsel_1_port, dout(0) => s2_pc_notsel_0_port)
                           ;
   MUX_WB_ADDR : Mux_DATA_SIZE5 port map( sel => s2_wr_addr_sel, din0(4) => 
                           istr_val(15), din0(3) => istr_val(14), din0(2) => 
                           istr_val(13), din0(1) => istr_val(12), din0(0) => 
                           istr_val(11), din1(4) => istr_val(20), din1(3) => 
                           istr_val(19), din1(2) => istr_val(18), din1(1) => 
                           istr_val(17), din1(0) => istr_val(16), dout(4) => 
                           s2_wr_addr_4_port, dout(3) => s2_wr_addr_3_port, 
                           dout(2) => s2_wr_addr_2_port, dout(1) => 
                           s2_wr_addr_1_port, dout(0) => s2_wr_addr_0_port);
   EXT_L : Extender_SRC_SIZE16_DEST_SIZE32 port map( s => cw(5), i(15) => 
                           istr_val(15), i(14) => istr_val(14), i(13) => 
                           istr_val(13), i(12) => istr_val(12), i(11) => 
                           istr_val(11), i(10) => istr_val(10), i(9) => 
                           istr_val(9), i(8) => istr_val(8), i(7) => 
                           istr_val(7), i(6) => istr_val(6), i(5) => 
                           istr_val(5), i(4) => istr_val(4), i(3) => 
                           istr_val(3), i(2) => istr_val(2), i(1) => 
                           istr_val(1), i(0) => istr_val(0), o(31) => 
                           s2_imm_l_ext_31_port, o(30) => net107975, o(29) => 
                           net107976, o(28) => net107977, o(27) => net107978, 
                           o(26) => net107979, o(25) => net107980, o(24) => 
                           net107981, o(23) => net107982, o(22) => net107983, 
                           o(21) => net107984, o(20) => net107985, o(19) => 
                           net107986, o(18) => net107987, o(17) => net107988, 
                           o(16) => net107989, o(15) => s2_imm_l_ext_15_port, 
                           o(14) => s2_imm_l_ext_14_port, o(13) => 
                           s2_imm_l_ext_13_port, o(12) => s2_imm_l_ext_12_port,
                           o(11) => s2_imm_l_ext_11_port, o(10) => 
                           s2_imm_l_ext_10_port, o(9) => s2_imm_l_ext_9_port, 
                           o(8) => s2_imm_l_ext_8_port, o(7) => 
                           s2_imm_l_ext_7_port, o(6) => s2_imm_l_ext_6_port, 
                           o(5) => s2_imm_l_ext_5_port, o(4) => 
                           s2_imm_l_ext_4_port, o(3) => s2_imm_l_ext_3_port, 
                           o(2) => s2_imm_l_ext_2_port, o(1) => 
                           s2_imm_l_ext_1_port, o(0) => s2_imm_l_ext_0_port);
   EXT_J : Extender_SRC_SIZE26_DEST_SIZE32 port map( s => X_Logic1_port, i(25) 
                           => istr_val(25), i(24) => istr_val(24), i(23) => 
                           istr_val(23), i(22) => istr_val(22), i(21) => 
                           istr_val(21), i(20) => istr_val(20), i(19) => 
                           istr_val(19), i(18) => istr_val(18), i(17) => 
                           istr_val(17), i(16) => istr_val(16), i(15) => 
                           istr_val(15), i(14) => istr_val(14), i(13) => 
                           istr_val(13), i(12) => istr_val(12), i(11) => 
                           istr_val(11), i(10) => istr_val(10), i(9) => 
                           istr_val(9), i(8) => istr_val(8), i(7) => 
                           istr_val(7), i(6) => istr_val(6), i(5) => 
                           istr_val(5), i(4) => istr_val(4), i(3) => 
                           istr_val(3), i(2) => istr_val(2), i(1) => 
                           istr_val(1), i(0) => istr_val(0), o(31) => 
                           s2_imm_j_ext_31_port, o(30) => s2_imm_j_ext_30_port,
                           o(29) => s2_imm_j_ext_29_port, o(28) => 
                           s2_imm_j_ext_28_port, o(27) => s2_imm_j_ext_27_port,
                           o(26) => s2_imm_j_ext_26_port, o(25) => 
                           s2_imm_j_ext_25_port, o(24) => s2_imm_j_ext_24_port,
                           o(23) => s2_imm_j_ext_23_port, o(22) => 
                           s2_imm_j_ext_22_port, o(21) => s2_imm_j_ext_21_port,
                           o(20) => s2_imm_j_ext_20_port, o(19) => 
                           s2_imm_j_ext_19_port, o(18) => s2_imm_j_ext_18_port,
                           o(17) => s2_imm_j_ext_17_port, o(16) => 
                           s2_imm_j_ext_16_port, o(15) => s2_imm_j_ext_15_port,
                           o(14) => s2_imm_j_ext_14_port, o(13) => 
                           s2_imm_j_ext_13_port, o(12) => s2_imm_j_ext_12_port,
                           o(11) => s2_imm_j_ext_11_port, o(10) => 
                           s2_imm_j_ext_10_port, o(9) => s2_imm_j_ext_9_port, 
                           o(8) => s2_imm_j_ext_8_port, o(7) => 
                           s2_imm_j_ext_7_port, o(6) => s2_imm_j_ext_6_port, 
                           o(5) => s2_imm_j_ext_5_port, o(4) => 
                           s2_imm_j_ext_4_port, o(3) => s2_imm_j_ext_3_port, 
                           o(2) => s2_imm_j_ext_2_port, o(1) => 
                           s2_imm_j_ext_1_port, o(0) => s2_imm_j_ext_0_port);
   RF0 : RegisterFile_DATA_SIZE32_REG_NUM32 port map( clk => clk, rst => rst, 
                           en => s2_rf_en, rd1_en => cw(6), rd2_en => cw(6), 
                           wr_en => cw(19), link_en => cw(4), rd1_addr(4) => 
                           istr_val(25), rd1_addr(3) => istr_val(24), 
                           rd1_addr(2) => istr_val(23), rd1_addr(1) => 
                           istr_val(22), rd1_addr(0) => istr_val(21), 
                           rd2_addr(4) => istr_val(20), rd2_addr(3) => 
                           istr_val(19), rd2_addr(2) => istr_val(18), 
                           rd2_addr(1) => istr_val(17), rd2_addr(0) => 
                           istr_val(16), wr_addr(4) => s5_wr_addr_4_port, 
                           wr_addr(3) => s5_wr_addr_3_port, wr_addr(2) => 
                           s5_wr_addr_2_port, wr_addr(1) => s5_wr_addr_1_port, 
                           wr_addr(0) => s5_wr_addr_0_port, d_out1(31) => 
                           s2_a_31_port, d_out1(30) => s2_a_30_port, d_out1(29)
                           => s2_a_29_port, d_out1(28) => s2_a_28_port, 
                           d_out1(27) => s2_a_27_port, d_out1(26) => 
                           s2_a_26_port, d_out1(25) => s2_a_25_port, d_out1(24)
                           => s2_a_24_port, d_out1(23) => s2_a_23_port, 
                           d_out1(22) => s2_a_22_port, d_out1(21) => 
                           s2_a_21_port, d_out1(20) => s2_a_20_port, d_out1(19)
                           => s2_a_19_port, d_out1(18) => s2_a_18_port, 
                           d_out1(17) => s2_a_17_port, d_out1(16) => 
                           s2_a_16_port, d_out1(15) => s2_a_15_port, d_out1(14)
                           => s2_a_14_port, d_out1(13) => s2_a_13_port, 
                           d_out1(12) => s2_a_12_port, d_out1(11) => 
                           s2_a_11_port, d_out1(10) => s2_a_10_port, d_out1(9) 
                           => s2_a_9_port, d_out1(8) => s2_a_8_port, d_out1(7) 
                           => s2_a_7_port, d_out1(6) => s2_a_6_port, d_out1(5) 
                           => s2_a_5_port, d_out1(4) => s2_a_4_port, d_out1(3) 
                           => s2_a_3_port, d_out1(2) => s2_a_2_port, d_out1(1) 
                           => s2_a_1_port, d_out1(0) => s2_a_0_port, d_out2(31)
                           => s2_b_31_port, d_out2(30) => s2_b_30_port, 
                           d_out2(29) => s2_b_29_port, d_out2(28) => 
                           s2_b_28_port, d_out2(27) => s2_b_27_port, d_out2(26)
                           => s2_b_26_port, d_out2(25) => s2_b_25_port, 
                           d_out2(24) => s2_b_24_port, d_out2(23) => 
                           s2_b_23_port, d_out2(22) => s2_b_22_port, d_out2(21)
                           => s2_b_21_port, d_out2(20) => s2_b_20_port, 
                           d_out2(19) => s2_b_19_port, d_out2(18) => 
                           s2_b_18_port, d_out2(17) => s2_b_17_port, d_out2(16)
                           => s2_b_16_port, d_out2(15) => s2_b_15_port, 
                           d_out2(14) => s2_b_14_port, d_out2(13) => 
                           s2_b_13_port, d_out2(12) => s2_b_12_port, d_out2(11)
                           => s2_b_11_port, d_out2(10) => s2_b_10_port, 
                           d_out2(9) => s2_b_9_port, d_out2(8) => s2_b_8_port, 
                           d_out2(7) => s2_b_7_port, d_out2(6) => s2_b_6_port, 
                           d_out2(5) => s2_b_5_port, d_out2(4) => s2_b_4_port, 
                           d_out2(3) => s2_b_3_port, d_out2(2) => s2_b_2_port, 
                           d_out2(1) => s2_b_1_port, d_out2(0) => s2_b_0_port, 
                           d_in(31) => s5_result_31_port, d_in(30) => 
                           s5_result_30_port, d_in(29) => s5_result_29_port, 
                           d_in(28) => s5_result_28_port, d_in(27) => 
                           s5_result_27_port, d_in(26) => s5_result_26_port, 
                           d_in(25) => s5_result_25_port, d_in(24) => 
                           s5_result_24_port, d_in(23) => s5_result_23_port, 
                           d_in(22) => s5_result_22_port, d_in(21) => 
                           s5_result_21_port, d_in(20) => s5_result_20_port, 
                           d_in(19) => s5_result_19_port, d_in(18) => 
                           s5_result_18_port, d_in(17) => s5_result_17_port, 
                           d_in(16) => s5_result_16_port, d_in(15) => 
                           s5_result_15_port, d_in(14) => s5_result_14_port, 
                           d_in(13) => s5_result_13_port, d_in(12) => 
                           s5_result_12_port, d_in(11) => s5_result_11_port, 
                           d_in(10) => s5_result_10_port, d_in(9) => 
                           s5_result_9_port, d_in(8) => s5_result_8_port, 
                           d_in(7) => s5_result_7_port, d_in(6) => 
                           s5_result_6_port, d_in(5) => s5_result_5_port, 
                           d_in(4) => s5_result_4_port, d_in(3) => 
                           s5_result_3_port, d_in(2) => s5_result_2_port, 
                           d_in(1) => s5_result_1_port, d_in(0) => 
                           s5_result_0_port, d_link(31) => s2_npc_31_port, 
                           d_link(30) => s2_npc_30_port, d_link(29) => 
                           s2_npc_29_port, d_link(28) => s2_npc_28_port, 
                           d_link(27) => s2_npc_27_port, d_link(26) => 
                           s2_npc_26_port, d_link(25) => s2_npc_25_port, 
                           d_link(24) => s2_npc_24_port, d_link(23) => 
                           s2_npc_23_port, d_link(22) => s2_npc_22_port, 
                           d_link(21) => s2_npc_21_port, d_link(20) => 
                           s2_npc_20_port, d_link(19) => s2_npc_19_port, 
                           d_link(18) => s2_npc_18_port, d_link(17) => 
                           s2_npc_17_port, d_link(16) => s2_npc_16_port, 
                           d_link(15) => s2_npc_15_port, d_link(14) => 
                           s2_npc_14_port, d_link(13) => s2_npc_13_port, 
                           d_link(12) => s2_npc_12_port, d_link(11) => 
                           s2_npc_11_port, d_link(10) => s2_npc_10_port, 
                           d_link(9) => s2_npc_9_port, d_link(8) => 
                           s2_npc_8_port, d_link(7) => s2_npc_7_port, d_link(6)
                           => s2_npc_6_port, d_link(5) => s2_npc_5_port, 
                           d_link(4) => s2_npc_4_port, d_link(3) => 
                           s2_npc_3_port, d_link(2) => s2_npc_2_port, d_link(1)
                           => s2_npc_1_port, d_link(0) => s2_npc_0_port);
   MUX_JPC0 : Mux_DATA_SIZE32_7 port map( sel => cw(2), din0(31) => 
                           s2_imm_i_ext_31_port, din0(30) => 
                           s2_imm_i_ext_30_port, din0(29) => 
                           s2_imm_i_ext_29_port, din0(28) => 
                           s2_imm_i_ext_28_port, din0(27) => 
                           s2_imm_i_ext_27_port, din0(26) => 
                           s2_imm_i_ext_26_port, din0(25) => 
                           s2_imm_i_ext_25_port, din0(24) => 
                           s2_imm_i_ext_24_port, din0(23) => 
                           s2_imm_i_ext_23_port, din0(22) => 
                           s2_imm_i_ext_22_port, din0(21) => 
                           s2_imm_i_ext_21_port, din0(20) => 
                           s2_imm_i_ext_20_port, din0(19) => 
                           s2_imm_i_ext_19_port, din0(18) => 
                           s2_imm_i_ext_18_port, din0(17) => 
                           s2_imm_i_ext_17_port, din0(16) => 
                           s2_imm_i_ext_16_port, din0(15) => 
                           s2_imm_i_ext_15_port, din0(14) => 
                           s2_imm_i_ext_14_port, din0(13) => 
                           s2_imm_i_ext_13_port, din0(12) => 
                           s2_imm_i_ext_12_port, din0(11) => 
                           s2_imm_i_ext_11_port, din0(10) => 
                           s2_imm_i_ext_10_port, din0(9) => s2_imm_i_ext_9_port
                           , din0(8) => s2_imm_i_ext_8_port, din0(7) => 
                           s2_imm_i_ext_7_port, din0(6) => s2_imm_i_ext_6_port,
                           din0(5) => s2_imm_i_ext_5_port, din0(4) => 
                           s2_imm_i_ext_4_port, din0(3) => s2_imm_i_ext_3_port,
                           din0(2) => s2_imm_i_ext_2_port, din0(1) => 
                           s2_imm_i_ext_1_port, din0(0) => s2_imm_i_ext_0_port,
                           din1(31) => s2_imm_j_ext_31_port, din1(30) => 
                           s2_imm_j_ext_30_port, din1(29) => 
                           s2_imm_j_ext_29_port, din1(28) => 
                           s2_imm_j_ext_28_port, din1(27) => 
                           s2_imm_j_ext_27_port, din1(26) => 
                           s2_imm_j_ext_26_port, din1(25) => 
                           s2_imm_j_ext_25_port, din1(24) => 
                           s2_imm_j_ext_24_port, din1(23) => 
                           s2_imm_j_ext_23_port, din1(22) => 
                           s2_imm_j_ext_22_port, din1(21) => 
                           s2_imm_j_ext_21_port, din1(20) => 
                           s2_imm_j_ext_20_port, din1(19) => 
                           s2_imm_j_ext_19_port, din1(18) => 
                           s2_imm_j_ext_18_port, din1(17) => 
                           s2_imm_j_ext_17_port, din1(16) => 
                           s2_imm_j_ext_16_port, din1(15) => 
                           s2_imm_j_ext_15_port, din1(14) => 
                           s2_imm_j_ext_14_port, din1(13) => 
                           s2_imm_j_ext_13_port, din1(12) => 
                           s2_imm_j_ext_12_port, din1(11) => 
                           s2_imm_j_ext_11_port, din1(10) => 
                           s2_imm_j_ext_10_port, din1(9) => s2_imm_j_ext_9_port
                           , din1(8) => s2_imm_j_ext_8_port, din1(7) => 
                           s2_imm_j_ext_7_port, din1(6) => s2_imm_j_ext_6_port,
                           din1(5) => s2_imm_j_ext_5_port, din1(4) => 
                           s2_imm_j_ext_4_port, din1(3) => s2_imm_j_ext_3_port,
                           din1(2) => s2_imm_j_ext_2_port, din1(1) => 
                           s2_imm_j_ext_1_port, din1(0) => s2_imm_j_ext_0_port,
                           dout(31) => s2_jump_addr_imm_31_port, dout(30) => 
                           s2_jump_addr_imm_30_port, dout(29) => 
                           s2_jump_addr_imm_29_port, dout(28) => 
                           s2_jump_addr_imm_28_port, dout(27) => 
                           s2_jump_addr_imm_27_port, dout(26) => 
                           s2_jump_addr_imm_26_port, dout(25) => 
                           s2_jump_addr_imm_25_port, dout(24) => 
                           s2_jump_addr_imm_24_port, dout(23) => 
                           s2_jump_addr_imm_23_port, dout(22) => 
                           s2_jump_addr_imm_22_port, dout(21) => 
                           s2_jump_addr_imm_21_port, dout(20) => 
                           s2_jump_addr_imm_20_port, dout(19) => 
                           s2_jump_addr_imm_19_port, dout(18) => 
                           s2_jump_addr_imm_18_port, dout(17) => 
                           s2_jump_addr_imm_17_port, dout(16) => 
                           s2_jump_addr_imm_16_port, dout(15) => 
                           s2_jump_addr_imm_15_port, dout(14) => 
                           s2_jump_addr_imm_14_port, dout(13) => 
                           s2_jump_addr_imm_13_port, dout(12) => 
                           s2_jump_addr_imm_12_port, dout(11) => 
                           s2_jump_addr_imm_11_port, dout(10) => 
                           s2_jump_addr_imm_10_port, dout(9) => 
                           s2_jump_addr_imm_9_port, dout(8) => 
                           s2_jump_addr_imm_8_port, dout(7) => 
                           s2_jump_addr_imm_7_port, dout(6) => 
                           s2_jump_addr_imm_6_port, dout(5) => 
                           s2_jump_addr_imm_5_port, dout(4) => 
                           s2_jump_addr_imm_4_port, dout(3) => 
                           s2_jump_addr_imm_3_port, dout(2) => 
                           s2_jump_addr_imm_2_port, dout(1) => 
                           s2_jump_addr_imm_1_port, dout(0) => 
                           s2_jump_addr_imm_0_port);
   ADDER_ADDR : Adder_DATA_SIZE32_7 port map( cin => X_Logic0_port, a(31) => 
                           s2_npc_31_port, a(30) => s2_npc_30_port, a(29) => 
                           s2_npc_29_port, a(28) => s2_npc_28_port, a(27) => 
                           s2_npc_27_port, a(26) => s2_npc_26_port, a(25) => 
                           s2_npc_25_port, a(24) => s2_npc_24_port, a(23) => 
                           s2_npc_23_port, a(22) => s2_npc_22_port, a(21) => 
                           s2_npc_21_port, a(20) => s2_npc_20_port, a(19) => 
                           s2_npc_19_port, a(18) => s2_npc_18_port, a(17) => 
                           s2_npc_17_port, a(16) => s2_npc_16_port, a(15) => 
                           s2_npc_15_port, a(14) => s2_npc_14_port, a(13) => 
                           s2_npc_13_port, a(12) => s2_npc_12_port, a(11) => 
                           s2_npc_11_port, a(10) => s2_npc_10_port, a(9) => 
                           s2_npc_9_port, a(8) => s2_npc_8_port, a(7) => 
                           s2_npc_7_port, a(6) => s2_npc_6_port, a(5) => 
                           s2_npc_5_port, a(4) => s2_npc_4_port, a(3) => 
                           s2_npc_3_port, a(2) => s2_npc_2_port, a(1) => 
                           s2_npc_1_port, a(0) => s2_npc_0_port, b(31) => 
                           s2_jump_addr_imm_31_port, b(30) => 
                           s2_jump_addr_imm_30_port, b(29) => 
                           s2_jump_addr_imm_29_port, b(28) => 
                           s2_jump_addr_imm_28_port, b(27) => 
                           s2_jump_addr_imm_27_port, b(26) => 
                           s2_jump_addr_imm_26_port, b(25) => 
                           s2_jump_addr_imm_25_port, b(24) => 
                           s2_jump_addr_imm_24_port, b(23) => 
                           s2_jump_addr_imm_23_port, b(22) => 
                           s2_jump_addr_imm_22_port, b(21) => 
                           s2_jump_addr_imm_21_port, b(20) => 
                           s2_jump_addr_imm_20_port, b(19) => 
                           s2_jump_addr_imm_19_port, b(18) => 
                           s2_jump_addr_imm_18_port, b(17) => 
                           s2_jump_addr_imm_17_port, b(16) => 
                           s2_jump_addr_imm_16_port, b(15) => 
                           s2_jump_addr_imm_15_port, b(14) => 
                           s2_jump_addr_imm_14_port, b(13) => 
                           s2_jump_addr_imm_13_port, b(12) => 
                           s2_jump_addr_imm_12_port, b(11) => 
                           s2_jump_addr_imm_11_port, b(10) => 
                           s2_jump_addr_imm_10_port, b(9) => 
                           s2_jump_addr_imm_9_port, b(8) => 
                           s2_jump_addr_imm_8_port, b(7) => 
                           s2_jump_addr_imm_7_port, b(6) => 
                           s2_jump_addr_imm_6_port, b(5) => 
                           s2_jump_addr_imm_5_port, b(4) => 
                           s2_jump_addr_imm_4_port, b(3) => 
                           s2_jump_addr_imm_3_port, b(2) => 
                           s2_jump_addr_imm_2_port, b(1) => 
                           s2_jump_addr_imm_1_port, b(0) => 
                           s2_jump_addr_imm_0_port, s(31) => 
                           s2_jump_addr_rel_31_port, s(30) => 
                           s2_jump_addr_rel_30_port, s(29) => 
                           s2_jump_addr_rel_29_port, s(28) => 
                           s2_jump_addr_rel_28_port, s(27) => 
                           s2_jump_addr_rel_27_port, s(26) => 
                           s2_jump_addr_rel_26_port, s(25) => 
                           s2_jump_addr_rel_25_port, s(24) => 
                           s2_jump_addr_rel_24_port, s(23) => 
                           s2_jump_addr_rel_23_port, s(22) => 
                           s2_jump_addr_rel_22_port, s(21) => 
                           s2_jump_addr_rel_21_port, s(20) => 
                           s2_jump_addr_rel_20_port, s(19) => 
                           s2_jump_addr_rel_19_port, s(18) => 
                           s2_jump_addr_rel_18_port, s(17) => 
                           s2_jump_addr_rel_17_port, s(16) => 
                           s2_jump_addr_rel_16_port, s(15) => 
                           s2_jump_addr_rel_15_port, s(14) => 
                           s2_jump_addr_rel_14_port, s(13) => 
                           s2_jump_addr_rel_13_port, s(12) => 
                           s2_jump_addr_rel_12_port, s(11) => 
                           s2_jump_addr_rel_11_port, s(10) => 
                           s2_jump_addr_rel_10_port, s(9) => 
                           s2_jump_addr_rel_9_port, s(8) => 
                           s2_jump_addr_rel_8_port, s(7) => 
                           s2_jump_addr_rel_7_port, s(6) => 
                           s2_jump_addr_rel_6_port, s(5) => 
                           s2_jump_addr_rel_5_port, s(4) => 
                           s2_jump_addr_rel_4_port, s(3) => 
                           s2_jump_addr_rel_3_port, s(2) => 
                           s2_jump_addr_rel_2_port, s(1) => 
                           s2_jump_addr_rel_1_port, s(0) => 
                           s2_jump_addr_rel_0_port, cout => net1293);
   MUX_JPC1 : Mux_DATA_SIZE32_6 port map( sel => cw(3), din0(31) => 
                           s2_jump_addr_rel_31_port, din0(30) => 
                           s2_jump_addr_rel_30_port, din0(29) => 
                           s2_jump_addr_rel_29_port, din0(28) => 
                           s2_jump_addr_rel_28_port, din0(27) => 
                           s2_jump_addr_rel_27_port, din0(26) => 
                           s2_jump_addr_rel_26_port, din0(25) => 
                           s2_jump_addr_rel_25_port, din0(24) => 
                           s2_jump_addr_rel_24_port, din0(23) => 
                           s2_jump_addr_rel_23_port, din0(22) => 
                           s2_jump_addr_rel_22_port, din0(21) => 
                           s2_jump_addr_rel_21_port, din0(20) => 
                           s2_jump_addr_rel_20_port, din0(19) => 
                           s2_jump_addr_rel_19_port, din0(18) => 
                           s2_jump_addr_rel_18_port, din0(17) => 
                           s2_jump_addr_rel_17_port, din0(16) => 
                           s2_jump_addr_rel_16_port, din0(15) => 
                           s2_jump_addr_rel_15_port, din0(14) => 
                           s2_jump_addr_rel_14_port, din0(13) => 
                           s2_jump_addr_rel_13_port, din0(12) => 
                           s2_jump_addr_rel_12_port, din0(11) => 
                           s2_jump_addr_rel_11_port, din0(10) => 
                           s2_jump_addr_rel_10_port, din0(9) => 
                           s2_jump_addr_rel_9_port, din0(8) => 
                           s2_jump_addr_rel_8_port, din0(7) => 
                           s2_jump_addr_rel_7_port, din0(6) => 
                           s2_jump_addr_rel_6_port, din0(5) => 
                           s2_jump_addr_rel_5_port, din0(4) => 
                           s2_jump_addr_rel_4_port, din0(3) => 
                           s2_jump_addr_rel_3_port, din0(2) => 
                           s2_jump_addr_rel_2_port, din0(1) => 
                           s2_jump_addr_rel_1_port, din0(0) => 
                           s2_jump_addr_rel_0_port, din1(31) => 
                           s2_jump_addr_reg_31_port, din1(30) => 
                           s2_jump_addr_reg_30_port, din1(29) => 
                           s2_jump_addr_reg_29_port, din1(28) => 
                           s2_jump_addr_reg_28_port, din1(27) => 
                           s2_jump_addr_reg_27_port, din1(26) => 
                           s2_jump_addr_reg_26_port, din1(25) => 
                           s2_jump_addr_reg_25_port, din1(24) => 
                           s2_jump_addr_reg_24_port, din1(23) => 
                           s2_jump_addr_reg_23_port, din1(22) => 
                           s2_jump_addr_reg_22_port, din1(21) => 
                           s2_jump_addr_reg_21_port, din1(20) => 
                           s2_jump_addr_reg_20_port, din1(19) => 
                           s2_jump_addr_reg_19_port, din1(18) => 
                           s2_jump_addr_reg_18_port, din1(17) => 
                           s2_jump_addr_reg_17_port, din1(16) => 
                           s2_jump_addr_reg_16_port, din1(15) => 
                           s2_jump_addr_reg_15_port, din1(14) => 
                           s2_jump_addr_reg_14_port, din1(13) => 
                           s2_jump_addr_reg_13_port, din1(12) => 
                           s2_jump_addr_reg_12_port, din1(11) => 
                           s2_jump_addr_reg_11_port, din1(10) => 
                           s2_jump_addr_reg_10_port, din1(9) => 
                           s2_jump_addr_reg_9_port, din1(8) => 
                           s2_jump_addr_reg_8_port, din1(7) => 
                           s2_jump_addr_reg_7_port, din1(6) => 
                           s2_jump_addr_reg_6_port, din1(5) => 
                           s2_jump_addr_reg_5_port, din1(4) => 
                           s2_jump_addr_reg_4_port, din1(3) => 
                           s2_jump_addr_reg_3_port, din1(2) => 
                           s2_jump_addr_reg_2_port, din1(1) => 
                           s2_jump_addr_reg_1_port, din1(0) => 
                           s2_jump_addr_reg_0_port, dout(31) => net1292, 
                           dout(30) => s2_jpc_30_port, dout(29) => 
                           s2_jpc_29_port, dout(28) => s2_jpc_28_port, dout(27)
                           => s2_jpc_27_port, dout(26) => s2_jpc_26_port, 
                           dout(25) => s2_jpc_25_port, dout(24) => 
                           s2_jpc_24_port, dout(23) => s2_jpc_23_port, dout(22)
                           => s2_jpc_22_port, dout(21) => s2_jpc_21_port, 
                           dout(20) => s2_jpc_20_port, dout(19) => 
                           s2_jpc_19_port, dout(18) => s2_jpc_18_port, dout(17)
                           => s2_jpc_17_port, dout(16) => s2_jpc_16_port, 
                           dout(15) => s2_jpc_15_port, dout(14) => 
                           s2_jpc_14_port, dout(13) => s2_jpc_13_port, dout(12)
                           => s2_jpc_12_port, dout(11) => s2_jpc_11_port, 
                           dout(10) => s2_jpc_10_port, dout(9) => s2_jpc_9_port
                           , dout(8) => s2_jpc_8_port, dout(7) => s2_jpc_7_port
                           , dout(6) => s2_jpc_6_port, dout(5) => s2_jpc_5_port
                           , dout(4) => s2_jpc_4_port, dout(3) => s2_jpc_3_port
                           , dout(2) => s2_jpc_2_port, dout(1) => s2_jpc_1_port
                           , dout(0) => s2_jpc_0_port);
   FWDMUX_2AB : FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_0 port map( reg_c(31) => 
                           s2_a_31_port, reg_c(30) => s2_a_30_port, reg_c(29) 
                           => s2_a_29_port, reg_c(28) => s2_a_28_port, 
                           reg_c(27) => s2_a_27_port, reg_c(26) => s2_a_26_port
                           , reg_c(25) => s2_a_25_port, reg_c(24) => 
                           s2_a_24_port, reg_c(23) => s2_a_23_port, reg_c(22) 
                           => s2_a_22_port, reg_c(21) => s2_a_21_port, 
                           reg_c(20) => s2_a_20_port, reg_c(19) => s2_a_19_port
                           , reg_c(18) => s2_a_18_port, reg_c(17) => 
                           s2_a_17_port, reg_c(16) => s2_a_16_port, reg_c(15) 
                           => s2_a_15_port, reg_c(14) => s2_a_14_port, 
                           reg_c(13) => s2_a_13_port, reg_c(12) => s2_a_12_port
                           , reg_c(11) => s2_a_11_port, reg_c(10) => 
                           s2_a_10_port, reg_c(9) => s2_a_9_port, reg_c(8) => 
                           s2_a_8_port, reg_c(7) => s2_a_7_port, reg_c(6) => 
                           s2_a_6_port, reg_c(5) => s2_a_5_port, reg_c(4) => 
                           s2_a_4_port, reg_c(3) => s2_a_3_port, reg_c(2) => 
                           s2_a_2_port, reg_c(1) => s2_a_1_port, reg_c(0) => 
                           s2_a_0_port, reg_f(31) => s3_exe_out_31_port, 
                           reg_f(30) => s3_exe_out_30_port, reg_f(29) => 
                           s3_exe_out_29_port, reg_f(28) => s3_exe_out_28_port,
                           reg_f(27) => s3_exe_out_27_port, reg_f(26) => 
                           s3_exe_out_26_port, reg_f(25) => s3_exe_out_25_port,
                           reg_f(24) => s3_exe_out_24_port, reg_f(23) => 
                           s3_exe_out_23_port, reg_f(22) => s3_exe_out_22_port,
                           reg_f(21) => s3_exe_out_21_port, reg_f(20) => 
                           s3_exe_out_20_port, reg_f(19) => s3_exe_out_19_port,
                           reg_f(18) => s3_exe_out_18_port, reg_f(17) => 
                           s3_exe_out_17_port, reg_f(16) => s3_exe_out_16_port,
                           reg_f(15) => s3_exe_out_15_port, reg_f(14) => 
                           s3_exe_out_14_port, reg_f(13) => s3_exe_out_13_port,
                           reg_f(12) => s3_exe_out_12_port, reg_f(11) => 
                           s3_exe_out_11_port, reg_f(10) => s3_exe_out_10_port,
                           reg_f(9) => s3_exe_out_9_port, reg_f(8) => 
                           s3_exe_out_8_port, reg_f(7) => s3_exe_out_7_port, 
                           reg_f(6) => s3_exe_out_6_port, reg_f(5) => 
                           s3_exe_out_5_port, reg_f(4) => s3_exe_out_4_port, 
                           reg_f(3) => s3_exe_out_3_port, reg_f(2) => 
                           s3_exe_out_2_port, reg_f(1) => s3_exe_out_1_port, 
                           reg_f(0) => s3_exe_out_0_port, reg_ff(31) => 
                           s4_result_31_port, reg_ff(30) => s4_result_30_port, 
                           reg_ff(29) => s4_result_29_port, reg_ff(28) => 
                           s4_result_28_port, reg_ff(27) => s4_result_27_port, 
                           reg_ff(26) => s4_result_26_port, reg_ff(25) => 
                           s4_result_25_port, reg_ff(24) => s4_result_24_port, 
                           reg_ff(23) => s4_result_23_port, reg_ff(22) => 
                           s4_result_22_port, reg_ff(21) => s4_result_21_port, 
                           reg_ff(20) => s4_result_20_port, reg_ff(19) => 
                           s4_result_19_port, reg_ff(18) => s4_result_18_port, 
                           reg_ff(17) => s4_result_17_port, reg_ff(16) => 
                           s4_result_16_port, reg_ff(15) => s4_result_15_port, 
                           reg_ff(14) => s4_result_14_port, reg_ff(13) => 
                           s4_result_13_port, reg_ff(12) => s4_result_12_port, 
                           reg_ff(11) => s4_result_11_port, reg_ff(10) => 
                           s4_result_10_port, reg_ff(9) => s4_result_9_port, 
                           reg_ff(8) => s4_result_8_port, reg_ff(7) => 
                           s4_result_7_port, reg_ff(6) => s4_result_6_port, 
                           reg_ff(5) => s4_result_5_port, reg_ff(4) => 
                           s4_result_4_port, reg_ff(3) => s4_result_3_port, 
                           reg_ff(2) => s4_result_2_port, reg_ff(1) => 
                           s4_result_1_port, reg_ff(0) => s4_result_0_port, 
                           addr_c(4) => istr_val(25), addr_c(3) => istr_val(24)
                           , addr_c(2) => istr_val(23), addr_c(1) => 
                           istr_val(22), addr_c(0) => istr_val(21), addr_f(4) 
                           => s3_wr_addr_4_port, addr_f(3) => s3_wr_addr_3_port
                           , addr_f(2) => s3_wr_addr_2_port, addr_f(1) => 
                           s3_wr_addr_1_port, addr_f(0) => s3_wr_addr_0_port, 
                           addr_ff(4) => s4_wr_addr_4_port, addr_ff(3) => 
                           s4_wr_addr_3_port, addr_ff(2) => s4_wr_addr_2_port, 
                           addr_ff(1) => s4_wr_addr_1_port, addr_ff(0) => 
                           s4_wr_addr_0_port, valid_f => s2_a_f_b_en, valid_ff 
                           => s2_a_ff_b_en, dirty_f => cw(8), dirty_ff => 
                           X_Logic0_port, en => X_Logic1_port, output(31) => 
                           reg_a_out(31), output(30) => reg_a_out(30), 
                           output(29) => reg_a_out(29), output(28) => 
                           reg_a_out(28), output(27) => reg_a_out(27), 
                           output(26) => reg_a_out(26), output(25) => 
                           reg_a_out(25), output(24) => reg_a_out(24), 
                           output(23) => reg_a_out(23), output(22) => 
                           reg_a_out(22), output(21) => reg_a_out(21), 
                           output(20) => reg_a_out(20), output(19) => 
                           reg_a_out(19), output(18) => reg_a_out(18), 
                           output(17) => reg_a_out(17), output(16) => 
                           reg_a_out(16), output(15) => reg_a_out(15), 
                           output(14) => reg_a_out(14), output(13) => 
                           reg_a_out(13), output(12) => reg_a_out(12), 
                           output(11) => reg_a_out(11), output(10) => 
                           reg_a_out(10), output(9) => reg_a_out(9), output(8) 
                           => reg_a_out(8), output(7) => reg_a_out(7), 
                           output(6) => reg_a_out(6), output(5) => reg_a_out(5)
                           , output(4) => reg_a_out(4), output(3) => 
                           reg_a_out(3), output(2) => reg_a_out(2), output(1) 
                           => reg_a_out(1), output(0) => reg_a_out(0), 
                           match_dirty_f => sig_bal, match_dirty_ff => net1291)
                           ;
   FWDMUX_2AJ : FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_4 port map( reg_c(31) => 
                           s2_a_31_port, reg_c(30) => s2_a_30_port, reg_c(29) 
                           => s2_a_29_port, reg_c(28) => s2_a_28_port, 
                           reg_c(27) => s2_a_27_port, reg_c(26) => s2_a_26_port
                           , reg_c(25) => s2_a_25_port, reg_c(24) => 
                           s2_a_24_port, reg_c(23) => s2_a_23_port, reg_c(22) 
                           => s2_a_22_port, reg_c(21) => s2_a_21_port, 
                           reg_c(20) => s2_a_20_port, reg_c(19) => s2_a_19_port
                           , reg_c(18) => s2_a_18_port, reg_c(17) => 
                           s2_a_17_port, reg_c(16) => s2_a_16_port, reg_c(15) 
                           => s2_a_15_port, reg_c(14) => s2_a_14_port, 
                           reg_c(13) => s2_a_13_port, reg_c(12) => s2_a_12_port
                           , reg_c(11) => s2_a_11_port, reg_c(10) => 
                           s2_a_10_port, reg_c(9) => s2_a_9_port, reg_c(8) => 
                           s2_a_8_port, reg_c(7) => s2_a_7_port, reg_c(6) => 
                           s2_a_6_port, reg_c(5) => s2_a_5_port, reg_c(4) => 
                           s2_a_4_port, reg_c(3) => s2_a_3_port, reg_c(2) => 
                           s2_a_2_port, reg_c(1) => s2_a_1_port, reg_c(0) => 
                           s2_a_0_port, reg_f(31) => s3_exe_out_31_port, 
                           reg_f(30) => s3_exe_out_30_port, reg_f(29) => 
                           s3_exe_out_29_port, reg_f(28) => s3_exe_out_28_port,
                           reg_f(27) => s3_exe_out_27_port, reg_f(26) => 
                           s3_exe_out_26_port, reg_f(25) => s3_exe_out_25_port,
                           reg_f(24) => s3_exe_out_24_port, reg_f(23) => 
                           s3_exe_out_23_port, reg_f(22) => s3_exe_out_22_port,
                           reg_f(21) => s3_exe_out_21_port, reg_f(20) => 
                           s3_exe_out_20_port, reg_f(19) => s3_exe_out_19_port,
                           reg_f(18) => s3_exe_out_18_port, reg_f(17) => 
                           s3_exe_out_17_port, reg_f(16) => s3_exe_out_16_port,
                           reg_f(15) => s3_exe_out_15_port, reg_f(14) => 
                           s3_exe_out_14_port, reg_f(13) => s3_exe_out_13_port,
                           reg_f(12) => s3_exe_out_12_port, reg_f(11) => 
                           s3_exe_out_11_port, reg_f(10) => s3_exe_out_10_port,
                           reg_f(9) => s3_exe_out_9_port, reg_f(8) => 
                           s3_exe_out_8_port, reg_f(7) => s3_exe_out_7_port, 
                           reg_f(6) => s3_exe_out_6_port, reg_f(5) => 
                           s3_exe_out_5_port, reg_f(4) => s3_exe_out_4_port, 
                           reg_f(3) => s3_exe_out_3_port, reg_f(2) => 
                           s3_exe_out_2_port, reg_f(1) => s3_exe_out_1_port, 
                           reg_f(0) => s3_exe_out_0_port, reg_ff(31) => 
                           s4_result_31_port, reg_ff(30) => s4_result_30_port, 
                           reg_ff(29) => s4_result_29_port, reg_ff(28) => 
                           s4_result_28_port, reg_ff(27) => s4_result_27_port, 
                           reg_ff(26) => s4_result_26_port, reg_ff(25) => 
                           s4_result_25_port, reg_ff(24) => s4_result_24_port, 
                           reg_ff(23) => s4_result_23_port, reg_ff(22) => 
                           s4_result_22_port, reg_ff(21) => s4_result_21_port, 
                           reg_ff(20) => s4_result_20_port, reg_ff(19) => 
                           s4_result_19_port, reg_ff(18) => s4_result_18_port, 
                           reg_ff(17) => s4_result_17_port, reg_ff(16) => 
                           s4_result_16_port, reg_ff(15) => s4_result_15_port, 
                           reg_ff(14) => s4_result_14_port, reg_ff(13) => 
                           s4_result_13_port, reg_ff(12) => s4_result_12_port, 
                           reg_ff(11) => s4_result_11_port, reg_ff(10) => 
                           s4_result_10_port, reg_ff(9) => s4_result_9_port, 
                           reg_ff(8) => s4_result_8_port, reg_ff(7) => 
                           s4_result_7_port, reg_ff(6) => s4_result_6_port, 
                           reg_ff(5) => s4_result_5_port, reg_ff(4) => 
                           s4_result_4_port, reg_ff(3) => s4_result_3_port, 
                           reg_ff(2) => s4_result_2_port, reg_ff(1) => 
                           s4_result_1_port, reg_ff(0) => s4_result_0_port, 
                           addr_c(4) => istr_val(25), addr_c(3) => istr_val(24)
                           , addr_c(2) => istr_val(23), addr_c(1) => 
                           istr_val(22), addr_c(0) => istr_val(21), addr_f(4) 
                           => s3_wr_addr_4_port, addr_f(3) => s3_wr_addr_3_port
                           , addr_f(2) => s3_wr_addr_2_port, addr_f(1) => 
                           s3_wr_addr_1_port, addr_f(0) => s3_wr_addr_0_port, 
                           addr_ff(4) => s4_wr_addr_4_port, addr_ff(3) => 
                           s4_wr_addr_3_port, addr_ff(2) => s4_wr_addr_2_port, 
                           addr_ff(1) => s4_wr_addr_1_port, addr_ff(0) => 
                           s4_wr_addr_0_port, valid_f => s2_a_f_j_en, valid_ff 
                           => s2_a_ff_j_en, dirty_f => cw(8), dirty_ff => 
                           X_Logic0_port, en => X_Logic1_port, output(31) => 
                           s2_jump_addr_reg_31_port, output(30) => 
                           s2_jump_addr_reg_30_port, output(29) => 
                           s2_jump_addr_reg_29_port, output(28) => 
                           s2_jump_addr_reg_28_port, output(27) => 
                           s2_jump_addr_reg_27_port, output(26) => 
                           s2_jump_addr_reg_26_port, output(25) => 
                           s2_jump_addr_reg_25_port, output(24) => 
                           s2_jump_addr_reg_24_port, output(23) => 
                           s2_jump_addr_reg_23_port, output(22) => 
                           s2_jump_addr_reg_22_port, output(21) => 
                           s2_jump_addr_reg_21_port, output(20) => 
                           s2_jump_addr_reg_20_port, output(19) => 
                           s2_jump_addr_reg_19_port, output(18) => 
                           s2_jump_addr_reg_18_port, output(17) => 
                           s2_jump_addr_reg_17_port, output(16) => 
                           s2_jump_addr_reg_16_port, output(15) => 
                           s2_jump_addr_reg_15_port, output(14) => 
                           s2_jump_addr_reg_14_port, output(13) => 
                           s2_jump_addr_reg_13_port, output(12) => 
                           s2_jump_addr_reg_12_port, output(11) => 
                           s2_jump_addr_reg_11_port, output(10) => 
                           s2_jump_addr_reg_10_port, output(9) => 
                           s2_jump_addr_reg_9_port, output(8) => 
                           s2_jump_addr_reg_8_port, output(7) => 
                           s2_jump_addr_reg_7_port, output(6) => 
                           s2_jump_addr_reg_6_port, output(5) => 
                           s2_jump_addr_reg_5_port, output(4) => 
                           s2_jump_addr_reg_4_port, output(3) => 
                           s2_jump_addr_reg_3_port, output(2) => 
                           s2_jump_addr_reg_2_port, output(1) => 
                           s2_jump_addr_reg_1_port, output(0) => 
                           s2_jump_addr_reg_0_port, match_dirty_f => sig_jral, 
                           match_dirty_ff => net1290);
   REG_A : Reg_DATA_SIZE32_11 port map( rst => rst, en => cw(6), clk => clk, 
                           din(31) => s2_a_31_port, din(30) => s2_a_30_port, 
                           din(29) => s2_a_29_port, din(28) => s2_a_28_port, 
                           din(27) => s2_a_27_port, din(26) => s2_a_26_port, 
                           din(25) => s2_a_25_port, din(24) => s2_a_24_port, 
                           din(23) => s2_a_23_port, din(22) => s2_a_22_port, 
                           din(21) => s2_a_21_port, din(20) => s2_a_20_port, 
                           din(19) => s2_a_19_port, din(18) => s2_a_18_port, 
                           din(17) => s2_a_17_port, din(16) => s2_a_16_port, 
                           din(15) => s2_a_15_port, din(14) => s2_a_14_port, 
                           din(13) => s2_a_13_port, din(12) => s2_a_12_port, 
                           din(11) => s2_a_11_port, din(10) => s2_a_10_port, 
                           din(9) => s2_a_9_port, din(8) => s2_a_8_port, din(7)
                           => s2_a_7_port, din(6) => s2_a_6_port, din(5) => 
                           s2_a_5_port, din(4) => s2_a_4_port, din(3) => 
                           s2_a_3_port, din(2) => s2_a_2_port, din(1) => 
                           s2_a_1_port, din(0) => s2_a_0_port, dout(31) => 
                           s3_a_31_port, dout(30) => s3_a_30_port, dout(29) => 
                           s3_a_29_port, dout(28) => s3_a_28_port, dout(27) => 
                           s3_a_27_port, dout(26) => s3_a_26_port, dout(25) => 
                           s3_a_25_port, dout(24) => s3_a_24_port, dout(23) => 
                           s3_a_23_port, dout(22) => s3_a_22_port, dout(21) => 
                           s3_a_21_port, dout(20) => s3_a_20_port, dout(19) => 
                           s3_a_19_port, dout(18) => s3_a_18_port, dout(17) => 
                           s3_a_17_port, dout(16) => s3_a_16_port, dout(15) => 
                           s3_a_15_port, dout(14) => s3_a_14_port, dout(13) => 
                           s3_a_13_port, dout(12) => s3_a_12_port, dout(11) => 
                           s3_a_11_port, dout(10) => s3_a_10_port, dout(9) => 
                           s3_a_9_port, dout(8) => s3_a_8_port, dout(7) => 
                           s3_a_7_port, dout(6) => s3_a_6_port, dout(5) => 
                           s3_a_5_port, dout(4) => s3_a_4_port, dout(3) => 
                           s3_a_3_port, dout(2) => s3_a_2_port, dout(1) => 
                           s3_a_1_port, dout(0) => s3_a_0_port);
   REG_B : Reg_DATA_SIZE32_10 port map( rst => rst, en => cw(6), clk => clk, 
                           din(31) => s2_b_31_port, din(30) => s2_b_30_port, 
                           din(29) => s2_b_29_port, din(28) => s2_b_28_port, 
                           din(27) => s2_b_27_port, din(26) => s2_b_26_port, 
                           din(25) => s2_b_25_port, din(24) => s2_b_24_port, 
                           din(23) => s2_b_23_port, din(22) => s2_b_22_port, 
                           din(21) => s2_b_21_port, din(20) => s2_b_20_port, 
                           din(19) => s2_b_19_port, din(18) => s2_b_18_port, 
                           din(17) => s2_b_17_port, din(16) => s2_b_16_port, 
                           din(15) => s2_b_15_port, din(14) => s2_b_14_port, 
                           din(13) => s2_b_13_port, din(12) => s2_b_12_port, 
                           din(11) => s2_b_11_port, din(10) => s2_b_10_port, 
                           din(9) => s2_b_9_port, din(8) => s2_b_8_port, din(7)
                           => s2_b_7_port, din(6) => s2_b_6_port, din(5) => 
                           s2_b_5_port, din(4) => s2_b_4_port, din(3) => 
                           s2_b_3_port, din(2) => s2_b_2_port, din(1) => 
                           s2_b_1_port, din(0) => s2_b_0_port, dout(31) => 
                           s3_b_31_port, dout(30) => s3_b_30_port, dout(29) => 
                           s3_b_29_port, dout(28) => s3_b_28_port, dout(27) => 
                           s3_b_27_port, dout(26) => s3_b_26_port, dout(25) => 
                           s3_b_25_port, dout(24) => s3_b_24_port, dout(23) => 
                           s3_b_23_port, dout(22) => s3_b_22_port, dout(21) => 
                           s3_b_21_port, dout(20) => s3_b_20_port, dout(19) => 
                           s3_b_19_port, dout(18) => s3_b_18_port, dout(17) => 
                           s3_b_17_port, dout(16) => s3_b_16_port, dout(15) => 
                           s3_b_15_port, dout(14) => s3_b_14_port, dout(13) => 
                           s3_b_13_port, dout(12) => s3_b_12_port, dout(11) => 
                           s3_b_11_port, dout(10) => s3_b_10_port, dout(9) => 
                           s3_b_9_port, dout(8) => s3_b_8_port, dout(7) => 
                           s3_b_7_port, dout(6) => s3_b_6_port, dout(5) => 
                           s3_b_5_port, dout(4) => s3_b_4_port, dout(3) => 
                           s3_b_3_port, dout(2) => s3_b_2_port, dout(1) => 
                           s3_b_1_port, dout(0) => s3_b_0_port);
   REG_I : Reg_DATA_SIZE32_9 port map( rst => rst, en => cw(6), clk => clk, 
                           din(31) => s2_imm_i_ext_31_port, din(30) => 
                           s2_imm_i_ext_30_port, din(29) => 
                           s2_imm_i_ext_29_port, din(28) => 
                           s2_imm_i_ext_28_port, din(27) => 
                           s2_imm_i_ext_27_port, din(26) => 
                           s2_imm_i_ext_26_port, din(25) => 
                           s2_imm_i_ext_25_port, din(24) => 
                           s2_imm_i_ext_24_port, din(23) => 
                           s2_imm_i_ext_23_port, din(22) => 
                           s2_imm_i_ext_22_port, din(21) => 
                           s2_imm_i_ext_21_port, din(20) => 
                           s2_imm_i_ext_20_port, din(19) => 
                           s2_imm_i_ext_19_port, din(18) => 
                           s2_imm_i_ext_18_port, din(17) => 
                           s2_imm_i_ext_17_port, din(16) => 
                           s2_imm_i_ext_16_port, din(15) => 
                           s2_imm_i_ext_15_port, din(14) => 
                           s2_imm_i_ext_14_port, din(13) => 
                           s2_imm_i_ext_13_port, din(12) => 
                           s2_imm_i_ext_12_port, din(11) => 
                           s2_imm_i_ext_11_port, din(10) => 
                           s2_imm_i_ext_10_port, din(9) => s2_imm_i_ext_9_port,
                           din(8) => s2_imm_i_ext_8_port, din(7) => 
                           s2_imm_i_ext_7_port, din(6) => s2_imm_i_ext_6_port, 
                           din(5) => s2_imm_i_ext_5_port, din(4) => 
                           s2_imm_i_ext_4_port, din(3) => s2_imm_i_ext_3_port, 
                           din(2) => s2_imm_i_ext_2_port, din(1) => 
                           s2_imm_i_ext_1_port, din(0) => s2_imm_i_ext_0_port, 
                           dout(31) => s3_imm_i_ext_31_port, dout(30) => 
                           s3_imm_i_ext_30_port, dout(29) => 
                           s3_imm_i_ext_29_port, dout(28) => 
                           s3_imm_i_ext_28_port, dout(27) => 
                           s3_imm_i_ext_27_port, dout(26) => 
                           s3_imm_i_ext_26_port, dout(25) => 
                           s3_imm_i_ext_25_port, dout(24) => 
                           s3_imm_i_ext_24_port, dout(23) => 
                           s3_imm_i_ext_23_port, dout(22) => 
                           s3_imm_i_ext_22_port, dout(21) => 
                           s3_imm_i_ext_21_port, dout(20) => 
                           s3_imm_i_ext_20_port, dout(19) => 
                           s3_imm_i_ext_19_port, dout(18) => 
                           s3_imm_i_ext_18_port, dout(17) => 
                           s3_imm_i_ext_17_port, dout(16) => 
                           s3_imm_i_ext_16_port, dout(15) => 
                           s3_imm_i_ext_15_port, dout(14) => 
                           s3_imm_i_ext_14_port, dout(13) => 
                           s3_imm_i_ext_13_port, dout(12) => 
                           s3_imm_i_ext_12_port, dout(11) => 
                           s3_imm_i_ext_11_port, dout(10) => 
                           s3_imm_i_ext_10_port, dout(9) => s3_imm_i_ext_9_port
                           , dout(8) => s3_imm_i_ext_8_port, dout(7) => 
                           s3_imm_i_ext_7_port, dout(6) => s3_imm_i_ext_6_port,
                           dout(5) => s3_imm_i_ext_5_port, dout(4) => 
                           s3_imm_i_ext_4_port, dout(3) => s3_imm_i_ext_3_port,
                           dout(2) => s3_imm_i_ext_2_port, dout(1) => 
                           s3_imm_i_ext_1_port, dout(0) => s3_imm_i_ext_0_port)
                           ;
   REG_WR2 : Reg_DATA_SIZE5_0 port map( rst => rst, en => cw(6), clk => clk, 
                           din(4) => s2_wr_addr_4_port, din(3) => 
                           s2_wr_addr_3_port, din(2) => s2_wr_addr_2_port, 
                           din(1) => s2_wr_addr_1_port, din(0) => 
                           s2_wr_addr_0_port, dout(4) => s3_wr_addr_4_port, 
                           dout(3) => s3_wr_addr_3_port, dout(2) => 
                           s3_wr_addr_2_port, dout(1) => s3_wr_addr_1_port, 
                           dout(0) => s3_wr_addr_0_port);
   REG_A_ADDR_2 : Reg_DATA_SIZE5_6 port map( rst => rst, en => cw(6), clk => 
                           clk, din(4) => istr_val(25), din(3) => istr_val(24),
                           din(2) => istr_val(23), din(1) => istr_val(22), 
                           din(0) => istr_val(21), dout(4) => 
                           s3_rd1_addr_4_port, dout(3) => s3_rd1_addr_3_port, 
                           dout(2) => s3_rd1_addr_2_port, dout(1) => 
                           s3_rd1_addr_1_port, dout(0) => s3_rd1_addr_0_port);
   REG_B_ADDR_2 : Reg_DATA_SIZE5_5 port map( rst => rst, en => cw(6), clk => 
                           clk, din(4) => istr_val(20), din(3) => istr_val(19),
                           din(2) => istr_val(18), din(1) => istr_val(17), 
                           din(0) => istr_val(16), dout(4) => 
                           s3_rd2_addr_4_port, dout(3) => s3_rd2_addr_3_port, 
                           dout(2) => s3_rd2_addr_2_port, dout(1) => 
                           s3_rd2_addr_1_port, dout(0) => s3_rd2_addr_0_port);
   REG_PC_NOT_SEL : Reg_DATA_SIZE32_8 port map( rst => rst, en => cw(6), clk =>
                           clk, din(31) => s2_pc_notsel_31_port, din(30) => 
                           s2_pc_notsel_30_port, din(29) => 
                           s2_pc_notsel_29_port, din(28) => 
                           s2_pc_notsel_28_port, din(27) => 
                           s2_pc_notsel_27_port, din(26) => 
                           s2_pc_notsel_26_port, din(25) => 
                           s2_pc_notsel_25_port, din(24) => 
                           s2_pc_notsel_24_port, din(23) => 
                           s2_pc_notsel_23_port, din(22) => 
                           s2_pc_notsel_22_port, din(21) => 
                           s2_pc_notsel_21_port, din(20) => 
                           s2_pc_notsel_20_port, din(19) => 
                           s2_pc_notsel_19_port, din(18) => 
                           s2_pc_notsel_18_port, din(17) => 
                           s2_pc_notsel_17_port, din(16) => 
                           s2_pc_notsel_16_port, din(15) => 
                           s2_pc_notsel_15_port, din(14) => 
                           s2_pc_notsel_14_port, din(13) => 
                           s2_pc_notsel_13_port, din(12) => 
                           s2_pc_notsel_12_port, din(11) => 
                           s2_pc_notsel_11_port, din(10) => 
                           s2_pc_notsel_10_port, din(9) => s2_pc_notsel_9_port,
                           din(8) => s2_pc_notsel_8_port, din(7) => 
                           s2_pc_notsel_7_port, din(6) => s2_pc_notsel_6_port, 
                           din(5) => s2_pc_notsel_5_port, din(4) => 
                           s2_pc_notsel_4_port, din(3) => s2_pc_notsel_3_port, 
                           din(2) => s2_pc_notsel_2_port, din(1) => 
                           s2_pc_notsel_1_port, din(0) => s2_pc_notsel_0_port, 
                           dout(31) => s3_pc_notsel_31_port, dout(30) => 
                           s3_pc_notsel_30_port, dout(29) => 
                           s3_pc_notsel_29_port, dout(28) => 
                           s3_pc_notsel_28_port, dout(27) => 
                           s3_pc_notsel_27_port, dout(26) => 
                           s3_pc_notsel_26_port, dout(25) => 
                           s3_pc_notsel_25_port, dout(24) => 
                           s3_pc_notsel_24_port, dout(23) => 
                           s3_pc_notsel_23_port, dout(22) => 
                           s3_pc_notsel_22_port, dout(21) => 
                           s3_pc_notsel_21_port, dout(20) => 
                           s3_pc_notsel_20_port, dout(19) => 
                           s3_pc_notsel_19_port, dout(18) => 
                           s3_pc_notsel_18_port, dout(17) => 
                           s3_pc_notsel_17_port, dout(16) => 
                           s3_pc_notsel_16_port, dout(15) => 
                           s3_pc_notsel_15_port, dout(14) => 
                           s3_pc_notsel_14_port, dout(13) => 
                           s3_pc_notsel_13_port, dout(12) => 
                           s3_pc_notsel_12_port, dout(11) => 
                           s3_pc_notsel_11_port, dout(10) => 
                           s3_pc_notsel_10_port, dout(9) => s3_pc_notsel_9_port
                           , dout(8) => s3_pc_notsel_8_port, dout(7) => 
                           s3_pc_notsel_7_port, dout(6) => s3_pc_notsel_6_port,
                           dout(5) => s3_pc_notsel_5_port, dout(4) => 
                           s3_pc_notsel_4_port, dout(3) => s3_pc_notsel_3_port,
                           dout(2) => s3_pc_notsel_2_port, dout(1) => 
                           s3_pc_notsel_1_port, dout(0) => s3_pc_notsel_0_port)
                           ;
   MUX_KEEP_A : Mux_DATA_SIZE32_5 port map( sel => s4_reg_b_wait, din0(31) => 
                           s3_a_31_port, din0(30) => s3_a_30_port, din0(29) => 
                           s3_a_29_port, din0(28) => s3_a_28_port, din0(27) => 
                           s3_a_27_port, din0(26) => s3_a_26_port, din0(25) => 
                           s3_a_25_port, din0(24) => s3_a_24_port, din0(23) => 
                           s3_a_23_port, din0(22) => s3_a_22_port, din0(21) => 
                           s3_a_21_port, din0(20) => s3_a_20_port, din0(19) => 
                           s3_a_19_port, din0(18) => s3_a_18_port, din0(17) => 
                           s3_a_17_port, din0(16) => s3_a_16_port, din0(15) => 
                           s3_a_15_port, din0(14) => s3_a_14_port, din0(13) => 
                           s3_a_13_port, din0(12) => s3_a_12_port, din0(11) => 
                           s3_a_11_port, din0(10) => s3_a_10_port, din0(9) => 
                           s3_a_9_port, din0(8) => s3_a_8_port, din0(7) => 
                           s3_a_7_port, din0(6) => s3_a_6_port, din0(5) => 
                           s3_a_5_port, din0(4) => s3_a_4_port, din0(3) => 
                           s3_a_3_port, din0(2) => s3_a_2_port, din0(1) => 
                           s3_a_1_port, din0(0) => s3_a_0_port, din1(31) => 
                           s4_a_31_port, din1(30) => s4_a_30_port, din1(29) => 
                           s4_a_29_port, din1(28) => s4_a_28_port, din1(27) => 
                           s4_a_27_port, din1(26) => s4_a_26_port, din1(25) => 
                           s4_a_25_port, din1(24) => s4_a_24_port, din1(23) => 
                           s4_a_23_port, din1(22) => s4_a_22_port, din1(21) => 
                           s4_a_21_port, din1(20) => s4_a_20_port, din1(19) => 
                           s4_a_19_port, din1(18) => s4_a_18_port, din1(17) => 
                           s4_a_17_port, din1(16) => s4_a_16_port, din1(15) => 
                           s4_a_15_port, din1(14) => s4_a_14_port, din1(13) => 
                           s4_a_13_port, din1(12) => s4_a_12_port, din1(11) => 
                           s4_a_11_port, din1(10) => s4_a_10_port, din1(9) => 
                           s4_a_9_port, din1(8) => s4_a_8_port, din1(7) => 
                           s4_a_7_port, din1(6) => s4_a_6_port, din1(5) => 
                           s4_a_5_port, din1(4) => s4_a_4_port, din1(3) => 
                           s4_a_3_port, din1(2) => s4_a_2_port, din1(1) => 
                           s4_a_1_port, din1(0) => s4_a_0_port, dout(31) => 
                           s3_a_keep_31_port, dout(30) => s3_a_keep_30_port, 
                           dout(29) => s3_a_keep_29_port, dout(28) => 
                           s3_a_keep_28_port, dout(27) => s3_a_keep_27_port, 
                           dout(26) => s3_a_keep_26_port, dout(25) => 
                           s3_a_keep_25_port, dout(24) => s3_a_keep_24_port, 
                           dout(23) => s3_a_keep_23_port, dout(22) => 
                           s3_a_keep_22_port, dout(21) => s3_a_keep_21_port, 
                           dout(20) => s3_a_keep_20_port, dout(19) => 
                           s3_a_keep_19_port, dout(18) => s3_a_keep_18_port, 
                           dout(17) => s3_a_keep_17_port, dout(16) => 
                           s3_a_keep_16_port, dout(15) => s3_a_keep_15_port, 
                           dout(14) => s3_a_keep_14_port, dout(13) => 
                           s3_a_keep_13_port, dout(12) => s3_a_keep_12_port, 
                           dout(11) => s3_a_keep_11_port, dout(10) => 
                           s3_a_keep_10_port, dout(9) => s3_a_keep_9_port, 
                           dout(8) => s3_a_keep_8_port, dout(7) => 
                           s3_a_keep_7_port, dout(6) => s3_a_keep_6_port, 
                           dout(5) => s3_a_keep_5_port, dout(4) => 
                           s3_a_keep_4_port, dout(3) => s3_a_keep_3_port, 
                           dout(2) => s3_a_keep_2_port, dout(1) => 
                           s3_a_keep_1_port, dout(0) => s3_a_keep_0_port);
   MUX_KEEP_B : Mux_DATA_SIZE32_4 port map( sel => s4_reg_a_wait, din0(31) => 
                           s3_b_31_port, din0(30) => s3_b_30_port, din0(29) => 
                           s3_b_29_port, din0(28) => s3_b_28_port, din0(27) => 
                           s3_b_27_port, din0(26) => s3_b_26_port, din0(25) => 
                           s3_b_25_port, din0(24) => s3_b_24_port, din0(23) => 
                           s3_b_23_port, din0(22) => s3_b_22_port, din0(21) => 
                           s3_b_21_port, din0(20) => s3_b_20_port, din0(19) => 
                           s3_b_19_port, din0(18) => s3_b_18_port, din0(17) => 
                           s3_b_17_port, din0(16) => s3_b_16_port, din0(15) => 
                           s3_b_15_port, din0(14) => s3_b_14_port, din0(13) => 
                           s3_b_13_port, din0(12) => s3_b_12_port, din0(11) => 
                           s3_b_11_port, din0(10) => s3_b_10_port, din0(9) => 
                           s3_b_9_port, din0(8) => s3_b_8_port, din0(7) => 
                           s3_b_7_port, din0(6) => s3_b_6_port, din0(5) => 
                           s3_b_5_port, din0(4) => s3_b_4_port, din0(3) => 
                           s3_b_3_port, din0(2) => s3_b_2_port, din0(1) => 
                           s3_b_1_port, din0(0) => s3_b_0_port, din1(31) => 
                           s4_b_31_port, din1(30) => s4_b_30_port, din1(29) => 
                           s4_b_29_port, din1(28) => s4_b_28_port, din1(27) => 
                           s4_b_27_port, din1(26) => s4_b_26_port, din1(25) => 
                           s4_b_25_port, din1(24) => s4_b_24_port, din1(23) => 
                           s4_b_23_port, din1(22) => s4_b_22_port, din1(21) => 
                           s4_b_21_port, din1(20) => s4_b_20_port, din1(19) => 
                           s4_b_19_port, din1(18) => s4_b_18_port, din1(17) => 
                           s4_b_17_port, din1(16) => s4_b_16_port, din1(15) => 
                           s4_b_15_port, din1(14) => s4_b_14_port, din1(13) => 
                           s4_b_13_port, din1(12) => s4_b_12_port, din1(11) => 
                           s4_b_11_port, din1(10) => s4_b_10_port, din1(9) => 
                           s4_b_9_port, din1(8) => s4_b_8_port, din1(7) => 
                           s4_b_7_port, din1(6) => s4_b_6_port, din1(5) => 
                           s4_b_5_port, din1(4) => s4_b_4_port, din1(3) => 
                           s4_b_3_port, din1(2) => s4_b_2_port, din1(1) => 
                           s4_b_1_port, din1(0) => s4_b_0_port, dout(31) => 
                           s3_b_keep_31_port, dout(30) => s3_b_keep_30_port, 
                           dout(29) => s3_b_keep_29_port, dout(28) => 
                           s3_b_keep_28_port, dout(27) => s3_b_keep_27_port, 
                           dout(26) => s3_b_keep_26_port, dout(25) => 
                           s3_b_keep_25_port, dout(24) => s3_b_keep_24_port, 
                           dout(23) => s3_b_keep_23_port, dout(22) => 
                           s3_b_keep_22_port, dout(21) => s3_b_keep_21_port, 
                           dout(20) => s3_b_keep_20_port, dout(19) => 
                           s3_b_keep_19_port, dout(18) => s3_b_keep_18_port, 
                           dout(17) => s3_b_keep_17_port, dout(16) => 
                           s3_b_keep_16_port, dout(15) => s3_b_keep_15_port, 
                           dout(14) => s3_b_keep_14_port, dout(13) => 
                           s3_b_keep_13_port, dout(12) => s3_b_keep_12_port, 
                           dout(11) => s3_b_keep_11_port, dout(10) => 
                           s3_b_keep_10_port, dout(9) => s3_b_keep_9_port, 
                           dout(8) => s3_b_keep_8_port, dout(7) => 
                           s3_b_keep_7_port, dout(6) => s3_b_keep_6_port, 
                           dout(5) => s3_b_keep_5_port, dout(4) => 
                           s3_b_keep_4_port, dout(3) => s3_b_keep_3_port, 
                           dout(2) => s3_b_keep_2_port, dout(1) => 
                           s3_b_keep_1_port, dout(0) => s3_b_keep_0_port);
   FWDMUX_A : FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_3 port map( reg_c(31) => 
                           s3_a_keep_31_port, reg_c(30) => s3_a_keep_30_port, 
                           reg_c(29) => s3_a_keep_29_port, reg_c(28) => 
                           s3_a_keep_28_port, reg_c(27) => s3_a_keep_27_port, 
                           reg_c(26) => s3_a_keep_26_port, reg_c(25) => 
                           s3_a_keep_25_port, reg_c(24) => s3_a_keep_24_port, 
                           reg_c(23) => s3_a_keep_23_port, reg_c(22) => 
                           s3_a_keep_22_port, reg_c(21) => s3_a_keep_21_port, 
                           reg_c(20) => s3_a_keep_20_port, reg_c(19) => 
                           s3_a_keep_19_port, reg_c(18) => s3_a_keep_18_port, 
                           reg_c(17) => s3_a_keep_17_port, reg_c(16) => 
                           s3_a_keep_16_port, reg_c(15) => s3_a_keep_15_port, 
                           reg_c(14) => s3_a_keep_14_port, reg_c(13) => 
                           s3_a_keep_13_port, reg_c(12) => s3_a_keep_12_port, 
                           reg_c(11) => s3_a_keep_11_port, reg_c(10) => 
                           s3_a_keep_10_port, reg_c(9) => s3_a_keep_9_port, 
                           reg_c(8) => s3_a_keep_8_port, reg_c(7) => 
                           s3_a_keep_7_port, reg_c(6) => s3_a_keep_6_port, 
                           reg_c(5) => s3_a_keep_5_port, reg_c(4) => 
                           s3_a_keep_4_port, reg_c(3) => s3_a_keep_3_port, 
                           reg_c(2) => s3_a_keep_2_port, reg_c(1) => 
                           s3_a_keep_1_port, reg_c(0) => s3_a_keep_0_port, 
                           reg_f(31) => data_addr_31_port, reg_f(30) => 
                           data_addr_30_port, reg_f(29) => data_addr_29_port, 
                           reg_f(28) => data_addr_28_port, reg_f(27) => 
                           data_addr_27_port, reg_f(26) => data_addr_26_port, 
                           reg_f(25) => data_addr_25_port, reg_f(24) => 
                           data_addr_24_port, reg_f(23) => data_addr_23_port, 
                           reg_f(22) => data_addr_22_port, reg_f(21) => 
                           data_addr_21_port, reg_f(20) => data_addr_20_port, 
                           reg_f(19) => data_addr_19_port, reg_f(18) => 
                           data_addr_18_port, reg_f(17) => data_addr_17_port, 
                           reg_f(16) => data_addr_16_port, reg_f(15) => 
                           data_addr_15_port, reg_f(14) => data_addr_14_port, 
                           reg_f(13) => data_addr_13_port, reg_f(12) => 
                           data_addr_12_port, reg_f(11) => data_addr_11_port, 
                           reg_f(10) => data_addr_10_port, reg_f(9) => 
                           data_addr_9_port, reg_f(8) => data_addr_8_port, 
                           reg_f(7) => data_addr_7_port, reg_f(6) => 
                           data_addr_6_port, reg_f(5) => data_addr_5_port, 
                           reg_f(4) => data_addr_4_port, reg_f(3) => 
                           data_addr_3_port, reg_f(2) => data_addr_2_port, 
                           reg_f(1) => data_addr_1_port, reg_f(0) => 
                           data_addr_0_port, reg_ff(31) => s5_result_31_port, 
                           reg_ff(30) => s5_result_30_port, reg_ff(29) => 
                           s5_result_29_port, reg_ff(28) => s5_result_28_port, 
                           reg_ff(27) => s5_result_27_port, reg_ff(26) => 
                           s5_result_26_port, reg_ff(25) => s5_result_25_port, 
                           reg_ff(24) => s5_result_24_port, reg_ff(23) => 
                           s5_result_23_port, reg_ff(22) => s5_result_22_port, 
                           reg_ff(21) => s5_result_21_port, reg_ff(20) => 
                           s5_result_20_port, reg_ff(19) => s5_result_19_port, 
                           reg_ff(18) => s5_result_18_port, reg_ff(17) => 
                           s5_result_17_port, reg_ff(16) => s5_result_16_port, 
                           reg_ff(15) => s5_result_15_port, reg_ff(14) => 
                           s5_result_14_port, reg_ff(13) => s5_result_13_port, 
                           reg_ff(12) => s5_result_12_port, reg_ff(11) => 
                           s5_result_11_port, reg_ff(10) => s5_result_10_port, 
                           reg_ff(9) => s5_result_9_port, reg_ff(8) => 
                           s5_result_8_port, reg_ff(7) => s5_result_7_port, 
                           reg_ff(6) => s5_result_6_port, reg_ff(5) => 
                           s5_result_5_port, reg_ff(4) => s5_result_4_port, 
                           reg_ff(3) => s5_result_3_port, reg_ff(2) => 
                           s5_result_2_port, reg_ff(1) => s5_result_1_port, 
                           reg_ff(0) => s5_result_0_port, addr_c(4) => 
                           s3_rd1_addr_4_port, addr_c(3) => s3_rd1_addr_3_port,
                           addr_c(2) => s3_rd1_addr_2_port, addr_c(1) => 
                           s3_rd1_addr_1_port, addr_c(0) => s3_rd1_addr_0_port,
                           addr_f(4) => s4_wr_addr_4_port, addr_f(3) => 
                           s4_wr_addr_3_port, addr_f(2) => s4_wr_addr_2_port, 
                           addr_f(1) => s4_wr_addr_1_port, addr_f(0) => 
                           s4_wr_addr_0_port, addr_ff(4) => s5_wr_addr_4_port, 
                           addr_ff(3) => s5_wr_addr_3_port, addr_ff(2) => 
                           s5_wr_addr_2_port, addr_ff(1) => s5_wr_addr_1_port, 
                           addr_ff(0) => s5_wr_addr_0_port, valid_f => 
                           s3_a_sel_f_en, valid_ff => s3_a_sel_ff_en, dirty_f 
                           => cw(16), dirty_ff => X_Logic0_port, en => 
                           X_Logic1_port, output(31) => s3_a_sel_31_port, 
                           output(30) => s3_a_sel_30_port, output(29) => 
                           s3_a_sel_29_port, output(28) => s3_a_sel_28_port, 
                           output(27) => s3_a_sel_27_port, output(26) => 
                           s3_a_sel_26_port, output(25) => s3_a_sel_25_port, 
                           output(24) => s3_a_sel_24_port, output(23) => 
                           s3_a_sel_23_port, output(22) => s3_a_sel_22_port, 
                           output(21) => s3_a_sel_21_port, output(20) => 
                           s3_a_sel_20_port, output(19) => s3_a_sel_19_port, 
                           output(18) => s3_a_sel_18_port, output(17) => 
                           s3_a_sel_17_port, output(16) => s3_a_sel_16_port, 
                           output(15) => s3_a_sel_15_port, output(14) => 
                           s3_a_sel_14_port, output(13) => s3_a_sel_13_port, 
                           output(12) => s3_a_sel_12_port, output(11) => 
                           s3_a_sel_11_port, output(10) => s3_a_sel_10_port, 
                           output(9) => s3_a_sel_9_port, output(8) => 
                           s3_a_sel_8_port, output(7) => s3_a_sel_7_port, 
                           output(6) => s3_a_sel_6_port, output(5) => 
                           s3_a_sel_5_port, output(4) => s3_a_sel_4_port, 
                           output(3) => s3_a_sel_3_port, output(2) => 
                           s3_a_sel_2_port, output(1) => s3_a_sel_1_port, 
                           output(0) => s3_a_sel_0_port, match_dirty_f => 
                           s3_reg_a_wait, match_dirty_ff => net1288);
   FWDMUX_B : FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_2 port map( reg_c(31) => 
                           s3_b_keep_31_port, reg_c(30) => s3_b_keep_30_port, 
                           reg_c(29) => s3_b_keep_29_port, reg_c(28) => 
                           s3_b_keep_28_port, reg_c(27) => s3_b_keep_27_port, 
                           reg_c(26) => s3_b_keep_26_port, reg_c(25) => 
                           s3_b_keep_25_port, reg_c(24) => s3_b_keep_24_port, 
                           reg_c(23) => s3_b_keep_23_port, reg_c(22) => 
                           s3_b_keep_22_port, reg_c(21) => s3_b_keep_21_port, 
                           reg_c(20) => s3_b_keep_20_port, reg_c(19) => 
                           s3_b_keep_19_port, reg_c(18) => s3_b_keep_18_port, 
                           reg_c(17) => s3_b_keep_17_port, reg_c(16) => 
                           s3_b_keep_16_port, reg_c(15) => s3_b_keep_15_port, 
                           reg_c(14) => s3_b_keep_14_port, reg_c(13) => 
                           s3_b_keep_13_port, reg_c(12) => s3_b_keep_12_port, 
                           reg_c(11) => s3_b_keep_11_port, reg_c(10) => 
                           s3_b_keep_10_port, reg_c(9) => s3_b_keep_9_port, 
                           reg_c(8) => s3_b_keep_8_port, reg_c(7) => 
                           s3_b_keep_7_port, reg_c(6) => s3_b_keep_6_port, 
                           reg_c(5) => s3_b_keep_5_port, reg_c(4) => 
                           s3_b_keep_4_port, reg_c(3) => s3_b_keep_3_port, 
                           reg_c(2) => s3_b_keep_2_port, reg_c(1) => 
                           s3_b_keep_1_port, reg_c(0) => s3_b_keep_0_port, 
                           reg_f(31) => data_addr_31_port, reg_f(30) => 
                           data_addr_30_port, reg_f(29) => data_addr_29_port, 
                           reg_f(28) => data_addr_28_port, reg_f(27) => 
                           data_addr_27_port, reg_f(26) => data_addr_26_port, 
                           reg_f(25) => data_addr_25_port, reg_f(24) => 
                           data_addr_24_port, reg_f(23) => data_addr_23_port, 
                           reg_f(22) => data_addr_22_port, reg_f(21) => 
                           data_addr_21_port, reg_f(20) => data_addr_20_port, 
                           reg_f(19) => data_addr_19_port, reg_f(18) => 
                           data_addr_18_port, reg_f(17) => data_addr_17_port, 
                           reg_f(16) => data_addr_16_port, reg_f(15) => 
                           data_addr_15_port, reg_f(14) => data_addr_14_port, 
                           reg_f(13) => data_addr_13_port, reg_f(12) => 
                           data_addr_12_port, reg_f(11) => data_addr_11_port, 
                           reg_f(10) => data_addr_10_port, reg_f(9) => 
                           data_addr_9_port, reg_f(8) => data_addr_8_port, 
                           reg_f(7) => data_addr_7_port, reg_f(6) => 
                           data_addr_6_port, reg_f(5) => data_addr_5_port, 
                           reg_f(4) => data_addr_4_port, reg_f(3) => 
                           data_addr_3_port, reg_f(2) => data_addr_2_port, 
                           reg_f(1) => data_addr_1_port, reg_f(0) => 
                           data_addr_0_port, reg_ff(31) => s5_result_31_port, 
                           reg_ff(30) => s5_result_30_port, reg_ff(29) => 
                           s5_result_29_port, reg_ff(28) => s5_result_28_port, 
                           reg_ff(27) => s5_result_27_port, reg_ff(26) => 
                           s5_result_26_port, reg_ff(25) => s5_result_25_port, 
                           reg_ff(24) => s5_result_24_port, reg_ff(23) => 
                           s5_result_23_port, reg_ff(22) => s5_result_22_port, 
                           reg_ff(21) => s5_result_21_port, reg_ff(20) => 
                           s5_result_20_port, reg_ff(19) => s5_result_19_port, 
                           reg_ff(18) => s5_result_18_port, reg_ff(17) => 
                           s5_result_17_port, reg_ff(16) => s5_result_16_port, 
                           reg_ff(15) => s5_result_15_port, reg_ff(14) => 
                           s5_result_14_port, reg_ff(13) => s5_result_13_port, 
                           reg_ff(12) => s5_result_12_port, reg_ff(11) => 
                           s5_result_11_port, reg_ff(10) => s5_result_10_port, 
                           reg_ff(9) => s5_result_9_port, reg_ff(8) => 
                           s5_result_8_port, reg_ff(7) => s5_result_7_port, 
                           reg_ff(6) => s5_result_6_port, reg_ff(5) => 
                           s5_result_5_port, reg_ff(4) => s5_result_4_port, 
                           reg_ff(3) => s5_result_3_port, reg_ff(2) => 
                           s5_result_2_port, reg_ff(1) => s5_result_1_port, 
                           reg_ff(0) => s5_result_0_port, addr_c(4) => 
                           s3_rd2_addr_4_port, addr_c(3) => s3_rd2_addr_3_port,
                           addr_c(2) => s3_rd2_addr_2_port, addr_c(1) => 
                           s3_rd2_addr_1_port, addr_c(0) => s3_rd2_addr_0_port,
                           addr_f(4) => s4_wr_addr_4_port, addr_f(3) => 
                           s4_wr_addr_3_port, addr_f(2) => s4_wr_addr_2_port, 
                           addr_f(1) => s4_wr_addr_1_port, addr_f(0) => 
                           s4_wr_addr_0_port, addr_ff(4) => s5_wr_addr_4_port, 
                           addr_ff(3) => s5_wr_addr_3_port, addr_ff(2) => 
                           s5_wr_addr_2_port, addr_ff(1) => s5_wr_addr_1_port, 
                           addr_ff(0) => s5_wr_addr_0_port, valid_f => 
                           s3_b_sel_f_en, valid_ff => s3_b_sel_ff_en, dirty_f 
                           => cw(16), dirty_ff => X_Logic0_port, en => 
                           X_Logic1_port, output(31) => s3_b_fwd_31_port, 
                           output(30) => s3_b_fwd_30_port, output(29) => 
                           s3_b_fwd_29_port, output(28) => s3_b_fwd_28_port, 
                           output(27) => s3_b_fwd_27_port, output(26) => 
                           s3_b_fwd_26_port, output(25) => s3_b_fwd_25_port, 
                           output(24) => s3_b_fwd_24_port, output(23) => 
                           s3_b_fwd_23_port, output(22) => s3_b_fwd_22_port, 
                           output(21) => s3_b_fwd_21_port, output(20) => 
                           s3_b_fwd_20_port, output(19) => s3_b_fwd_19_port, 
                           output(18) => s3_b_fwd_18_port, output(17) => 
                           s3_b_fwd_17_port, output(16) => s3_b_fwd_16_port, 
                           output(15) => s3_b_fwd_15_port, output(14) => 
                           s3_b_fwd_14_port, output(13) => s3_b_fwd_13_port, 
                           output(12) => s3_b_fwd_12_port, output(11) => 
                           s3_b_fwd_11_port, output(10) => s3_b_fwd_10_port, 
                           output(9) => s3_b_fwd_9_port, output(8) => 
                           s3_b_fwd_8_port, output(7) => s3_b_fwd_7_port, 
                           output(6) => s3_b_fwd_6_port, output(5) => 
                           s3_b_fwd_5_port, output(4) => s3_b_fwd_4_port, 
                           output(3) => s3_b_fwd_3_port, output(2) => 
                           s3_b_fwd_2_port, output(1) => s3_b_fwd_1_port, 
                           output(0) => s3_b_fwd_0_port, match_dirty_f => 
                           s3_reg_b_wait, match_dirty_ff => net1287);
   MUXB : Mux_DATA_SIZE32_3 port map( sel => cw(7), din0(31) => 
                           s3_b_fwd_31_port, din0(30) => s3_b_fwd_30_port, 
                           din0(29) => s3_b_fwd_29_port, din0(28) => 
                           s3_b_fwd_28_port, din0(27) => s3_b_fwd_27_port, 
                           din0(26) => s3_b_fwd_26_port, din0(25) => 
                           s3_b_fwd_25_port, din0(24) => s3_b_fwd_24_port, 
                           din0(23) => s3_b_fwd_23_port, din0(22) => 
                           s3_b_fwd_22_port, din0(21) => s3_b_fwd_21_port, 
                           din0(20) => s3_b_fwd_20_port, din0(19) => 
                           s3_b_fwd_19_port, din0(18) => s3_b_fwd_18_port, 
                           din0(17) => s3_b_fwd_17_port, din0(16) => 
                           s3_b_fwd_16_port, din0(15) => s3_b_fwd_15_port, 
                           din0(14) => s3_b_fwd_14_port, din0(13) => 
                           s3_b_fwd_13_port, din0(12) => s3_b_fwd_12_port, 
                           din0(11) => s3_b_fwd_11_port, din0(10) => 
                           s3_b_fwd_10_port, din0(9) => s3_b_fwd_9_port, 
                           din0(8) => s3_b_fwd_8_port, din0(7) => 
                           s3_b_fwd_7_port, din0(6) => s3_b_fwd_6_port, din0(5)
                           => s3_b_fwd_5_port, din0(4) => s3_b_fwd_4_port, 
                           din0(3) => s3_b_fwd_3_port, din0(2) => 
                           s3_b_fwd_2_port, din0(1) => s3_b_fwd_1_port, din0(0)
                           => s3_b_fwd_0_port, din1(31) => s3_imm_i_ext_31_port
                           , din1(30) => s3_imm_i_ext_30_port, din1(29) => 
                           s3_imm_i_ext_29_port, din1(28) => 
                           s3_imm_i_ext_28_port, din1(27) => 
                           s3_imm_i_ext_27_port, din1(26) => 
                           s3_imm_i_ext_26_port, din1(25) => 
                           s3_imm_i_ext_25_port, din1(24) => 
                           s3_imm_i_ext_24_port, din1(23) => 
                           s3_imm_i_ext_23_port, din1(22) => 
                           s3_imm_i_ext_22_port, din1(21) => 
                           s3_imm_i_ext_21_port, din1(20) => 
                           s3_imm_i_ext_20_port, din1(19) => 
                           s3_imm_i_ext_19_port, din1(18) => 
                           s3_imm_i_ext_18_port, din1(17) => 
                           s3_imm_i_ext_17_port, din1(16) => 
                           s3_imm_i_ext_16_port, din1(15) => 
                           s3_imm_i_ext_15_port, din1(14) => 
                           s3_imm_i_ext_14_port, din1(13) => 
                           s3_imm_i_ext_13_port, din1(12) => 
                           s3_imm_i_ext_12_port, din1(11) => 
                           s3_imm_i_ext_11_port, din1(10) => 
                           s3_imm_i_ext_10_port, din1(9) => s3_imm_i_ext_9_port
                           , din1(8) => s3_imm_i_ext_8_port, din1(7) => 
                           s3_imm_i_ext_7_port, din1(6) => s3_imm_i_ext_6_port,
                           din1(5) => s3_imm_i_ext_5_port, din1(4) => 
                           s3_imm_i_ext_4_port, din1(3) => s3_imm_i_ext_3_port,
                           din1(2) => s3_imm_i_ext_2_port, din1(1) => 
                           s3_imm_i_ext_1_port, din1(0) => s3_imm_i_ext_0_port,
                           dout(31) => s3_b_sel_31_port, dout(30) => 
                           s3_b_sel_30_port, dout(29) => s3_b_sel_29_port, 
                           dout(28) => s3_b_sel_28_port, dout(27) => 
                           s3_b_sel_27_port, dout(26) => s3_b_sel_26_port, 
                           dout(25) => s3_b_sel_25_port, dout(24) => 
                           s3_b_sel_24_port, dout(23) => s3_b_sel_23_port, 
                           dout(22) => s3_b_sel_22_port, dout(21) => 
                           s3_b_sel_21_port, dout(20) => s3_b_sel_20_port, 
                           dout(19) => s3_b_sel_19_port, dout(18) => 
                           s3_b_sel_18_port, dout(17) => s3_b_sel_17_port, 
                           dout(16) => s3_b_sel_16_port, dout(15) => 
                           s3_b_sel_15_port, dout(14) => s3_b_sel_14_port, 
                           dout(13) => s3_b_sel_13_port, dout(12) => 
                           s3_b_sel_12_port, dout(11) => s3_b_sel_11_port, 
                           dout(10) => s3_b_sel_10_port, dout(9) => 
                           s3_b_sel_9_port, dout(8) => s3_b_sel_8_port, dout(7)
                           => s3_b_sel_7_port, dout(6) => s3_b_sel_6_port, 
                           dout(5) => s3_b_sel_5_port, dout(4) => 
                           s3_b_sel_4_port, dout(3) => s3_b_sel_3_port, dout(2)
                           => s3_b_sel_2_port, dout(1) => s3_b_sel_1_port, 
                           dout(0) => s3_b_sel_0_port);
   ALU0 : Alu_DATA_SIZE32 port map( f(4) => calu(4), f(3) => calu(3), f(2) => 
                           calu(2), f(1) => calu(1), f(0) => calu(0), a(31) => 
                           s3_a_sel_31_port, a(30) => s3_a_sel_30_port, a(29) 
                           => s3_a_sel_29_port, a(28) => s3_a_sel_28_port, 
                           a(27) => s3_a_sel_27_port, a(26) => s3_a_sel_26_port
                           , a(25) => s3_a_sel_25_port, a(24) => 
                           s3_a_sel_24_port, a(23) => s3_a_sel_23_port, a(22) 
                           => s3_a_sel_22_port, a(21) => s3_a_sel_21_port, 
                           a(20) => s3_a_sel_20_port, a(19) => s3_a_sel_19_port
                           , a(18) => s3_a_sel_18_port, a(17) => 
                           s3_a_sel_17_port, a(16) => s3_a_sel_16_port, a(15) 
                           => s3_a_sel_15_port, a(14) => s3_a_sel_14_port, 
                           a(13) => s3_a_sel_13_port, a(12) => s3_a_sel_12_port
                           , a(11) => s3_a_sel_11_port, a(10) => 
                           s3_a_sel_10_port, a(9) => s3_a_sel_9_port, a(8) => 
                           s3_a_sel_8_port, a(7) => s3_a_sel_7_port, a(6) => 
                           s3_a_sel_6_port, a(5) => s3_a_sel_5_port, a(4) => 
                           s3_a_sel_4_port, a(3) => s3_a_sel_3_port, a(2) => 
                           s3_a_sel_2_port, a(1) => s3_a_sel_1_port, a(0) => 
                           s3_a_sel_0_port, b(31) => s3_b_sel_31_port, b(30) =>
                           s3_b_sel_30_port, b(29) => s3_b_sel_29_port, b(28) 
                           => s3_b_sel_28_port, b(27) => s3_b_sel_27_port, 
                           b(26) => s3_b_sel_26_port, b(25) => s3_b_sel_25_port
                           , b(24) => s3_b_sel_24_port, b(23) => 
                           s3_b_sel_23_port, b(22) => s3_b_sel_22_port, b(21) 
                           => s3_b_sel_21_port, b(20) => s3_b_sel_20_port, 
                           b(19) => s3_b_sel_19_port, b(18) => s3_b_sel_18_port
                           , b(17) => s3_b_sel_17_port, b(16) => 
                           s3_b_sel_16_port, b(15) => s3_b_sel_15_port, b(14) 
                           => s3_b_sel_14_port, b(13) => s3_b_sel_13_port, 
                           b(12) => s3_b_sel_12_port, b(11) => s3_b_sel_11_port
                           , b(10) => s3_b_sel_10_port, b(9) => s3_b_sel_9_port
                           , b(8) => s3_b_sel_8_port, b(7) => s3_b_sel_7_port, 
                           b(6) => s3_b_sel_6_port, b(5) => s3_b_sel_5_port, 
                           b(4) => s3_b_sel_4_port, b(3) => s3_b_sel_3_port, 
                           b(2) => s3_b_sel_2_port, b(1) => s3_b_sel_1_port, 
                           b(0) => s3_b_sel_0_port, o(31) => s3_alu_out_31_port
                           , o(30) => s3_alu_out_30_port, o(29) => 
                           s3_alu_out_29_port, o(28) => s3_alu_out_28_port, 
                           o(27) => s3_alu_out_27_port, o(26) => 
                           s3_alu_out_26_port, o(25) => s3_alu_out_25_port, 
                           o(24) => s3_alu_out_24_port, o(23) => 
                           s3_alu_out_23_port, o(22) => s3_alu_out_22_port, 
                           o(21) => s3_alu_out_21_port, o(20) => 
                           s3_alu_out_20_port, o(19) => s3_alu_out_19_port, 
                           o(18) => s3_alu_out_18_port, o(17) => 
                           s3_alu_out_17_port, o(16) => s3_alu_out_16_port, 
                           o(15) => s3_alu_out_15_port, o(14) => 
                           s3_alu_out_14_port, o(13) => s3_alu_out_13_port, 
                           o(12) => s3_alu_out_12_port, o(11) => 
                           s3_alu_out_11_port, o(10) => s3_alu_out_10_port, 
                           o(9) => s3_alu_out_9_port, o(8) => s3_alu_out_8_port
                           , o(7) => s3_alu_out_7_port, o(6) => 
                           s3_alu_out_6_port, o(5) => s3_alu_out_5_port, o(4) 
                           => s3_alu_out_4_port, o(3) => s3_alu_out_3_port, 
                           o(2) => s3_alu_out_2_port, o(1) => s3_alu_out_1_port
                           , o(0) => s3_alu_out_0_port);
   MUL0 : Mul_DATA_SIZE16_STAGE10 port map( rst => rst, clk => clk, en => 
                           sig_mul_port, lock => sig_ral_port, sign => 
                           s3_mul_sign, a(15) => s3_a_sel_15_port, a(14) => 
                           s3_a_sel_14_port, a(13) => s3_a_sel_13_port, a(12) 
                           => s3_a_sel_12_port, a(11) => s3_a_sel_11_port, 
                           a(10) => s3_a_sel_10_port, a(9) => s3_a_sel_9_port, 
                           a(8) => s3_a_sel_8_port, a(7) => s3_a_sel_7_port, 
                           a(6) => s3_a_sel_6_port, a(5) => s3_a_sel_5_port, 
                           a(4) => s3_a_sel_4_port, a(3) => s3_a_sel_3_port, 
                           a(2) => s3_a_sel_2_port, a(1) => s3_a_sel_1_port, 
                           a(0) => s3_a_sel_0_port, b(15) => s3_b_sel_15_port, 
                           b(14) => s3_b_sel_14_port, b(13) => s3_b_sel_13_port
                           , b(12) => s3_b_sel_12_port, b(11) => 
                           s3_b_sel_11_port, b(10) => s3_b_sel_10_port, b(9) =>
                           s3_b_sel_9_port, b(8) => s3_b_sel_8_port, b(7) => 
                           s3_b_sel_7_port, b(6) => s3_b_sel_6_port, b(5) => 
                           s3_b_sel_5_port, b(4) => s3_b_sel_4_port, b(3) => 
                           s3_b_sel_3_port, b(2) => s3_b_sel_2_port, b(1) => 
                           s3_b_sel_1_port, b(0) => s3_b_sel_0_port, o(31) => 
                           s3_mul_out_31_port, o(30) => s3_mul_out_30_port, 
                           o(29) => s3_mul_out_29_port, o(28) => 
                           s3_mul_out_28_port, o(27) => s3_mul_out_27_port, 
                           o(26) => s3_mul_out_26_port, o(25) => 
                           s3_mul_out_25_port, o(24) => s3_mul_out_24_port, 
                           o(23) => s3_mul_out_23_port, o(22) => 
                           s3_mul_out_22_port, o(21) => s3_mul_out_21_port, 
                           o(20) => s3_mul_out_20_port, o(19) => 
                           s3_mul_out_19_port, o(18) => s3_mul_out_18_port, 
                           o(17) => s3_mul_out_17_port, o(16) => 
                           s3_mul_out_16_port, o(15) => s3_mul_out_15_port, 
                           o(14) => s3_mul_out_14_port, o(13) => 
                           s3_mul_out_13_port, o(12) => s3_mul_out_12_port, 
                           o(11) => s3_mul_out_11_port, o(10) => 
                           s3_mul_out_10_port, o(9) => s3_mul_out_9_port, o(8) 
                           => s3_mul_out_8_port, o(7) => s3_mul_out_7_port, 
                           o(6) => s3_mul_out_6_port, o(5) => s3_mul_out_5_port
                           , o(4) => s3_mul_out_4_port, o(3) => 
                           s3_mul_out_3_port, o(2) => s3_mul_out_2_port, o(1) 
                           => s3_mul_out_1_port, o(0) => s3_mul_out_0_port);
   DIV0 : Div_DATA_SIZE32_DIV_STAGE34_SQRT_STAGE18 port map( rst => rst, clk =>
                           clk, en => s3_exe_sel_1_port, lock => sig_ral_port, 
                           sign => s3_div_sign, func => sig_sqrt_port, a(31) =>
                           s3_a_sel_31_port, a(30) => s3_a_sel_30_port, a(29) 
                           => s3_a_sel_29_port, a(28) => s3_a_sel_28_port, 
                           a(27) => s3_a_sel_27_port, a(26) => s3_a_sel_26_port
                           , a(25) => s3_a_sel_25_port, a(24) => 
                           s3_a_sel_24_port, a(23) => s3_a_sel_23_port, a(22) 
                           => s3_a_sel_22_port, a(21) => s3_a_sel_21_port, 
                           a(20) => s3_a_sel_20_port, a(19) => s3_a_sel_19_port
                           , a(18) => s3_a_sel_18_port, a(17) => 
                           s3_a_sel_17_port, a(16) => s3_a_sel_16_port, a(15) 
                           => s3_a_sel_15_port, a(14) => s3_a_sel_14_port, 
                           a(13) => s3_a_sel_13_port, a(12) => s3_a_sel_12_port
                           , a(11) => s3_a_sel_11_port, a(10) => 
                           s3_a_sel_10_port, a(9) => s3_a_sel_9_port, a(8) => 
                           s3_a_sel_8_port, a(7) => s3_a_sel_7_port, a(6) => 
                           s3_a_sel_6_port, a(5) => s3_a_sel_5_port, a(4) => 
                           s3_a_sel_4_port, a(3) => s3_a_sel_3_port, a(2) => 
                           s3_a_sel_2_port, a(1) => s3_a_sel_1_port, a(0) => 
                           s3_a_sel_0_port, b(31) => s3_b_sel_31_port, b(30) =>
                           s3_b_sel_30_port, b(29) => s3_b_sel_29_port, b(28) 
                           => s3_b_sel_28_port, b(27) => s3_b_sel_27_port, 
                           b(26) => s3_b_sel_26_port, b(25) => s3_b_sel_25_port
                           , b(24) => s3_b_sel_24_port, b(23) => 
                           s3_b_sel_23_port, b(22) => s3_b_sel_22_port, b(21) 
                           => s3_b_sel_21_port, b(20) => s3_b_sel_20_port, 
                           b(19) => s3_b_sel_19_port, b(18) => s3_b_sel_18_port
                           , b(17) => s3_b_sel_17_port, b(16) => 
                           s3_b_sel_16_port, b(15) => s3_b_sel_15_port, b(14) 
                           => s3_b_sel_14_port, b(13) => s3_b_sel_13_port, 
                           b(12) => s3_b_sel_12_port, b(11) => s3_b_sel_11_port
                           , b(10) => s3_b_sel_10_port, b(9) => s3_b_sel_9_port
                           , b(8) => s3_b_sel_8_port, b(7) => s3_b_sel_7_port, 
                           b(6) => s3_b_sel_6_port, b(5) => s3_b_sel_5_port, 
                           b(4) => s3_b_sel_4_port, b(3) => s3_b_sel_3_port, 
                           b(2) => s3_b_sel_2_port, b(1) => s3_b_sel_1_port, 
                           b(0) => s3_b_sel_0_port, o(31) => s3_div_out_31_port
                           , o(30) => s3_div_out_30_port, o(29) => 
                           s3_div_out_29_port, o(28) => s3_div_out_28_port, 
                           o(27) => s3_div_out_27_port, o(26) => 
                           s3_div_out_26_port, o(25) => s3_div_out_25_port, 
                           o(24) => s3_div_out_24_port, o(23) => 
                           s3_div_out_23_port, o(22) => s3_div_out_22_port, 
                           o(21) => s3_div_out_21_port, o(20) => 
                           s3_div_out_20_port, o(19) => s3_div_out_19_port, 
                           o(18) => s3_div_out_18_port, o(17) => 
                           s3_div_out_17_port, o(16) => s3_div_out_16_port, 
                           o(15) => s3_div_out_15_port, o(14) => 
                           s3_div_out_14_port, o(13) => s3_div_out_13_port, 
                           o(12) => s3_div_out_12_port, o(11) => 
                           s3_div_out_11_port, o(10) => s3_div_out_10_port, 
                           o(9) => s3_div_out_9_port, o(8) => s3_div_out_8_port
                           , o(7) => s3_div_out_7_port, o(6) => 
                           s3_div_out_6_port, o(5) => s3_div_out_5_port, o(4) 
                           => s3_div_out_4_port, o(3) => s3_div_out_3_port, 
                           o(2) => s3_div_out_2_port, o(1) => s3_div_out_1_port
                           , o(0) => s3_div_out_0_port);
   MUXEXE : Mux4_DATA_SIZE32 port map( sel(1) => s3_exe_sel_1_port, sel(0) => 
                           sig_mul_port, din0(31) => s3_alu_out_31_port, 
                           din0(30) => s3_alu_out_30_port, din0(29) => 
                           s3_alu_out_29_port, din0(28) => s3_alu_out_28_port, 
                           din0(27) => s3_alu_out_27_port, din0(26) => 
                           s3_alu_out_26_port, din0(25) => s3_alu_out_25_port, 
                           din0(24) => s3_alu_out_24_port, din0(23) => 
                           s3_alu_out_23_port, din0(22) => s3_alu_out_22_port, 
                           din0(21) => s3_alu_out_21_port, din0(20) => 
                           s3_alu_out_20_port, din0(19) => s3_alu_out_19_port, 
                           din0(18) => s3_alu_out_18_port, din0(17) => 
                           s3_alu_out_17_port, din0(16) => s3_alu_out_16_port, 
                           din0(15) => s3_alu_out_15_port, din0(14) => 
                           s3_alu_out_14_port, din0(13) => s3_alu_out_13_port, 
                           din0(12) => s3_alu_out_12_port, din0(11) => 
                           s3_alu_out_11_port, din0(10) => s3_alu_out_10_port, 
                           din0(9) => s3_alu_out_9_port, din0(8) => 
                           s3_alu_out_8_port, din0(7) => s3_alu_out_7_port, 
                           din0(6) => s3_alu_out_6_port, din0(5) => 
                           s3_alu_out_5_port, din0(4) => s3_alu_out_4_port, 
                           din0(3) => s3_alu_out_3_port, din0(2) => 
                           s3_alu_out_2_port, din0(1) => s3_alu_out_1_port, 
                           din0(0) => s3_alu_out_0_port, din1(31) => 
                           s3_mul_out_31_port, din1(30) => s3_mul_out_30_port, 
                           din1(29) => s3_mul_out_29_port, din1(28) => 
                           s3_mul_out_28_port, din1(27) => s3_mul_out_27_port, 
                           din1(26) => s3_mul_out_26_port, din1(25) => 
                           s3_mul_out_25_port, din1(24) => s3_mul_out_24_port, 
                           din1(23) => s3_mul_out_23_port, din1(22) => 
                           s3_mul_out_22_port, din1(21) => s3_mul_out_21_port, 
                           din1(20) => s3_mul_out_20_port, din1(19) => 
                           s3_mul_out_19_port, din1(18) => s3_mul_out_18_port, 
                           din1(17) => s3_mul_out_17_port, din1(16) => 
                           s3_mul_out_16_port, din1(15) => s3_mul_out_15_port, 
                           din1(14) => s3_mul_out_14_port, din1(13) => 
                           s3_mul_out_13_port, din1(12) => s3_mul_out_12_port, 
                           din1(11) => s3_mul_out_11_port, din1(10) => 
                           s3_mul_out_10_port, din1(9) => s3_mul_out_9_port, 
                           din1(8) => s3_mul_out_8_port, din1(7) => 
                           s3_mul_out_7_port, din1(6) => s3_mul_out_6_port, 
                           din1(5) => s3_mul_out_5_port, din1(4) => 
                           s3_mul_out_4_port, din1(3) => s3_mul_out_3_port, 
                           din1(2) => s3_mul_out_2_port, din1(1) => 
                           s3_mul_out_1_port, din1(0) => s3_mul_out_0_port, 
                           din2(31) => s3_div_out_31_port, din2(30) => 
                           s3_div_out_30_port, din2(29) => s3_div_out_29_port, 
                           din2(28) => s3_div_out_28_port, din2(27) => 
                           s3_div_out_27_port, din2(26) => s3_div_out_26_port, 
                           din2(25) => s3_div_out_25_port, din2(24) => 
                           s3_div_out_24_port, din2(23) => s3_div_out_23_port, 
                           din2(22) => s3_div_out_22_port, din2(21) => 
                           s3_div_out_21_port, din2(20) => s3_div_out_20_port, 
                           din2(19) => s3_div_out_19_port, din2(18) => 
                           s3_div_out_18_port, din2(17) => s3_div_out_17_port, 
                           din2(16) => s3_div_out_16_port, din2(15) => 
                           s3_div_out_15_port, din2(14) => s3_div_out_14_port, 
                           din2(13) => s3_div_out_13_port, din2(12) => 
                           s3_div_out_12_port, din2(11) => s3_div_out_11_port, 
                           din2(10) => s3_div_out_10_port, din2(9) => 
                           s3_div_out_9_port, din2(8) => s3_div_out_8_port, 
                           din2(7) => s3_div_out_7_port, din2(6) => 
                           s3_div_out_6_port, din2(5) => s3_div_out_5_port, 
                           din2(4) => s3_div_out_4_port, din2(3) => 
                           s3_div_out_3_port, din2(2) => s3_div_out_2_port, 
                           din2(1) => s3_div_out_1_port, din2(0) => 
                           s3_div_out_0_port, din3(31) => X_Logic0_port, 
                           din3(30) => X_Logic0_port, din3(29) => X_Logic0_port
                           , din3(28) => X_Logic0_port, din3(27) => 
                           X_Logic0_port, din3(26) => X_Logic0_port, din3(25) 
                           => X_Logic0_port, din3(24) => X_Logic0_port, 
                           din3(23) => X_Logic0_port, din3(22) => X_Logic0_port
                           , din3(21) => X_Logic0_port, din3(20) => 
                           X_Logic0_port, din3(19) => X_Logic0_port, din3(18) 
                           => X_Logic0_port, din3(17) => X_Logic0_port, 
                           din3(16) => X_Logic0_port, din3(15) => X_Logic0_port
                           , din3(14) => X_Logic0_port, din3(13) => 
                           X_Logic0_port, din3(12) => X_Logic0_port, din3(11) 
                           => X_Logic0_port, din3(10) => X_Logic0_port, din3(9)
                           => X_Logic0_port, din3(8) => X_Logic0_port, din3(7) 
                           => X_Logic0_port, din3(6) => X_Logic0_port, din3(5) 
                           => X_Logic0_port, din3(4) => X_Logic0_port, din3(3) 
                           => X_Logic0_port, din3(2) => X_Logic0_port, din3(1) 
                           => X_Logic0_port, din3(0) => X_Logic0_port, dout(31)
                           => s3_exe_out_31_port, dout(30) => 
                           s3_exe_out_30_port, dout(29) => s3_exe_out_29_port, 
                           dout(28) => s3_exe_out_28_port, dout(27) => 
                           s3_exe_out_27_port, dout(26) => s3_exe_out_26_port, 
                           dout(25) => s3_exe_out_25_port, dout(24) => 
                           s3_exe_out_24_port, dout(23) => s3_exe_out_23_port, 
                           dout(22) => s3_exe_out_22_port, dout(21) => 
                           s3_exe_out_21_port, dout(20) => s3_exe_out_20_port, 
                           dout(19) => s3_exe_out_19_port, dout(18) => 
                           s3_exe_out_18_port, dout(17) => s3_exe_out_17_port, 
                           dout(16) => s3_exe_out_16_port, dout(15) => 
                           s3_exe_out_15_port, dout(14) => s3_exe_out_14_port, 
                           dout(13) => s3_exe_out_13_port, dout(12) => 
                           s3_exe_out_12_port, dout(11) => s3_exe_out_11_port, 
                           dout(10) => s3_exe_out_10_port, dout(9) => 
                           s3_exe_out_9_port, dout(8) => s3_exe_out_8_port, 
                           dout(7) => s3_exe_out_7_port, dout(6) => 
                           s3_exe_out_6_port, dout(5) => s3_exe_out_5_port, 
                           dout(4) => s3_exe_out_4_port, dout(3) => 
                           s3_exe_out_3_port, dout(2) => s3_exe_out_2_port, 
                           dout(1) => s3_exe_out_1_port, dout(0) => 
                           s3_exe_out_0_port);
   REG_ALU : Reg_DATA_SIZE32_7 port map( rst => rst, en => cw(10), clk => clk, 
                           din(31) => s3_exe_out_31_port, din(30) => 
                           s3_exe_out_30_port, din(29) => s3_exe_out_29_port, 
                           din(28) => s3_exe_out_28_port, din(27) => 
                           s3_exe_out_27_port, din(26) => s3_exe_out_26_port, 
                           din(25) => s3_exe_out_25_port, din(24) => 
                           s3_exe_out_24_port, din(23) => s3_exe_out_23_port, 
                           din(22) => s3_exe_out_22_port, din(21) => 
                           s3_exe_out_21_port, din(20) => s3_exe_out_20_port, 
                           din(19) => s3_exe_out_19_port, din(18) => 
                           s3_exe_out_18_port, din(17) => s3_exe_out_17_port, 
                           din(16) => s3_exe_out_16_port, din(15) => 
                           s3_exe_out_15_port, din(14) => s3_exe_out_14_port, 
                           din(13) => s3_exe_out_13_port, din(12) => 
                           s3_exe_out_12_port, din(11) => s3_exe_out_11_port, 
                           din(10) => s3_exe_out_10_port, din(9) => 
                           s3_exe_out_9_port, din(8) => s3_exe_out_8_port, 
                           din(7) => s3_exe_out_7_port, din(6) => 
                           s3_exe_out_6_port, din(5) => s3_exe_out_5_port, 
                           din(4) => s3_exe_out_4_port, din(3) => 
                           s3_exe_out_3_port, din(2) => s3_exe_out_2_port, 
                           din(1) => s3_exe_out_1_port, din(0) => 
                           s3_exe_out_0_port, dout(31) => data_addr_31_port, 
                           dout(30) => data_addr_30_port, dout(29) => 
                           data_addr_29_port, dout(28) => data_addr_28_port, 
                           dout(27) => data_addr_27_port, dout(26) => 
                           data_addr_26_port, dout(25) => data_addr_25_port, 
                           dout(24) => data_addr_24_port, dout(23) => 
                           data_addr_23_port, dout(22) => data_addr_22_port, 
                           dout(21) => data_addr_21_port, dout(20) => 
                           data_addr_20_port, dout(19) => data_addr_19_port, 
                           dout(18) => data_addr_18_port, dout(17) => 
                           data_addr_17_port, dout(16) => data_addr_16_port, 
                           dout(15) => data_addr_15_port, dout(14) => 
                           data_addr_14_port, dout(13) => data_addr_13_port, 
                           dout(12) => data_addr_12_port, dout(11) => 
                           data_addr_11_port, dout(10) => data_addr_10_port, 
                           dout(9) => data_addr_9_port, dout(8) => 
                           data_addr_8_port, dout(7) => data_addr_7_port, 
                           dout(6) => data_addr_6_port, dout(5) => 
                           data_addr_5_port, dout(4) => data_addr_4_port, 
                           dout(3) => data_addr_3_port, dout(2) => 
                           data_addr_2_port, dout(1) => data_addr_1_port, 
                           dout(0) => data_addr_0_port);
   REG_BB : Reg_DATA_SIZE32_6 port map( rst => rst, en => cw(10), clk => clk, 
                           din(31) => s3_b_fwd_31_port, din(30) => 
                           s3_b_fwd_30_port, din(29) => s3_b_fwd_29_port, 
                           din(28) => s3_b_fwd_28_port, din(27) => 
                           s3_b_fwd_27_port, din(26) => s3_b_fwd_26_port, 
                           din(25) => s3_b_fwd_25_port, din(24) => 
                           s3_b_fwd_24_port, din(23) => s3_b_fwd_23_port, 
                           din(22) => s3_b_fwd_22_port, din(21) => 
                           s3_b_fwd_21_port, din(20) => s3_b_fwd_20_port, 
                           din(19) => s3_b_fwd_19_port, din(18) => 
                           s3_b_fwd_18_port, din(17) => s3_b_fwd_17_port, 
                           din(16) => s3_b_fwd_16_port, din(15) => 
                           s3_b_fwd_15_port, din(14) => s3_b_fwd_14_port, 
                           din(13) => s3_b_fwd_13_port, din(12) => 
                           s3_b_fwd_12_port, din(11) => s3_b_fwd_11_port, 
                           din(10) => s3_b_fwd_10_port, din(9) => 
                           s3_b_fwd_9_port, din(8) => s3_b_fwd_8_port, din(7) 
                           => s3_b_fwd_7_port, din(6) => s3_b_fwd_6_port, 
                           din(5) => s3_b_fwd_5_port, din(4) => s3_b_fwd_4_port
                           , din(3) => s3_b_fwd_3_port, din(2) => 
                           s3_b_fwd_2_port, din(1) => s3_b_fwd_1_port, din(0) 
                           => s3_b_fwd_0_port, dout(31) => s4_b_fwd_31_port, 
                           dout(30) => s4_b_fwd_30_port, dout(29) => 
                           s4_b_fwd_29_port, dout(28) => s4_b_fwd_28_port, 
                           dout(27) => s4_b_fwd_27_port, dout(26) => 
                           s4_b_fwd_26_port, dout(25) => s4_b_fwd_25_port, 
                           dout(24) => s4_b_fwd_24_port, dout(23) => 
                           s4_b_fwd_23_port, dout(22) => s4_b_fwd_22_port, 
                           dout(21) => s4_b_fwd_21_port, dout(20) => 
                           s4_b_fwd_20_port, dout(19) => s4_b_fwd_19_port, 
                           dout(18) => s4_b_fwd_18_port, dout(17) => 
                           s4_b_fwd_17_port, dout(16) => s4_b_fwd_16_port, 
                           dout(15) => s4_b_fwd_15_port, dout(14) => 
                           s4_b_fwd_14_port, dout(13) => s4_b_fwd_13_port, 
                           dout(12) => s4_b_fwd_12_port, dout(11) => 
                           s4_b_fwd_11_port, dout(10) => s4_b_fwd_10_port, 
                           dout(9) => s4_b_fwd_9_port, dout(8) => 
                           s4_b_fwd_8_port, dout(7) => s4_b_fwd_7_port, dout(6)
                           => s4_b_fwd_6_port, dout(5) => s4_b_fwd_5_port, 
                           dout(4) => s4_b_fwd_4_port, dout(3) => 
                           s4_b_fwd_3_port, dout(2) => s4_b_fwd_2_port, dout(1)
                           => s4_b_fwd_1_port, dout(0) => s4_b_fwd_0_port);
   REG_B_ADDR_3 : Reg_DATA_SIZE5_4 port map( rst => rst, en => cw(10), clk => 
                           clk, din(4) => s3_rd2_addr_4_port, din(3) => 
                           s3_rd2_addr_3_port, din(2) => s3_rd2_addr_2_port, 
                           din(1) => s3_rd2_addr_1_port, din(0) => 
                           s3_rd2_addr_0_port, dout(4) => s4_rd2_addr_4_port, 
                           dout(3) => s4_rd2_addr_3_port, dout(2) => 
                           s4_rd2_addr_2_port, dout(1) => s4_rd2_addr_1_port, 
                           dout(0) => s4_rd2_addr_0_port);
   REG_WR3 : Reg_DATA_SIZE5_3 port map( rst => rst, en => cw(10), clk => clk, 
                           din(4) => s3_wr_addr_4_port, din(3) => 
                           s3_wr_addr_3_port, din(2) => s3_wr_addr_2_port, 
                           din(1) => s3_wr_addr_1_port, din(0) => 
                           s3_wr_addr_0_port, dout(4) => s4_wr_addr_4_port, 
                           dout(3) => s4_wr_addr_3_port, dout(2) => 
                           s4_wr_addr_2_port, dout(1) => s4_wr_addr_1_port, 
                           dout(0) => s4_wr_addr_0_port);
   REG_OPRD_A_WAIT : Reg_DATA_SIZE32_5 port map( rst => rst, en => 
                           X_Logic1_port, clk => clk, din(31) => 
                           s3_a_sel_31_port, din(30) => s3_a_sel_30_port, 
                           din(29) => s3_a_sel_29_port, din(28) => 
                           s3_a_sel_28_port, din(27) => s3_a_sel_27_port, 
                           din(26) => s3_a_sel_26_port, din(25) => 
                           s3_a_sel_25_port, din(24) => s3_a_sel_24_port, 
                           din(23) => s3_a_sel_23_port, din(22) => 
                           s3_a_sel_22_port, din(21) => s3_a_sel_21_port, 
                           din(20) => s3_a_sel_20_port, din(19) => 
                           s3_a_sel_19_port, din(18) => s3_a_sel_18_port, 
                           din(17) => s3_a_sel_17_port, din(16) => 
                           s3_a_sel_16_port, din(15) => s3_a_sel_15_port, 
                           din(14) => s3_a_sel_14_port, din(13) => 
                           s3_a_sel_13_port, din(12) => s3_a_sel_12_port, 
                           din(11) => s3_a_sel_11_port, din(10) => 
                           s3_a_sel_10_port, din(9) => s3_a_sel_9_port, din(8) 
                           => s3_a_sel_8_port, din(7) => s3_a_sel_7_port, 
                           din(6) => s3_a_sel_6_port, din(5) => s3_a_sel_5_port
                           , din(4) => s3_a_sel_4_port, din(3) => 
                           s3_a_sel_3_port, din(2) => s3_a_sel_2_port, din(1) 
                           => s3_a_sel_1_port, din(0) => s3_a_sel_0_port, 
                           dout(31) => s4_a_31_port, dout(30) => s4_a_30_port, 
                           dout(29) => s4_a_29_port, dout(28) => s4_a_28_port, 
                           dout(27) => s4_a_27_port, dout(26) => s4_a_26_port, 
                           dout(25) => s4_a_25_port, dout(24) => s4_a_24_port, 
                           dout(23) => s4_a_23_port, dout(22) => s4_a_22_port, 
                           dout(21) => s4_a_21_port, dout(20) => s4_a_20_port, 
                           dout(19) => s4_a_19_port, dout(18) => s4_a_18_port, 
                           dout(17) => s4_a_17_port, dout(16) => s4_a_16_port, 
                           dout(15) => s4_a_15_port, dout(14) => s4_a_14_port, 
                           dout(13) => s4_a_13_port, dout(12) => s4_a_12_port, 
                           dout(11) => s4_a_11_port, dout(10) => s4_a_10_port, 
                           dout(9) => s4_a_9_port, dout(8) => s4_a_8_port, 
                           dout(7) => s4_a_7_port, dout(6) => s4_a_6_port, 
                           dout(5) => s4_a_5_port, dout(4) => s4_a_4_port, 
                           dout(3) => s4_a_3_port, dout(2) => s4_a_2_port, 
                           dout(1) => s4_a_1_port, dout(0) => s4_a_0_port);
   REG_OPRD_B_WAIT : Reg_DATA_SIZE32_4 port map( rst => rst, en => 
                           X_Logic1_port, clk => clk, din(31) => 
                           s3_b_sel_31_port, din(30) => s3_b_sel_30_port, 
                           din(29) => s3_b_sel_29_port, din(28) => 
                           s3_b_sel_28_port, din(27) => s3_b_sel_27_port, 
                           din(26) => s3_b_sel_26_port, din(25) => 
                           s3_b_sel_25_port, din(24) => s3_b_sel_24_port, 
                           din(23) => s3_b_sel_23_port, din(22) => 
                           s3_b_sel_22_port, din(21) => s3_b_sel_21_port, 
                           din(20) => s3_b_sel_20_port, din(19) => 
                           s3_b_sel_19_port, din(18) => s3_b_sel_18_port, 
                           din(17) => s3_b_sel_17_port, din(16) => 
                           s3_b_sel_16_port, din(15) => s3_b_sel_15_port, 
                           din(14) => s3_b_sel_14_port, din(13) => 
                           s3_b_sel_13_port, din(12) => s3_b_sel_12_port, 
                           din(11) => s3_b_sel_11_port, din(10) => 
                           s3_b_sel_10_port, din(9) => s3_b_sel_9_port, din(8) 
                           => s3_b_sel_8_port, din(7) => s3_b_sel_7_port, 
                           din(6) => s3_b_sel_6_port, din(5) => s3_b_sel_5_port
                           , din(4) => s3_b_sel_4_port, din(3) => 
                           s3_b_sel_3_port, din(2) => s3_b_sel_2_port, din(1) 
                           => s3_b_sel_1_port, din(0) => s3_b_sel_0_port, 
                           dout(31) => s4_b_31_port, dout(30) => s4_b_30_port, 
                           dout(29) => s4_b_29_port, dout(28) => s4_b_28_port, 
                           dout(27) => s4_b_27_port, dout(26) => s4_b_26_port, 
                           dout(25) => s4_b_25_port, dout(24) => s4_b_24_port, 
                           dout(23) => s4_b_23_port, dout(22) => s4_b_22_port, 
                           dout(21) => s4_b_21_port, dout(20) => s4_b_20_port, 
                           dout(19) => s4_b_19_port, dout(18) => s4_b_18_port, 
                           dout(17) => s4_b_17_port, dout(16) => s4_b_16_port, 
                           dout(15) => s4_b_15_port, dout(14) => s4_b_14_port, 
                           dout(13) => s4_b_13_port, dout(12) => s4_b_12_port, 
                           dout(11) => s4_b_11_port, dout(10) => s4_b_10_port, 
                           dout(9) => s4_b_9_port, dout(8) => s4_b_8_port, 
                           dout(7) => s4_b_7_port, dout(6) => s4_b_6_port, 
                           dout(5) => s4_b_5_port, dout(4) => s4_b_4_port, 
                           dout(3) => s4_b_3_port, dout(2) => s4_b_2_port, 
                           dout(1) => s4_b_1_port, dout(0) => s4_b_0_port);
   FWDMUX_BB : FwdMux2_DATA_SIZE32_REG_ADDR_SIZE5_1 port map( reg_c(31) => 
                           s4_b_fwd_31_port, reg_c(30) => s4_b_fwd_30_port, 
                           reg_c(29) => s4_b_fwd_29_port, reg_c(28) => 
                           s4_b_fwd_28_port, reg_c(27) => s4_b_fwd_27_port, 
                           reg_c(26) => s4_b_fwd_26_port, reg_c(25) => 
                           s4_b_fwd_25_port, reg_c(24) => s4_b_fwd_24_port, 
                           reg_c(23) => s4_b_fwd_23_port, reg_c(22) => 
                           s4_b_fwd_22_port, reg_c(21) => s4_b_fwd_21_port, 
                           reg_c(20) => s4_b_fwd_20_port, reg_c(19) => 
                           s4_b_fwd_19_port, reg_c(18) => s4_b_fwd_18_port, 
                           reg_c(17) => s4_b_fwd_17_port, reg_c(16) => 
                           s4_b_fwd_16_port, reg_c(15) => s4_b_fwd_15_port, 
                           reg_c(14) => s4_b_fwd_14_port, reg_c(13) => 
                           s4_b_fwd_13_port, reg_c(12) => s4_b_fwd_12_port, 
                           reg_c(11) => s4_b_fwd_11_port, reg_c(10) => 
                           s4_b_fwd_10_port, reg_c(9) => s4_b_fwd_9_port, 
                           reg_c(8) => s4_b_fwd_8_port, reg_c(7) => 
                           s4_b_fwd_7_port, reg_c(6) => s4_b_fwd_6_port, 
                           reg_c(5) => s4_b_fwd_5_port, reg_c(4) => 
                           s4_b_fwd_4_port, reg_c(3) => s4_b_fwd_3_port, 
                           reg_c(2) => s4_b_fwd_2_port, reg_c(1) => 
                           s4_b_fwd_1_port, reg_c(0) => s4_b_fwd_0_port, 
                           reg_f(31) => s5_result_31_port, reg_f(30) => 
                           s5_result_30_port, reg_f(29) => s5_result_29_port, 
                           reg_f(28) => s5_result_28_port, reg_f(27) => 
                           s5_result_27_port, reg_f(26) => s5_result_26_port, 
                           reg_f(25) => s5_result_25_port, reg_f(24) => 
                           s5_result_24_port, reg_f(23) => s5_result_23_port, 
                           reg_f(22) => s5_result_22_port, reg_f(21) => 
                           s5_result_21_port, reg_f(20) => s5_result_20_port, 
                           reg_f(19) => s5_result_19_port, reg_f(18) => 
                           s5_result_18_port, reg_f(17) => s5_result_17_port, 
                           reg_f(16) => s5_result_16_port, reg_f(15) => 
                           s5_result_15_port, reg_f(14) => s5_result_14_port, 
                           reg_f(13) => s5_result_13_port, reg_f(12) => 
                           s5_result_12_port, reg_f(11) => s5_result_11_port, 
                           reg_f(10) => s5_result_10_port, reg_f(9) => 
                           s5_result_9_port, reg_f(8) => s5_result_8_port, 
                           reg_f(7) => s5_result_7_port, reg_f(6) => 
                           s5_result_6_port, reg_f(5) => s5_result_5_port, 
                           reg_f(4) => s5_result_4_port, reg_f(3) => 
                           s5_result_3_port, reg_f(2) => s5_result_2_port, 
                           reg_f(1) => s5_result_1_port, reg_f(0) => 
                           s5_result_0_port, reg_ff(31) => s6_result_31_port, 
                           reg_ff(30) => s6_result_30_port, reg_ff(29) => 
                           s6_result_29_port, reg_ff(28) => s6_result_28_port, 
                           reg_ff(27) => s6_result_27_port, reg_ff(26) => 
                           s6_result_26_port, reg_ff(25) => s6_result_25_port, 
                           reg_ff(24) => s6_result_24_port, reg_ff(23) => 
                           s6_result_23_port, reg_ff(22) => s6_result_22_port, 
                           reg_ff(21) => s6_result_21_port, reg_ff(20) => 
                           s6_result_20_port, reg_ff(19) => s6_result_19_port, 
                           reg_ff(18) => s6_result_18_port, reg_ff(17) => 
                           s6_result_17_port, reg_ff(16) => s6_result_16_port, 
                           reg_ff(15) => s6_result_15_port, reg_ff(14) => 
                           s6_result_14_port, reg_ff(13) => s6_result_13_port, 
                           reg_ff(12) => s6_result_12_port, reg_ff(11) => 
                           s6_result_11_port, reg_ff(10) => s6_result_10_port, 
                           reg_ff(9) => s6_result_9_port, reg_ff(8) => 
                           s6_result_8_port, reg_ff(7) => s6_result_7_port, 
                           reg_ff(6) => s6_result_6_port, reg_ff(5) => 
                           s6_result_5_port, reg_ff(4) => s6_result_4_port, 
                           reg_ff(3) => s6_result_3_port, reg_ff(2) => 
                           s6_result_2_port, reg_ff(1) => s6_result_1_port, 
                           reg_ff(0) => s6_result_0_port, addr_c(4) => 
                           s4_rd2_addr_4_port, addr_c(3) => s4_rd2_addr_3_port,
                           addr_c(2) => s4_rd2_addr_2_port, addr_c(1) => 
                           s4_rd2_addr_1_port, addr_c(0) => s4_rd2_addr_0_port,
                           addr_f(4) => s5_wr_addr_4_port, addr_f(3) => 
                           s5_wr_addr_3_port, addr_f(2) => s5_wr_addr_2_port, 
                           addr_f(1) => s5_wr_addr_1_port, addr_f(0) => 
                           s5_wr_addr_0_port, addr_ff(4) => s6_wr_addr_4_port, 
                           addr_ff(3) => s6_wr_addr_3_port, addr_ff(2) => 
                           s6_wr_addr_2_port, addr_ff(1) => s6_wr_addr_1_port, 
                           addr_ff(0) => s6_wr_addr_0_port, valid_f => cw(19), 
                           valid_ff => s6_en_wb, dirty_f => X_Logic0_port, 
                           dirty_ff => X_Logic0_port, en => cw(14), output(31) 
                           => data_o_val(31), output(30) => data_o_val(30), 
                           output(29) => data_o_val(29), output(28) => 
                           data_o_val(28), output(27) => data_o_val(27), 
                           output(26) => data_o_val(26), output(25) => 
                           data_o_val(25), output(24) => data_o_val(24), 
                           output(23) => data_o_val(23), output(22) => 
                           data_o_val(22), output(21) => data_o_val(21), 
                           output(20) => data_o_val(20), output(19) => 
                           data_o_val(19), output(18) => data_o_val(18), 
                           output(17) => data_o_val(17), output(16) => 
                           data_o_val(16), output(15) => data_o_val(15), 
                           output(14) => data_o_val(14), output(13) => 
                           data_o_val(13), output(12) => data_o_val(12), 
                           output(11) => data_o_val(11), output(10) => 
                           data_o_val(10), output(9) => data_o_val(9), 
                           output(8) => data_o_val(8), output(7) => 
                           data_o_val(7), output(6) => data_o_val(6), output(5)
                           => data_o_val(5), output(4) => data_o_val(4), 
                           output(3) => data_o_val(3), output(2) => 
                           data_o_val(2), output(1) => data_o_val(1), output(0)
                           => data_o_val(0), match_dirty_f => net1283, 
                           match_dirty_ff => net1284);
   MUX_RESULT : Mux_DATA_SIZE32_2 port map( sel => cw(15), din0(31) => 
                           data_addr_31_port, din0(30) => data_addr_30_port, 
                           din0(29) => data_addr_29_port, din0(28) => 
                           data_addr_28_port, din0(27) => data_addr_27_port, 
                           din0(26) => data_addr_26_port, din0(25) => 
                           data_addr_25_port, din0(24) => data_addr_24_port, 
                           din0(23) => data_addr_23_port, din0(22) => 
                           data_addr_22_port, din0(21) => data_addr_21_port, 
                           din0(20) => data_addr_20_port, din0(19) => 
                           data_addr_19_port, din0(18) => data_addr_18_port, 
                           din0(17) => data_addr_17_port, din0(16) => 
                           data_addr_16_port, din0(15) => data_addr_15_port, 
                           din0(14) => data_addr_14_port, din0(13) => 
                           data_addr_13_port, din0(12) => data_addr_12_port, 
                           din0(11) => data_addr_11_port, din0(10) => 
                           data_addr_10_port, din0(9) => data_addr_9_port, 
                           din0(8) => data_addr_8_port, din0(7) => 
                           data_addr_7_port, din0(6) => data_addr_6_port, 
                           din0(5) => data_addr_5_port, din0(4) => 
                           data_addr_4_port, din0(3) => data_addr_3_port, 
                           din0(2) => data_addr_2_port, din0(1) => 
                           data_addr_1_port, din0(0) => data_addr_0_port, 
                           din1(31) => data_i_val(31), din1(30) => 
                           data_i_val(30), din1(29) => data_i_val(29), din1(28)
                           => data_i_val(28), din1(27) => data_i_val(27), 
                           din1(26) => data_i_val(26), din1(25) => 
                           data_i_val(25), din1(24) => data_i_val(24), din1(23)
                           => data_i_val(23), din1(22) => data_i_val(22), 
                           din1(21) => data_i_val(21), din1(20) => 
                           data_i_val(20), din1(19) => data_i_val(19), din1(18)
                           => data_i_val(18), din1(17) => data_i_val(17), 
                           din1(16) => data_i_val(16), din1(15) => 
                           data_i_val(15), din1(14) => data_i_val(14), din1(13)
                           => data_i_val(13), din1(12) => data_i_val(12), 
                           din1(11) => data_i_val(11), din1(10) => 
                           data_i_val(10), din1(9) => data_i_val(9), din1(8) =>
                           data_i_val(8), din1(7) => data_i_val(7), din1(6) => 
                           data_i_val(6), din1(5) => data_i_val(5), din1(4) => 
                           data_i_val(4), din1(3) => data_i_val(3), din1(2) => 
                           data_i_val(2), din1(1) => data_i_val(1), din1(0) => 
                           data_i_val(0), dout(31) => s4_result_31_port, 
                           dout(30) => s4_result_30_port, dout(29) => 
                           s4_result_29_port, dout(28) => s4_result_28_port, 
                           dout(27) => s4_result_27_port, dout(26) => 
                           s4_result_26_port, dout(25) => s4_result_25_port, 
                           dout(24) => s4_result_24_port, dout(23) => 
                           s4_result_23_port, dout(22) => s4_result_22_port, 
                           dout(21) => s4_result_21_port, dout(20) => 
                           s4_result_20_port, dout(19) => s4_result_19_port, 
                           dout(18) => s4_result_18_port, dout(17) => 
                           s4_result_17_port, dout(16) => s4_result_16_port, 
                           dout(15) => s4_result_15_port, dout(14) => 
                           s4_result_14_port, dout(13) => s4_result_13_port, 
                           dout(12) => s4_result_12_port, dout(11) => 
                           s4_result_11_port, dout(10) => s4_result_10_port, 
                           dout(9) => s4_result_9_port, dout(8) => 
                           s4_result_8_port, dout(7) => s4_result_7_port, 
                           dout(6) => s4_result_6_port, dout(5) => 
                           s4_result_5_port, dout(4) => s4_result_4_port, 
                           dout(3) => s4_result_3_port, dout(2) => 
                           s4_result_2_port, dout(1) => s4_result_1_port, 
                           dout(0) => s4_result_0_port);
   REG_RESULT : Reg_DATA_SIZE32_3 port map( rst => rst, en => cw(18), clk => 
                           clk, din(31) => s4_result_31_port, din(30) => 
                           s4_result_30_port, din(29) => s4_result_29_port, 
                           din(28) => s4_result_28_port, din(27) => 
                           s4_result_27_port, din(26) => s4_result_26_port, 
                           din(25) => s4_result_25_port, din(24) => 
                           s4_result_24_port, din(23) => s4_result_23_port, 
                           din(22) => s4_result_22_port, din(21) => 
                           s4_result_21_port, din(20) => s4_result_20_port, 
                           din(19) => s4_result_19_port, din(18) => 
                           s4_result_18_port, din(17) => s4_result_17_port, 
                           din(16) => s4_result_16_port, din(15) => 
                           s4_result_15_port, din(14) => s4_result_14_port, 
                           din(13) => s4_result_13_port, din(12) => 
                           s4_result_12_port, din(11) => s4_result_11_port, 
                           din(10) => s4_result_10_port, din(9) => 
                           s4_result_9_port, din(8) => s4_result_8_port, din(7)
                           => s4_result_7_port, din(6) => s4_result_6_port, 
                           din(5) => s4_result_5_port, din(4) => 
                           s4_result_4_port, din(3) => s4_result_3_port, din(2)
                           => s4_result_2_port, din(1) => s4_result_1_port, 
                           din(0) => s4_result_0_port, dout(31) => 
                           s5_result_31_port, dout(30) => s5_result_30_port, 
                           dout(29) => s5_result_29_port, dout(28) => 
                           s5_result_28_port, dout(27) => s5_result_27_port, 
                           dout(26) => s5_result_26_port, dout(25) => 
                           s5_result_25_port, dout(24) => s5_result_24_port, 
                           dout(23) => s5_result_23_port, dout(22) => 
                           s5_result_22_port, dout(21) => s5_result_21_port, 
                           dout(20) => s5_result_20_port, dout(19) => 
                           s5_result_19_port, dout(18) => s5_result_18_port, 
                           dout(17) => s5_result_17_port, dout(16) => 
                           s5_result_16_port, dout(15) => s5_result_15_port, 
                           dout(14) => s5_result_14_port, dout(13) => 
                           s5_result_13_port, dout(12) => s5_result_12_port, 
                           dout(11) => s5_result_11_port, dout(10) => 
                           s5_result_10_port, dout(9) => s5_result_9_port, 
                           dout(8) => s5_result_8_port, dout(7) => 
                           s5_result_7_port, dout(6) => s5_result_6_port, 
                           dout(5) => s5_result_5_port, dout(4) => 
                           s5_result_4_port, dout(3) => s5_result_3_port, 
                           dout(2) => s5_result_2_port, dout(1) => 
                           s5_result_1_port, dout(0) => s5_result_0_port);
   REG_WR4 : Reg_DATA_SIZE5_2 port map( rst => rst, en => cw(18), clk => clk, 
                           din(4) => s4_wr_addr_4_port, din(3) => 
                           s4_wr_addr_3_port, din(2) => s4_wr_addr_2_port, 
                           din(1) => s4_wr_addr_1_port, din(0) => 
                           s4_wr_addr_0_port, dout(4) => s5_wr_addr_4_port, 
                           dout(3) => s5_wr_addr_3_port, dout(2) => 
                           s5_wr_addr_2_port, dout(1) => s5_wr_addr_1_port, 
                           dout(0) => s5_wr_addr_0_port);
   REG_RESULT5 : Reg_DATA_SIZE32_2 port map( rst => rst, en => cw(19), clk => 
                           clk, din(31) => s5_result_31_port, din(30) => 
                           s5_result_30_port, din(29) => s5_result_29_port, 
                           din(28) => s5_result_28_port, din(27) => 
                           s5_result_27_port, din(26) => s5_result_26_port, 
                           din(25) => s5_result_25_port, din(24) => 
                           s5_result_24_port, din(23) => s5_result_23_port, 
                           din(22) => s5_result_22_port, din(21) => 
                           s5_result_21_port, din(20) => s5_result_20_port, 
                           din(19) => s5_result_19_port, din(18) => 
                           s5_result_18_port, din(17) => s5_result_17_port, 
                           din(16) => s5_result_16_port, din(15) => 
                           s5_result_15_port, din(14) => s5_result_14_port, 
                           din(13) => s5_result_13_port, din(12) => 
                           s5_result_12_port, din(11) => s5_result_11_port, 
                           din(10) => s5_result_10_port, din(9) => 
                           s5_result_9_port, din(8) => s5_result_8_port, din(7)
                           => s5_result_7_port, din(6) => s5_result_6_port, 
                           din(5) => s5_result_5_port, din(4) => 
                           s5_result_4_port, din(3) => s5_result_3_port, din(2)
                           => s5_result_2_port, din(1) => s5_result_1_port, 
                           din(0) => s5_result_0_port, dout(31) => 
                           s6_result_31_port, dout(30) => s6_result_30_port, 
                           dout(29) => s6_result_29_port, dout(28) => 
                           s6_result_28_port, dout(27) => s6_result_27_port, 
                           dout(26) => s6_result_26_port, dout(25) => 
                           s6_result_25_port, dout(24) => s6_result_24_port, 
                           dout(23) => s6_result_23_port, dout(22) => 
                           s6_result_22_port, dout(21) => s6_result_21_port, 
                           dout(20) => s6_result_20_port, dout(19) => 
                           s6_result_19_port, dout(18) => s6_result_18_port, 
                           dout(17) => s6_result_17_port, dout(16) => 
                           s6_result_16_port, dout(15) => s6_result_15_port, 
                           dout(14) => s6_result_14_port, dout(13) => 
                           s6_result_13_port, dout(12) => s6_result_12_port, 
                           dout(11) => s6_result_11_port, dout(10) => 
                           s6_result_10_port, dout(9) => s6_result_9_port, 
                           dout(8) => s6_result_8_port, dout(7) => 
                           s6_result_7_port, dout(6) => s6_result_6_port, 
                           dout(5) => s6_result_5_port, dout(4) => 
                           s6_result_4_port, dout(3) => s6_result_3_port, 
                           dout(2) => s6_result_2_port, dout(1) => 
                           s6_result_1_port, dout(0) => s6_result_0_port);
   REG_WR5 : Reg_DATA_SIZE5_1 port map( rst => rst, en => cw(19), clk => clk, 
                           din(4) => s5_wr_addr_4_port, din(3) => 
                           s5_wr_addr_3_port, din(2) => s5_wr_addr_2_port, 
                           din(1) => s5_wr_addr_1_port, din(0) => 
                           s5_wr_addr_0_port, dout(4) => s6_wr_addr_4_port, 
                           dout(3) => s6_wr_addr_3_port, dout(2) => 
                           s6_wr_addr_2_port, dout(1) => s6_wr_addr_1_port, 
                           dout(0) => s6_wr_addr_0_port);
   s4_reg_a_wait_reg : DFF_X2 port map( D => s3_reg_a_wait, CK => clk, Q => 
                           s4_reg_a_wait, QN => n2);
   s4_reg_b_wait_reg : DFF_X2 port map( D => s3_reg_b_wait, CK => clk, Q => 
                           s4_reg_b_wait, QN => n1);
   U3 : NAND4_X2 port map( A1 => n18, A2 => n37, A3 => istr_val(26), A4 => n38,
                           ZN => n19);
   U4 : INV_X1 port map( A => n3, ZN => sig_sqrt_port);
   U5 : OR2_X1 port map( A1 => s3_reg_a_wait, A2 => s3_reg_b_wait, ZN => 
                           sig_ral_port);
   U6 : INV_X1 port map( A => n4, ZN => sig_mul_port);
   U7 : INV_X1 port map( A => n5, ZN => sig_div);
   U8 : NOR2_X1 port map( A1 => n4, A2 => n6, ZN => s3_mul_sign);
   U9 : NAND3_X1 port map( A1 => n7, A2 => n8, A3 => n9, ZN => n4);
   U10 : NAND2_X1 port map( A1 => n3, A2 => n5, ZN => s3_exe_sel_1_port);
   U11 : NAND4_X1 port map( A1 => calu(2), A2 => n9, A3 => n6, A4 => n7, ZN => 
                           n3);
   U12 : INV_X1 port map( A => calu(1), ZN => n7);
   U13 : NOR2_X1 port map( A1 => n6, A2 => n5, ZN => s3_div_sign);
   U14 : NAND3_X1 port map( A1 => n9, A2 => n8, A3 => calu(1), ZN => n5);
   U15 : INV_X1 port map( A => calu(2), ZN => n8);
   U16 : NOR2_X1 port map( A1 => n10, A2 => calu(4), ZN => n9);
   U17 : INV_X1 port map( A => calu(3), ZN => n10);
   U18 : INV_X1 port map( A => calu(0), ZN => n6);
   U19 : NOR2_X1 port map( A1 => cw(7), A2 => n11, ZN => s3_b_sel_ff_en);
   U20 : INV_X1 port map( A => s3_a_sel_ff_en, ZN => n11);
   U21 : NOR2_X1 port map( A1 => cw(7), A2 => n12, ZN => s3_b_sel_f_en);
   U22 : INV_X1 port map( A => s3_a_sel_f_en, ZN => n12);
   U23 : NOR2_X1 port map( A1 => n13, A2 => s3_jump_flag, ZN => s3_a_sel_ff_en)
                           ;
   U24 : NOR2_X1 port map( A1 => n14, A2 => s3_jump_flag, ZN => s3_a_sel_f_en);
   U25 : NAND4_X1 port map( A1 => n15, A2 => n16, A3 => n17, A4 => n18, ZN => 
                           s2_wr_addr_sel);
   U26 : OR2_X1 port map( A1 => cw(19), A2 => cw(6), ZN => s2_rf_en);
   U27 : AND2_X1 port map( A1 => s2_imm_l_ext_9_port, A2 => n19, ZN => 
                           s2_imm_i_ext_9_port);
   U28 : AND2_X1 port map( A1 => s2_imm_l_ext_8_port, A2 => n19, ZN => 
                           s2_imm_i_ext_8_port);
   U29 : AND2_X1 port map( A1 => s2_imm_l_ext_7_port, A2 => n19, ZN => 
                           s2_imm_i_ext_7_port);
   U30 : AND2_X1 port map( A1 => s2_imm_l_ext_6_port, A2 => n19, ZN => 
                           s2_imm_i_ext_6_port);
   U31 : AND2_X1 port map( A1 => s2_imm_l_ext_5_port, A2 => n19, ZN => 
                           s2_imm_i_ext_5_port);
   U32 : AND2_X1 port map( A1 => s2_imm_l_ext_4_port, A2 => n19, ZN => 
                           s2_imm_i_ext_4_port);
   U33 : AND2_X1 port map( A1 => s2_imm_l_ext_3_port, A2 => n19, ZN => 
                           s2_imm_i_ext_3_port);
   U34 : OAI21_X1 port map( B1 => n19, B2 => n20, A => n21, ZN => 
                           s2_imm_i_ext_31_port);
   U35 : INV_X1 port map( A => istr_val(15), ZN => n20);
   U36 : OAI21_X1 port map( B1 => n19, B2 => n22, A => n21, ZN => 
                           s2_imm_i_ext_30_port);
   U37 : INV_X1 port map( A => istr_val(14), ZN => n22);
   U38 : AND2_X1 port map( A1 => s2_imm_l_ext_2_port, A2 => n19, ZN => 
                           s2_imm_i_ext_2_port);
   U39 : OAI21_X1 port map( B1 => n19, B2 => n23, A => n21, ZN => 
                           s2_imm_i_ext_29_port);
   U40 : INV_X1 port map( A => istr_val(13), ZN => n23);
   U41 : OAI21_X1 port map( B1 => n19, B2 => n24, A => n21, ZN => 
                           s2_imm_i_ext_28_port);
   U42 : INV_X1 port map( A => istr_val(12), ZN => n24);
   U43 : OAI21_X1 port map( B1 => n19, B2 => n25, A => n21, ZN => 
                           s2_imm_i_ext_27_port);
   U44 : INV_X1 port map( A => istr_val(11), ZN => n25);
   U45 : OAI21_X1 port map( B1 => n19, B2 => n26, A => n21, ZN => 
                           s2_imm_i_ext_26_port);
   U46 : INV_X1 port map( A => istr_val(10), ZN => n26);
   U47 : OAI21_X1 port map( B1 => n19, B2 => n27, A => n21, ZN => 
                           s2_imm_i_ext_25_port);
   U48 : INV_X1 port map( A => istr_val(9), ZN => n27);
   U49 : OAI21_X1 port map( B1 => n19, B2 => n28, A => n21, ZN => 
                           s2_imm_i_ext_24_port);
   U50 : INV_X1 port map( A => istr_val(8), ZN => n28);
   U51 : OAI21_X1 port map( B1 => n19, B2 => n29, A => n21, ZN => 
                           s2_imm_i_ext_23_port);
   U52 : INV_X1 port map( A => istr_val(7), ZN => n29);
   U53 : OAI21_X1 port map( B1 => n19, B2 => n30, A => n21, ZN => 
                           s2_imm_i_ext_22_port);
   U54 : INV_X1 port map( A => istr_val(6), ZN => n30);
   U55 : OAI21_X1 port map( B1 => n19, B2 => n31, A => n21, ZN => 
                           s2_imm_i_ext_21_port);
   U56 : INV_X1 port map( A => istr_val(5), ZN => n31);
   U57 : OAI21_X1 port map( B1 => n19, B2 => n32, A => n21, ZN => 
                           s2_imm_i_ext_20_port);
   U58 : INV_X1 port map( A => istr_val(4), ZN => n32);
   U59 : AND2_X1 port map( A1 => s2_imm_l_ext_1_port, A2 => n19, ZN => 
                           s2_imm_i_ext_1_port);
   U60 : OAI21_X1 port map( B1 => n19, B2 => n33, A => n21, ZN => 
                           s2_imm_i_ext_19_port);
   U61 : INV_X1 port map( A => istr_val(3), ZN => n33);
   U62 : OAI21_X1 port map( B1 => n19, B2 => n34, A => n21, ZN => 
                           s2_imm_i_ext_18_port);
   U63 : INV_X1 port map( A => istr_val(2), ZN => n34);
   U64 : OAI21_X1 port map( B1 => n19, B2 => n35, A => n21, ZN => 
                           s2_imm_i_ext_17_port);
   U65 : INV_X1 port map( A => istr_val(1), ZN => n35);
   U66 : OAI21_X1 port map( B1 => n19, B2 => n36, A => n21, ZN => 
                           s2_imm_i_ext_16_port);
   U67 : NAND2_X1 port map( A1 => s2_imm_l_ext_31_port, A2 => n19, ZN => n21);
   U68 : INV_X1 port map( A => istr_val(0), ZN => n36);
   U69 : AND2_X1 port map( A1 => s2_imm_l_ext_15_port, A2 => n19, ZN => 
                           s2_imm_i_ext_15_port);
   U70 : AND2_X1 port map( A1 => s2_imm_l_ext_14_port, A2 => n19, ZN => 
                           s2_imm_i_ext_14_port);
   U71 : AND2_X1 port map( A1 => s2_imm_l_ext_13_port, A2 => n19, ZN => 
                           s2_imm_i_ext_13_port);
   U72 : AND2_X1 port map( A1 => s2_imm_l_ext_12_port, A2 => n19, ZN => 
                           s2_imm_i_ext_12_port);
   U73 : AND2_X1 port map( A1 => s2_imm_l_ext_11_port, A2 => n19, ZN => 
                           s2_imm_i_ext_11_port);
   U74 : AND2_X1 port map( A1 => s2_imm_l_ext_10_port, A2 => n19, ZN => 
                           s2_imm_i_ext_10_port);
   U75 : AND2_X1 port map( A1 => s2_imm_l_ext_0_port, A2 => n19, ZN => 
                           s2_imm_i_ext_0_port);
   U76 : AND3_X1 port map( A1 => istr_val(29), A2 => istr_val(27), A3 => 
                           istr_val(28), ZN => n38);
   U77 : INV_X1 port map( A => istr_val(31), ZN => n37);
   U78 : NOR2_X1 port map( A1 => n14, A2 => n39, ZN => s2_a_ff_j_en);
   U79 : NOR3_X1 port map( A1 => n40, A2 => n14, A3 => n41, ZN => s2_a_ff_b_en)
                           ;
   U80 : INV_X1 port map( A => cw(17), ZN => n14);
   U81 : NOR2_X1 port map( A1 => n39, A2 => n42, ZN => s2_a_f_j_en);
   U82 : NAND4_X1 port map( A1 => istr_val(30), A2 => istr_val(27), A3 => n15, 
                           A4 => n17, ZN => n39);
   U83 : NOR3_X1 port map( A1 => n42, A2 => n41, A3 => n40, ZN => s2_a_f_b_en);
   U84 : INV_X1 port map( A => cw(9), ZN => n42);
   U85 : MUX2_X1 port map( A => s3_jump_flag, B => n43, S => cw(6), Z => n48);
   U86 : AOI21_X1 port map( B1 => n40, B2 => n46, A => n41, ZN => n43);
   U87 : INV_X1 port map( A => n15, ZN => n41);
   U88 : NOR2_X1 port map( A1 => istr_val(29), A2 => istr_val(31), ZN => n15);
   U89 : NAND2_X1 port map( A1 => istr_val(27), A2 => n17, ZN => n46);
   U90 : INV_X1 port map( A => istr_val(28), ZN => n17);
   U91 : NAND3_X1 port map( A1 => n16, A2 => n18, A3 => istr_val(28), ZN => n40
                           );
   U92 : INV_X1 port map( A => istr_val(30), ZN => n18);
   U93 : INV_X1 port map( A => istr_val(27), ZN => n16);
   U94 : NAND2_X1 port map( A1 => n44, A2 => n13, ZN => n45);
   U95 : INV_X1 port map( A => cw(19), ZN => n13);

end SYN_data_path_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity 
   ControlUnit_ISTR_SIZE32_DATA_SIZE32_OPCD_SIZE6_FUNC_SIZE11_CWRD_SIZE20_CALU_SIZE5_ADDR_SIZE32 
   is

   port( clk, rst : in std_logic;  ir, pc, reg_a, ld_a : in std_logic_vector 
         (31 downto 0);  sig_bal : in std_logic;  sig_bpw : out std_logic;  
         sig_jral, sig_ral, sig_mul, sig_div, sig_sqrt : in std_logic;  cw : 
         out std_logic_vector (19 downto 0);  calu : out std_logic_vector (4 
         downto 0));

end 
   ControlUnit_ISTR_SIZE32_DATA_SIZE32_OPCD_SIZE6_FUNC_SIZE11_CWRD_SIZE20_CALU_SIZE5_ADDR_SIZE32;

architecture SYN_control_unit_arch of 
   ControlUnit_ISTR_SIZE32_DATA_SIZE32_OPCD_SIZE6_FUNC_SIZE11_CWRD_SIZE20_CALU_SIZE5_ADDR_SIZE32 
   is

   component Branch_DATA_SIZE32_OPCD_SIZE6_ADDR_SIZE32
      port( rst, clk : in std_logic;  reg_a, ld_a : in std_logic_vector (31 
            downto 0);  opcd : in std_logic_vector (5 downto 0);  addr : in 
            std_logic_vector (31 downto 0);  sig_bal : in std_logic;  sig_bpw, 
            sig_brt : out std_logic);
   end component;
   
   component StallGenerator_CWRD_SIZE20
      port( rst, clk, sig_ral, sig_bpw, sig_jral, sig_mul, sig_div, sig_sqrt : 
            in std_logic;  stall_flag : out std_logic_vector (4 downto 0));
   end component;
   
   component 
      CwGenerator_DATA_SIZE32_OPCD_SIZE6_FUNC_SIZE11_CWRD_SIZE20_CALU_SIZE5
      port( clk, rst : in std_logic;  opcd : in std_logic_vector (5 downto 0); 
            func : in std_logic_vector (10 downto 0);  stall_flag : in 
            std_logic_vector (4 downto 0);  taken : in std_logic;  cw : out 
            std_logic_vector (19 downto 0);  calu : out std_logic_vector (4 
            downto 0));
   end component;
   
   signal sig_bpw_port, stall_flag_4_port, stall_flag_3_port, stall_flag_2_port
      , stall_flag_1_port, stall_flag_0_port, sig_brt, net107957, net107958, 
      net107959, net107960, net107961, net107962, net107963, net107964, 
      net107965, net107966, net107967, net107968, net107969, net107970, 
      net107971, net107972, net107973, net107974 : std_logic;

begin
   sig_bpw <= sig_bpw_port;
   
   CW_GEN : 
                           CwGenerator_DATA_SIZE32_OPCD_SIZE6_FUNC_SIZE11_CWRD_SIZE20_CALU_SIZE5 
                           port map( clk => clk, rst => rst, opcd(5) => ir(31),
                           opcd(4) => ir(30), opcd(3) => ir(29), opcd(2) => 
                           ir(28), opcd(1) => ir(27), opcd(0) => ir(26), 
                           func(10) => ir(10), func(9) => ir(9), func(8) => 
                           ir(8), func(7) => ir(7), func(6) => ir(6), func(5) 
                           => ir(5), func(4) => ir(4), func(3) => ir(3), 
                           func(2) => ir(2), func(1) => ir(1), func(0) => ir(0)
                           , stall_flag(4) => stall_flag_4_port, stall_flag(3) 
                           => stall_flag_3_port, stall_flag(2) => 
                           stall_flag_2_port, stall_flag(1) => 
                           stall_flag_1_port, stall_flag(0) => 
                           stall_flag_0_port, taken => sig_brt, cw(19) => 
                           net107957, cw(18) => net107958, cw(17) => net107959,
                           cw(16) => net107960, cw(15) => net107961, cw(14) => 
                           net107962, cw(13) => net107963, cw(12) => net107964,
                           cw(11) => net107965, cw(10) => net107966, cw(9) => 
                           net107967, cw(8) => net107968, cw(7) => net107969, 
                           cw(6) => net107970, cw(5) => net107971, cw(4) => 
                           net107972, cw(3) => net107973, cw(2) => net107974, 
                           cw(1) => cw(1), cw(0) => cw(0), calu(4) => calu(4), 
                           calu(3) => calu(3), calu(2) => calu(2), calu(1) => 
                           calu(1), calu(0) => calu(0));
   S_GEN : StallGenerator_CWRD_SIZE20 port map( rst => rst, clk => clk, sig_ral
                           => sig_ral, sig_bpw => sig_bpw_port, sig_jral => 
                           sig_jral, sig_mul => sig_mul, sig_div => sig_div, 
                           sig_sqrt => sig_sqrt, stall_flag(4) => 
                           stall_flag_4_port, stall_flag(3) => 
                           stall_flag_3_port, stall_flag(2) => 
                           stall_flag_2_port, stall_flag(1) => 
                           stall_flag_1_port, stall_flag(0) => 
                           stall_flag_0_port);
   BR : Branch_DATA_SIZE32_OPCD_SIZE6_ADDR_SIZE32 port map( rst => rst, clk => 
                           clk, reg_a(31) => reg_a(31), reg_a(30) => reg_a(30),
                           reg_a(29) => reg_a(29), reg_a(28) => reg_a(28), 
                           reg_a(27) => reg_a(27), reg_a(26) => reg_a(26), 
                           reg_a(25) => reg_a(25), reg_a(24) => reg_a(24), 
                           reg_a(23) => reg_a(23), reg_a(22) => reg_a(22), 
                           reg_a(21) => reg_a(21), reg_a(20) => reg_a(20), 
                           reg_a(19) => reg_a(19), reg_a(18) => reg_a(18), 
                           reg_a(17) => reg_a(17), reg_a(16) => reg_a(16), 
                           reg_a(15) => reg_a(15), reg_a(14) => reg_a(14), 
                           reg_a(13) => reg_a(13), reg_a(12) => reg_a(12), 
                           reg_a(11) => reg_a(11), reg_a(10) => reg_a(10), 
                           reg_a(9) => reg_a(9), reg_a(8) => reg_a(8), reg_a(7)
                           => reg_a(7), reg_a(6) => reg_a(6), reg_a(5) => 
                           reg_a(5), reg_a(4) => reg_a(4), reg_a(3) => reg_a(3)
                           , reg_a(2) => reg_a(2), reg_a(1) => reg_a(1), 
                           reg_a(0) => reg_a(0), ld_a(31) => ld_a(31), ld_a(30)
                           => ld_a(30), ld_a(29) => ld_a(29), ld_a(28) => 
                           ld_a(28), ld_a(27) => ld_a(27), ld_a(26) => ld_a(26)
                           , ld_a(25) => ld_a(25), ld_a(24) => ld_a(24), 
                           ld_a(23) => ld_a(23), ld_a(22) => ld_a(22), ld_a(21)
                           => ld_a(21), ld_a(20) => ld_a(20), ld_a(19) => 
                           ld_a(19), ld_a(18) => ld_a(18), ld_a(17) => ld_a(17)
                           , ld_a(16) => ld_a(16), ld_a(15) => ld_a(15), 
                           ld_a(14) => ld_a(14), ld_a(13) => ld_a(13), ld_a(12)
                           => ld_a(12), ld_a(11) => ld_a(11), ld_a(10) => 
                           ld_a(10), ld_a(9) => ld_a(9), ld_a(8) => ld_a(8), 
                           ld_a(7) => ld_a(7), ld_a(6) => ld_a(6), ld_a(5) => 
                           ld_a(5), ld_a(4) => ld_a(4), ld_a(3) => ld_a(3), 
                           ld_a(2) => ld_a(2), ld_a(1) => ld_a(1), ld_a(0) => 
                           ld_a(0), opcd(5) => ir(31), opcd(4) => ir(30), 
                           opcd(3) => ir(29), opcd(2) => ir(28), opcd(1) => 
                           ir(27), opcd(0) => ir(26), addr(31) => pc(31), 
                           addr(30) => pc(30), addr(29) => pc(29), addr(28) => 
                           pc(28), addr(27) => pc(27), addr(26) => pc(26), 
                           addr(25) => pc(25), addr(24) => pc(24), addr(23) => 
                           pc(23), addr(22) => pc(22), addr(21) => pc(21), 
                           addr(20) => pc(20), addr(19) => pc(19), addr(18) => 
                           pc(18), addr(17) => pc(17), addr(16) => pc(16), 
                           addr(15) => pc(15), addr(14) => pc(14), addr(13) => 
                           pc(13), addr(12) => pc(12), addr(11) => pc(11), 
                           addr(10) => pc(10), addr(9) => pc(9), addr(8) => 
                           pc(8), addr(7) => pc(7), addr(6) => pc(6), addr(5) 
                           => pc(5), addr(4) => pc(4), addr(3) => pc(3), 
                           addr(2) => pc(2), addr(1) => pc(1), addr(0) => pc(0)
                           , sig_bal => sig_bal, sig_bpw => sig_bpw_port, 
                           sig_brt => sig_brt);
   cw(2) <= '0';
   cw(3) <= '0';
   cw(4) <= '0';
   cw(5) <= '0';
   cw(6) <= '0';
   cw(7) <= '0';
   cw(8) <= '0';
   cw(9) <= '0';
   cw(10) <= '0';
   cw(11) <= '0';
   cw(12) <= '0';
   cw(13) <= '0';
   cw(14) <= '0';
   cw(15) <= '0';
   cw(16) <= '0';
   cw(17) <= '0';
   cw(18) <= '0';
   cw(19) <= '0';

end SYN_control_unit_arch;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4.all;

entity Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4 is

   port( clk, rst : in std_logic;  en_iram : out std_logic;  pc_bus : out 
         std_logic_vector (31 downto 0);  ir_bus : in std_logic_vector (31 
         downto 0);  en_dram : out std_logic;  addr_bus, di_bus : out 
         std_logic_vector (31 downto 0);  do_bus : in std_logic_vector (31 
         downto 0);  dr_cw : out std_logic_vector (3 downto 0));

end Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4;

architecture SYN_dlx_arch of Dlx_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_DRCW_SIZE4
   is

   component 
      DataPath_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_OPCD_SIZE6_IMME_SIZE16_CWRD_SIZE20_CALU_SIZE5_DRCW_SIZE4
      port( clk, rst : in std_logic;  istr_addr : out std_logic_vector (31 
            downto 0);  istr_val : in std_logic_vector (31 downto 0);  ir_out, 
            pc_out, reg_a_out, ld_a_out, data_addr : out std_logic_vector (31 
            downto 0);  data_i_val : in std_logic_vector (31 downto 0);  
            data_o_val : out std_logic_vector (31 downto 0);  cw : in 
            std_logic_vector (19 downto 0);  dr_cw : out std_logic_vector (3 
            downto 0);  calu : in std_logic_vector (4 downto 0);  sig_bal : out
            std_logic;  sig_bpw : in std_logic;  sig_jral, sig_ral, sig_mul, 
            sig_div, sig_sqrt : out std_logic);
   end component;
   
   component 
      ControlUnit_ISTR_SIZE32_DATA_SIZE32_OPCD_SIZE6_FUNC_SIZE11_CWRD_SIZE20_CALU_SIZE5_ADDR_SIZE32
      port( clk, rst : in std_logic;  ir, pc, reg_a, ld_a : in std_logic_vector
            (31 downto 0);  sig_bal : in std_logic;  sig_bpw : out std_logic;  
            sig_jral, sig_ral, sig_mul, sig_div, sig_sqrt : in std_logic;  cw :
            out std_logic_vector (19 downto 0);  calu : out std_logic_vector (4
            downto 0));
   end component;
   
   signal en_iram_port, ir_31_port, ir_30_port, ir_29_port, ir_28_port, 
      ir_27_port, ir_26_port, ir_25_port, ir_24_port, ir_23_port, ir_22_port, 
      ir_21_port, ir_20_port, ir_19_port, ir_18_port, ir_17_port, ir_16_port, 
      ir_15_port, ir_14_port, ir_13_port, ir_12_port, ir_11_port, ir_10_port, 
      ir_9_port, ir_8_port, ir_7_port, ir_6_port, ir_5_port, ir_4_port, 
      ir_3_port, ir_2_port, ir_1_port, ir_0_port, pc_31_port, pc_30_port, 
      pc_29_port, pc_28_port, pc_27_port, pc_26_port, pc_25_port, pc_24_port, 
      pc_23_port, pc_22_port, pc_21_port, pc_20_port, pc_19_port, pc_18_port, 
      pc_17_port, pc_16_port, pc_15_port, pc_14_port, pc_13_port, pc_12_port, 
      pc_11_port, pc_10_port, pc_9_port, pc_8_port, pc_7_port, pc_6_port, 
      pc_5_port, pc_4_port, pc_3_port, pc_2_port, pc_1_port, pc_0_port, 
      reg_a_val_31_port, reg_a_val_30_port, reg_a_val_29_port, 
      reg_a_val_28_port, reg_a_val_27_port, reg_a_val_26_port, 
      reg_a_val_25_port, reg_a_val_24_port, reg_a_val_23_port, 
      reg_a_val_22_port, reg_a_val_21_port, reg_a_val_20_port, 
      reg_a_val_19_port, reg_a_val_18_port, reg_a_val_17_port, 
      reg_a_val_16_port, reg_a_val_15_port, reg_a_val_14_port, 
      reg_a_val_13_port, reg_a_val_12_port, reg_a_val_11_port, 
      reg_a_val_10_port, reg_a_val_9_port, reg_a_val_8_port, reg_a_val_7_port, 
      reg_a_val_6_port, reg_a_val_5_port, reg_a_val_4_port, reg_a_val_3_port, 
      reg_a_val_2_port, reg_a_val_1_port, reg_a_val_0_port, ld_a_val_31_port, 
      ld_a_val_30_port, ld_a_val_29_port, ld_a_val_28_port, ld_a_val_27_port, 
      ld_a_val_26_port, ld_a_val_25_port, ld_a_val_24_port, ld_a_val_23_port, 
      ld_a_val_22_port, ld_a_val_21_port, ld_a_val_20_port, ld_a_val_19_port, 
      ld_a_val_18_port, ld_a_val_17_port, ld_a_val_16_port, ld_a_val_15_port, 
      ld_a_val_14_port, ld_a_val_13_port, ld_a_val_12_port, ld_a_val_11_port, 
      ld_a_val_10_port, ld_a_val_9_port, ld_a_val_8_port, ld_a_val_7_port, 
      ld_a_val_6_port, ld_a_val_5_port, ld_a_val_4_port, ld_a_val_3_port, 
      ld_a_val_2_port, ld_a_val_1_port, ld_a_val_0_port, sig_bal, sig_bpw, 
      sig_jral, sig_ral, sig_mul, sig_div, sig_sqrt, cw_19_port, cw_18_port, 
      cw_17_port, cw_16_port, cw_15_port, cw_14_port, cw_13_port, cw_12_port, 
      cw_11_port, cw_10_port, cw_9_port, cw_8_port, cw_7_port, cw_6_port, 
      cw_5_port, cw_4_port, cw_3_port, cw_2_port, cw_1_port, calu_4_port, 
      calu_3_port, calu_2_port, calu_1_port, calu_0_port, net107939, net107940,
      net107941, net107942, net107943, net107944, net107945, net107946, 
      net107947, net107948, net107949, net107950, net107951, net107952, 
      net107953, net107954, net107955, net107956 : std_logic;

begin
   en_iram <= en_iram_port;
   
   en_dram <= '1';
   CU0 : 
                           ControlUnit_ISTR_SIZE32_DATA_SIZE32_OPCD_SIZE6_FUNC_SIZE11_CWRD_SIZE20_CALU_SIZE5_ADDR_SIZE32 
                           port map( clk => clk, rst => rst, ir(31) => 
                           ir_31_port, ir(30) => ir_30_port, ir(29) => 
                           ir_29_port, ir(28) => ir_28_port, ir(27) => 
                           ir_27_port, ir(26) => ir_26_port, ir(25) => 
                           ir_25_port, ir(24) => ir_24_port, ir(23) => 
                           ir_23_port, ir(22) => ir_22_port, ir(21) => 
                           ir_21_port, ir(20) => ir_20_port, ir(19) => 
                           ir_19_port, ir(18) => ir_18_port, ir(17) => 
                           ir_17_port, ir(16) => ir_16_port, ir(15) => 
                           ir_15_port, ir(14) => ir_14_port, ir(13) => 
                           ir_13_port, ir(12) => ir_12_port, ir(11) => 
                           ir_11_port, ir(10) => ir_10_port, ir(9) => ir_9_port
                           , ir(8) => ir_8_port, ir(7) => ir_7_port, ir(6) => 
                           ir_6_port, ir(5) => ir_5_port, ir(4) => ir_4_port, 
                           ir(3) => ir_3_port, ir(2) => ir_2_port, ir(1) => 
                           ir_1_port, ir(0) => ir_0_port, pc(31) => pc_31_port,
                           pc(30) => pc_30_port, pc(29) => pc_29_port, pc(28) 
                           => pc_28_port, pc(27) => pc_27_port, pc(26) => 
                           pc_26_port, pc(25) => pc_25_port, pc(24) => 
                           pc_24_port, pc(23) => pc_23_port, pc(22) => 
                           pc_22_port, pc(21) => pc_21_port, pc(20) => 
                           pc_20_port, pc(19) => pc_19_port, pc(18) => 
                           pc_18_port, pc(17) => pc_17_port, pc(16) => 
                           pc_16_port, pc(15) => pc_15_port, pc(14) => 
                           pc_14_port, pc(13) => pc_13_port, pc(12) => 
                           pc_12_port, pc(11) => pc_11_port, pc(10) => 
                           pc_10_port, pc(9) => pc_9_port, pc(8) => pc_8_port, 
                           pc(7) => pc_7_port, pc(6) => pc_6_port, pc(5) => 
                           pc_5_port, pc(4) => pc_4_port, pc(3) => pc_3_port, 
                           pc(2) => pc_2_port, pc(1) => pc_1_port, pc(0) => 
                           pc_0_port, reg_a(31) => reg_a_val_31_port, reg_a(30)
                           => reg_a_val_30_port, reg_a(29) => reg_a_val_29_port
                           , reg_a(28) => reg_a_val_28_port, reg_a(27) => 
                           reg_a_val_27_port, reg_a(26) => reg_a_val_26_port, 
                           reg_a(25) => reg_a_val_25_port, reg_a(24) => 
                           reg_a_val_24_port, reg_a(23) => reg_a_val_23_port, 
                           reg_a(22) => reg_a_val_22_port, reg_a(21) => 
                           reg_a_val_21_port, reg_a(20) => reg_a_val_20_port, 
                           reg_a(19) => reg_a_val_19_port, reg_a(18) => 
                           reg_a_val_18_port, reg_a(17) => reg_a_val_17_port, 
                           reg_a(16) => reg_a_val_16_port, reg_a(15) => 
                           reg_a_val_15_port, reg_a(14) => reg_a_val_14_port, 
                           reg_a(13) => reg_a_val_13_port, reg_a(12) => 
                           reg_a_val_12_port, reg_a(11) => reg_a_val_11_port, 
                           reg_a(10) => reg_a_val_10_port, reg_a(9) => 
                           reg_a_val_9_port, reg_a(8) => reg_a_val_8_port, 
                           reg_a(7) => reg_a_val_7_port, reg_a(6) => 
                           reg_a_val_6_port, reg_a(5) => reg_a_val_5_port, 
                           reg_a(4) => reg_a_val_4_port, reg_a(3) => 
                           reg_a_val_3_port, reg_a(2) => reg_a_val_2_port, 
                           reg_a(1) => reg_a_val_1_port, reg_a(0) => 
                           reg_a_val_0_port, ld_a(31) => ld_a_val_31_port, 
                           ld_a(30) => ld_a_val_30_port, ld_a(29) => 
                           ld_a_val_29_port, ld_a(28) => ld_a_val_28_port, 
                           ld_a(27) => ld_a_val_27_port, ld_a(26) => 
                           ld_a_val_26_port, ld_a(25) => ld_a_val_25_port, 
                           ld_a(24) => ld_a_val_24_port, ld_a(23) => 
                           ld_a_val_23_port, ld_a(22) => ld_a_val_22_port, 
                           ld_a(21) => ld_a_val_21_port, ld_a(20) => 
                           ld_a_val_20_port, ld_a(19) => ld_a_val_19_port, 
                           ld_a(18) => ld_a_val_18_port, ld_a(17) => 
                           ld_a_val_17_port, ld_a(16) => ld_a_val_16_port, 
                           ld_a(15) => ld_a_val_15_port, ld_a(14) => 
                           ld_a_val_14_port, ld_a(13) => ld_a_val_13_port, 
                           ld_a(12) => ld_a_val_12_port, ld_a(11) => 
                           ld_a_val_11_port, ld_a(10) => ld_a_val_10_port, 
                           ld_a(9) => ld_a_val_9_port, ld_a(8) => 
                           ld_a_val_8_port, ld_a(7) => ld_a_val_7_port, ld_a(6)
                           => ld_a_val_6_port, ld_a(5) => ld_a_val_5_port, 
                           ld_a(4) => ld_a_val_4_port, ld_a(3) => 
                           ld_a_val_3_port, ld_a(2) => ld_a_val_2_port, ld_a(1)
                           => ld_a_val_1_port, ld_a(0) => ld_a_val_0_port, 
                           sig_bal => sig_bal, sig_bpw => sig_bpw, sig_jral => 
                           sig_jral, sig_ral => sig_ral, sig_mul => sig_mul, 
                           sig_div => sig_div, sig_sqrt => sig_sqrt, cw(19) => 
                           net107939, cw(18) => net107940, cw(17) => net107941,
                           cw(16) => net107942, cw(15) => net107943, cw(14) => 
                           net107944, cw(13) => net107945, cw(12) => net107946,
                           cw(11) => net107947, cw(10) => net107948, cw(9) => 
                           net107949, cw(8) => net107950, cw(7) => net107951, 
                           cw(6) => net107952, cw(5) => net107953, cw(4) => 
                           net107954, cw(3) => net107955, cw(2) => net107956, 
                           cw(1) => cw_1_port, cw(0) => en_iram_port, calu(4) 
                           => calu_4_port, calu(3) => calu_3_port, calu(2) => 
                           calu_2_port, calu(1) => calu_1_port, calu(0) => 
                           calu_0_port);
   DP0 : 
                           DataPath_ADDR_SIZE32_DATA_SIZE32_ISTR_SIZE32_OPCD_SIZE6_IMME_SIZE16_CWRD_SIZE20_CALU_SIZE5_DRCW_SIZE4 
                           port map( clk => clk, rst => rst, istr_addr(31) => 
                           pc_bus(31), istr_addr(30) => pc_bus(30), 
                           istr_addr(29) => pc_bus(29), istr_addr(28) => 
                           pc_bus(28), istr_addr(27) => pc_bus(27), 
                           istr_addr(26) => pc_bus(26), istr_addr(25) => 
                           pc_bus(25), istr_addr(24) => pc_bus(24), 
                           istr_addr(23) => pc_bus(23), istr_addr(22) => 
                           pc_bus(22), istr_addr(21) => pc_bus(21), 
                           istr_addr(20) => pc_bus(20), istr_addr(19) => 
                           pc_bus(19), istr_addr(18) => pc_bus(18), 
                           istr_addr(17) => pc_bus(17), istr_addr(16) => 
                           pc_bus(16), istr_addr(15) => pc_bus(15), 
                           istr_addr(14) => pc_bus(14), istr_addr(13) => 
                           pc_bus(13), istr_addr(12) => pc_bus(12), 
                           istr_addr(11) => pc_bus(11), istr_addr(10) => 
                           pc_bus(10), istr_addr(9) => pc_bus(9), istr_addr(8) 
                           => pc_bus(8), istr_addr(7) => pc_bus(7), 
                           istr_addr(6) => pc_bus(6), istr_addr(5) => pc_bus(5)
                           , istr_addr(4) => pc_bus(4), istr_addr(3) => 
                           pc_bus(3), istr_addr(2) => pc_bus(2), istr_addr(1) 
                           => pc_bus(1), istr_addr(0) => pc_bus(0), 
                           istr_val(31) => ir_bus(31), istr_val(30) => 
                           ir_bus(30), istr_val(29) => ir_bus(29), istr_val(28)
                           => ir_bus(28), istr_val(27) => ir_bus(27), 
                           istr_val(26) => ir_bus(26), istr_val(25) => 
                           ir_bus(25), istr_val(24) => ir_bus(24), istr_val(23)
                           => ir_bus(23), istr_val(22) => ir_bus(22), 
                           istr_val(21) => ir_bus(21), istr_val(20) => 
                           ir_bus(20), istr_val(19) => ir_bus(19), istr_val(18)
                           => ir_bus(18), istr_val(17) => ir_bus(17), 
                           istr_val(16) => ir_bus(16), istr_val(15) => 
                           ir_bus(15), istr_val(14) => ir_bus(14), istr_val(13)
                           => ir_bus(13), istr_val(12) => ir_bus(12), 
                           istr_val(11) => ir_bus(11), istr_val(10) => 
                           ir_bus(10), istr_val(9) => ir_bus(9), istr_val(8) =>
                           ir_bus(8), istr_val(7) => ir_bus(7), istr_val(6) => 
                           ir_bus(6), istr_val(5) => ir_bus(5), istr_val(4) => 
                           ir_bus(4), istr_val(3) => ir_bus(3), istr_val(2) => 
                           ir_bus(2), istr_val(1) => ir_bus(1), istr_val(0) => 
                           ir_bus(0), ir_out(31) => ir_31_port, ir_out(30) => 
                           ir_30_port, ir_out(29) => ir_29_port, ir_out(28) => 
                           ir_28_port, ir_out(27) => ir_27_port, ir_out(26) => 
                           ir_26_port, ir_out(25) => ir_25_port, ir_out(24) => 
                           ir_24_port, ir_out(23) => ir_23_port, ir_out(22) => 
                           ir_22_port, ir_out(21) => ir_21_port, ir_out(20) => 
                           ir_20_port, ir_out(19) => ir_19_port, ir_out(18) => 
                           ir_18_port, ir_out(17) => ir_17_port, ir_out(16) => 
                           ir_16_port, ir_out(15) => ir_15_port, ir_out(14) => 
                           ir_14_port, ir_out(13) => ir_13_port, ir_out(12) => 
                           ir_12_port, ir_out(11) => ir_11_port, ir_out(10) => 
                           ir_10_port, ir_out(9) => ir_9_port, ir_out(8) => 
                           ir_8_port, ir_out(7) => ir_7_port, ir_out(6) => 
                           ir_6_port, ir_out(5) => ir_5_port, ir_out(4) => 
                           ir_4_port, ir_out(3) => ir_3_port, ir_out(2) => 
                           ir_2_port, ir_out(1) => ir_1_port, ir_out(0) => 
                           ir_0_port, pc_out(31) => pc_31_port, pc_out(30) => 
                           pc_30_port, pc_out(29) => pc_29_port, pc_out(28) => 
                           pc_28_port, pc_out(27) => pc_27_port, pc_out(26) => 
                           pc_26_port, pc_out(25) => pc_25_port, pc_out(24) => 
                           pc_24_port, pc_out(23) => pc_23_port, pc_out(22) => 
                           pc_22_port, pc_out(21) => pc_21_port, pc_out(20) => 
                           pc_20_port, pc_out(19) => pc_19_port, pc_out(18) => 
                           pc_18_port, pc_out(17) => pc_17_port, pc_out(16) => 
                           pc_16_port, pc_out(15) => pc_15_port, pc_out(14) => 
                           pc_14_port, pc_out(13) => pc_13_port, pc_out(12) => 
                           pc_12_port, pc_out(11) => pc_11_port, pc_out(10) => 
                           pc_10_port, pc_out(9) => pc_9_port, pc_out(8) => 
                           pc_8_port, pc_out(7) => pc_7_port, pc_out(6) => 
                           pc_6_port, pc_out(5) => pc_5_port, pc_out(4) => 
                           pc_4_port, pc_out(3) => pc_3_port, pc_out(2) => 
                           pc_2_port, pc_out(1) => pc_1_port, pc_out(0) => 
                           pc_0_port, reg_a_out(31) => reg_a_val_31_port, 
                           reg_a_out(30) => reg_a_val_30_port, reg_a_out(29) =>
                           reg_a_val_29_port, reg_a_out(28) => 
                           reg_a_val_28_port, reg_a_out(27) => 
                           reg_a_val_27_port, reg_a_out(26) => 
                           reg_a_val_26_port, reg_a_out(25) => 
                           reg_a_val_25_port, reg_a_out(24) => 
                           reg_a_val_24_port, reg_a_out(23) => 
                           reg_a_val_23_port, reg_a_out(22) => 
                           reg_a_val_22_port, reg_a_out(21) => 
                           reg_a_val_21_port, reg_a_out(20) => 
                           reg_a_val_20_port, reg_a_out(19) => 
                           reg_a_val_19_port, reg_a_out(18) => 
                           reg_a_val_18_port, reg_a_out(17) => 
                           reg_a_val_17_port, reg_a_out(16) => 
                           reg_a_val_16_port, reg_a_out(15) => 
                           reg_a_val_15_port, reg_a_out(14) => 
                           reg_a_val_14_port, reg_a_out(13) => 
                           reg_a_val_13_port, reg_a_out(12) => 
                           reg_a_val_12_port, reg_a_out(11) => 
                           reg_a_val_11_port, reg_a_out(10) => 
                           reg_a_val_10_port, reg_a_out(9) => reg_a_val_9_port,
                           reg_a_out(8) => reg_a_val_8_port, reg_a_out(7) => 
                           reg_a_val_7_port, reg_a_out(6) => reg_a_val_6_port, 
                           reg_a_out(5) => reg_a_val_5_port, reg_a_out(4) => 
                           reg_a_val_4_port, reg_a_out(3) => reg_a_val_3_port, 
                           reg_a_out(2) => reg_a_val_2_port, reg_a_out(1) => 
                           reg_a_val_1_port, reg_a_out(0) => reg_a_val_0_port, 
                           ld_a_out(31) => ld_a_val_31_port, ld_a_out(30) => 
                           ld_a_val_30_port, ld_a_out(29) => ld_a_val_29_port, 
                           ld_a_out(28) => ld_a_val_28_port, ld_a_out(27) => 
                           ld_a_val_27_port, ld_a_out(26) => ld_a_val_26_port, 
                           ld_a_out(25) => ld_a_val_25_port, ld_a_out(24) => 
                           ld_a_val_24_port, ld_a_out(23) => ld_a_val_23_port, 
                           ld_a_out(22) => ld_a_val_22_port, ld_a_out(21) => 
                           ld_a_val_21_port, ld_a_out(20) => ld_a_val_20_port, 
                           ld_a_out(19) => ld_a_val_19_port, ld_a_out(18) => 
                           ld_a_val_18_port, ld_a_out(17) => ld_a_val_17_port, 
                           ld_a_out(16) => ld_a_val_16_port, ld_a_out(15) => 
                           ld_a_val_15_port, ld_a_out(14) => ld_a_val_14_port, 
                           ld_a_out(13) => ld_a_val_13_port, ld_a_out(12) => 
                           ld_a_val_12_port, ld_a_out(11) => ld_a_val_11_port, 
                           ld_a_out(10) => ld_a_val_10_port, ld_a_out(9) => 
                           ld_a_val_9_port, ld_a_out(8) => ld_a_val_8_port, 
                           ld_a_out(7) => ld_a_val_7_port, ld_a_out(6) => 
                           ld_a_val_6_port, ld_a_out(5) => ld_a_val_5_port, 
                           ld_a_out(4) => ld_a_val_4_port, ld_a_out(3) => 
                           ld_a_val_3_port, ld_a_out(2) => ld_a_val_2_port, 
                           ld_a_out(1) => ld_a_val_1_port, ld_a_out(0) => 
                           ld_a_val_0_port, data_addr(31) => addr_bus(31), 
                           data_addr(30) => addr_bus(30), data_addr(29) => 
                           addr_bus(29), data_addr(28) => addr_bus(28), 
                           data_addr(27) => addr_bus(27), data_addr(26) => 
                           addr_bus(26), data_addr(25) => addr_bus(25), 
                           data_addr(24) => addr_bus(24), data_addr(23) => 
                           addr_bus(23), data_addr(22) => addr_bus(22), 
                           data_addr(21) => addr_bus(21), data_addr(20) => 
                           addr_bus(20), data_addr(19) => addr_bus(19), 
                           data_addr(18) => addr_bus(18), data_addr(17) => 
                           addr_bus(17), data_addr(16) => addr_bus(16), 
                           data_addr(15) => addr_bus(15), data_addr(14) => 
                           addr_bus(14), data_addr(13) => addr_bus(13), 
                           data_addr(12) => addr_bus(12), data_addr(11) => 
                           addr_bus(11), data_addr(10) => addr_bus(10), 
                           data_addr(9) => addr_bus(9), data_addr(8) => 
                           addr_bus(8), data_addr(7) => addr_bus(7), 
                           data_addr(6) => addr_bus(6), data_addr(5) => 
                           addr_bus(5), data_addr(4) => addr_bus(4), 
                           data_addr(3) => addr_bus(3), data_addr(2) => 
                           addr_bus(2), data_addr(1) => addr_bus(1), 
                           data_addr(0) => addr_bus(0), data_i_val(31) => 
                           do_bus(31), data_i_val(30) => do_bus(30), 
                           data_i_val(29) => do_bus(29), data_i_val(28) => 
                           do_bus(28), data_i_val(27) => do_bus(27), 
                           data_i_val(26) => do_bus(26), data_i_val(25) => 
                           do_bus(25), data_i_val(24) => do_bus(24), 
                           data_i_val(23) => do_bus(23), data_i_val(22) => 
                           do_bus(22), data_i_val(21) => do_bus(21), 
                           data_i_val(20) => do_bus(20), data_i_val(19) => 
                           do_bus(19), data_i_val(18) => do_bus(18), 
                           data_i_val(17) => do_bus(17), data_i_val(16) => 
                           do_bus(16), data_i_val(15) => do_bus(15), 
                           data_i_val(14) => do_bus(14), data_i_val(13) => 
                           do_bus(13), data_i_val(12) => do_bus(12), 
                           data_i_val(11) => do_bus(11), data_i_val(10) => 
                           do_bus(10), data_i_val(9) => do_bus(9), 
                           data_i_val(8) => do_bus(8), data_i_val(7) => 
                           do_bus(7), data_i_val(6) => do_bus(6), data_i_val(5)
                           => do_bus(5), data_i_val(4) => do_bus(4), 
                           data_i_val(3) => do_bus(3), data_i_val(2) => 
                           do_bus(2), data_i_val(1) => do_bus(1), data_i_val(0)
                           => do_bus(0), data_o_val(31) => di_bus(31), 
                           data_o_val(30) => di_bus(30), data_o_val(29) => 
                           di_bus(29), data_o_val(28) => di_bus(28), 
                           data_o_val(27) => di_bus(27), data_o_val(26) => 
                           di_bus(26), data_o_val(25) => di_bus(25), 
                           data_o_val(24) => di_bus(24), data_o_val(23) => 
                           di_bus(23), data_o_val(22) => di_bus(22), 
                           data_o_val(21) => di_bus(21), data_o_val(20) => 
                           di_bus(20), data_o_val(19) => di_bus(19), 
                           data_o_val(18) => di_bus(18), data_o_val(17) => 
                           di_bus(17), data_o_val(16) => di_bus(16), 
                           data_o_val(15) => di_bus(15), data_o_val(14) => 
                           di_bus(14), data_o_val(13) => di_bus(13), 
                           data_o_val(12) => di_bus(12), data_o_val(11) => 
                           di_bus(11), data_o_val(10) => di_bus(10), 
                           data_o_val(9) => di_bus(9), data_o_val(8) => 
                           di_bus(8), data_o_val(7) => di_bus(7), data_o_val(6)
                           => di_bus(6), data_o_val(5) => di_bus(5), 
                           data_o_val(4) => di_bus(4), data_o_val(3) => 
                           di_bus(3), data_o_val(2) => di_bus(2), data_o_val(1)
                           => di_bus(1), data_o_val(0) => di_bus(0), cw(19) => 
                           cw_19_port, cw(18) => cw_18_port, cw(17) => 
                           cw_17_port, cw(16) => cw_16_port, cw(15) => 
                           cw_15_port, cw(14) => cw_14_port, cw(13) => 
                           cw_13_port, cw(12) => cw_12_port, cw(11) => 
                           cw_11_port, cw(10) => cw_10_port, cw(9) => cw_9_port
                           , cw(8) => cw_8_port, cw(7) => cw_7_port, cw(6) => 
                           cw_6_port, cw(5) => cw_5_port, cw(4) => cw_4_port, 
                           cw(3) => cw_3_port, cw(2) => cw_2_port, cw(1) => 
                           cw_1_port, cw(0) => en_iram_port, dr_cw(3) => 
                           dr_cw(3), dr_cw(2) => dr_cw(2), dr_cw(1) => dr_cw(1)
                           , dr_cw(0) => dr_cw(0), calu(4) => calu_4_port, 
                           calu(3) => calu_3_port, calu(2) => calu_2_port, 
                           calu(1) => calu_1_port, calu(0) => calu_0_port, 
                           sig_bal => sig_bal, sig_bpw => sig_bpw, sig_jral => 
                           sig_jral, sig_ral => sig_ral, sig_mul => sig_mul, 
                           sig_div => sig_div, sig_sqrt => sig_sqrt);
   cw_2_port <= '0';
   cw_3_port <= '0';
   cw_4_port <= '0';
   cw_5_port <= '0';
   cw_6_port <= '0';
   cw_7_port <= '0';
   cw_8_port <= '0';
   cw_9_port <= '0';
   cw_10_port <= '0';
   cw_11_port <= '0';
   cw_12_port <= '0';
   cw_13_port <= '0';
   cw_14_port <= '0';
   cw_15_port <= '0';
   cw_16_port <= '0';
   cw_17_port <= '0';
   cw_18_port <= '0';
   cw_19_port <= '0';

end SYN_dlx_arch;
