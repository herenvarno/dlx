--------------------------------------------------------------------------------
-- FILE: Types
-- DESC: Define all types.
--
-- Author:
-- Create: 2015-05-20
-- Update: 2015-05-20
-- Status: TESTED
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

package Types is

end Types;

